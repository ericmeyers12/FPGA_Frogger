module images/lilypad_sprite(output logic [9:0] rgb[0:39][0:39]);
assign rgb = '{
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd380,9'd380,9'd380,9'd380,9'd380,9'd380,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
},
'{
9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379,9'd379
}};
endmodule
