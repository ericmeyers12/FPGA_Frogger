module logo(output logic [5:0] rgb[0:152][0:39]);
assign rgb = '{
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
}};
endmodule
