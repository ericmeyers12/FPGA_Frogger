module InvShiftRows(input logic [0:127] in, output logic[0:127] out);
   assign out = {
                 in[0:7], in[104:111], in[80:87], in[56:63],
                 in[32:39], in[8:15], in[112:119], in[88:95],
                 in[64:71], in[40:47], in[16:23], in[120:127],
                 in[96:103], in[72:79], in[48:55], in[24:31]
                 };
endmodule
