module palette(output logic [7:0] palette[0:18][0:2]);
assign palette = '{'{8'd0,8'd0,8'd0},'{8'd30,8'd130,8'd0},'{8'd0,8'd20,8'd0},'{8'd30,8'd150,8'd0},'{8'd50,8'd150,8'd20},'{8'd40,8'd150,8'd10},'{8'd20,8'd90,8'd0},'{8'd30,8'd140,8'd0},'{8'd40,8'd140,8'd0},'{8'd160,8'd40,8'd0},'{8'd250,8'd0,8'd0},'{8'd70,8'd70,8'd70},'{8'd250,8'd40,8'd0},'{8'd0,8'd80,8'd250},'{8'd250,8'd250,8'd250},'{8'd250,8'd230,8'd0},'{8'd180,8'd140,8'd20},'{8'd250,8'd10,8'd10},'{8'd0,8'd0,8'd0}};
endmodule
