module images/car_left(output logic [17:0] rgb[0:79][0:39]);
assign rgb = '{
'{
17'd0,17'd0,17'd0,17'd0,17'd0,17'd0,17'd67641,17'd67642,17'd67643,17'd67644,17'd67645,17'd67646,17'd67647,17'd67648,17'd67649,17'd67650,17'd67651,17'd67652,17'd67653,17'd67654,17'd67655,17'd67656,17'd67657,17'd67658,17'd67659,17'd67660,17'd67661,17'd67662,17'd67663,17'd67664,17'd67665,17'd67666,17'd67667,17'd0,17'd0,17'd0,17'd0,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd0,17'd0,17'd0,17'd0,17'd67668,17'd67669,17'd67670,17'd67671,17'd67672,17'd67673,17'd67674,17'd67675,17'd67676,17'd67677,17'd67678,17'd67679,17'd67680,17'd67681,17'd67682,17'd67683,17'd67684,17'd67685,17'd67686,17'd67687,17'd67688,17'd67689,17'd67690,17'd67691,17'd67692,17'd67693,17'd67694,17'd49164,17'd0,17'd0,17'd0,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd0,17'd0,17'd0,17'd67695,17'd67696,17'd67697,17'd67698,17'd67699,17'd67700,17'd67701,17'd67702,17'd67703,17'd67704,17'd67705,17'd67706,17'd67707,17'd67708,17'd67709,17'd67710,17'd67711,17'd67712,17'd67713,17'd67714,17'd67715,17'd67716,17'd67717,17'd67718,17'd67719,17'd67720,17'd67721,17'd67722,17'd67723,17'd0,17'd0,17'd0,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd0,17'd0,17'd67724,17'd67725,17'd67726,17'd67727,17'd67728,17'd67729,17'd67730,17'd67731,17'd67732,17'd67733,17'd67734,17'd67735,17'd67736,17'd67737,17'd67738,17'd67739,17'd67740,17'd67741,17'd67742,17'd67743,17'd67744,17'd67745,17'd67746,17'd67747,17'd67748,17'd67749,17'd67750,17'd67751,17'd67752,17'd67753,17'd67754,17'd0,17'd0,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd67755,17'd67756,17'd67757,17'd67758,17'd67759,17'd67760,17'd67761,17'd67762,17'd67763,17'd67764,17'd67765,17'd67766,17'd67766,17'd67767,17'd67768,17'd67769,17'd67770,17'd67771,17'd67740,17'd67772,17'd67773,17'd67774,17'd67775,17'd67776,17'd67777,17'd67778,17'd67779,17'd67780,17'd67781,17'd67782,17'd67783,17'd67784,17'd67785,17'd0,17'd0,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd67786,17'd67787,17'd67788,17'd67789,17'd67790,17'd67791,17'd67792,17'd67793,17'd67766,17'd67794,17'd67794,17'd67794,17'd67795,17'd67764,17'd67767,17'd67796,17'd67797,17'd67798,17'd67799,17'd67800,17'd67801,17'd67802,17'd67803,17'd67804,17'd67805,17'd67806,17'd67807,17'd67808,17'd67809,17'd67810,17'd63671,17'd67811,17'd67812,17'd67813,17'd0,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd67814,17'd67815,17'd67816,17'd67817,17'd67818,17'd67819,17'd67820,17'd67821,17'd67765,17'd67794,17'd67794,17'd67794,17'd67795,17'd67764,17'd67822,17'd67822,17'd67823,17'd67824,17'd67825,17'd67826,17'd67827,17'd67828,17'd67829,17'd67830,17'd67831,17'd67832,17'd67833,17'd67834,17'd67835,17'd67836,17'd67837,17'd67838,17'd67839,17'd67840,17'd0,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd67841,17'd67842,17'd67843,17'd67844,17'd67845,17'd67846,17'd67847,17'd67848,17'd67794,17'd67794,17'd67794,17'd67794,17'd67794,17'd67795,17'd67795,17'd67795,17'd67849,17'd67850,17'd67851,17'd67852,17'd67853,17'd67854,17'd67855,17'd67856,17'd67857,17'd67858,17'd67859,17'd67860,17'd67861,17'd67862,17'd67863,17'd67864,17'd67865,17'd67866,17'd67867,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd67868,17'd67869,17'd67870,17'd67871,17'd67872,17'd67873,17'd67874,17'd67875,17'd67874,17'd67848,17'd67794,17'd67794,17'd67794,17'd67794,17'd67764,17'd67795,17'd67849,17'd67850,17'd67851,17'd67876,17'd67877,17'd67878,17'd67879,17'd67880,17'd67881,17'd67882,17'd67883,17'd67884,17'd67885,17'd67886,17'd67887,17'd67888,17'd67889,17'd67890,17'd67891,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd67892,17'd67893,17'd67894,17'd67895,17'd67895,17'd67896,17'd67897,17'd67898,17'd67899,17'd67875,17'd67848,17'd67794,17'd67794,17'd67794,17'd67764,17'd67795,17'd67849,17'd67850,17'd67851,17'd67876,17'd67877,17'd67900,17'd67901,17'd67902,17'd67903,17'd67904,17'd67905,17'd67906,17'd67907,17'd67908,17'd67909,17'd67910,17'd67911,17'd67912,17'd67913,17'd67914,17'd0,17'd0
},
'{
17'd0,17'd0,17'd67915,17'd67916,17'd67917,17'd67896,17'd67896,17'd67874,17'd67918,17'd67919,17'd67920,17'd67875,17'd67794,17'd67794,17'd67794,17'd67794,17'd67764,17'd67795,17'd67849,17'd67921,17'd67851,17'd67876,17'd67877,17'd67900,17'd67901,17'd67880,17'd67922,17'd67923,17'd67924,17'd67925,17'd67926,17'd67927,17'd67928,17'd67929,17'd67930,17'd67931,17'd67932,17'd67933,17'd0,17'd0
},
'{
17'd0,17'd0,17'd67934,17'd67935,17'd67936,17'd67766,17'd67795,17'd67848,17'd67874,17'd67937,17'd67938,17'd67794,17'd67794,17'd67794,17'd67794,17'd67794,17'd67764,17'd67795,17'd67939,17'd67921,17'd67851,17'd67876,17'd67877,17'd67900,17'd67901,17'd67880,17'd67940,17'd67941,17'd67942,17'd67943,17'd67944,17'd67945,17'd67946,17'd67947,17'd67948,17'd67949,17'd67950,17'd67951,17'd0,17'd0
},
'{
17'd0,17'd0,17'd67952,17'd67953,17'd67954,17'd67764,17'd67848,17'd67874,17'd67955,17'd67899,17'd67956,17'd67874,17'd67794,17'd67794,17'd67794,17'd67794,17'd67764,17'd67795,17'd67849,17'd67921,17'd67851,17'd67876,17'd67877,17'd67900,17'd67901,17'd67957,17'd67958,17'd67959,17'd67960,17'd67961,17'd67962,17'd67963,17'd67964,17'd67778,17'd67965,17'd67966,17'd67967,17'd56726,17'd0,17'd0
},
'{
17'd0,17'd0,17'd67968,17'd67969,17'd67970,17'd67795,17'd67794,17'd67874,17'd67918,17'd67971,17'd67920,17'd67875,17'd67794,17'd67794,17'd67794,17'd67794,17'd67764,17'd67795,17'd67849,17'd67921,17'd67851,17'd67876,17'd67877,17'd67900,17'd67901,17'd67957,17'd67972,17'd67973,17'd67974,17'd67975,17'd67976,17'd67977,17'd67978,17'd67979,17'd67980,17'd67981,17'd43262,17'd67982,17'd0,17'd0
},
'{
17'd0,17'd0,17'd67983,17'd67984,17'd67942,17'd67795,17'd67794,17'd67848,17'd67875,17'd67985,17'd67938,17'd67794,17'd67794,17'd67794,17'd67794,17'd67794,17'd67764,17'd67795,17'd67849,17'd67850,17'd67851,17'd67876,17'd67877,17'd67900,17'd67901,17'd67986,17'd67987,17'd67988,17'd67985,17'd67989,17'd67990,17'd67991,17'd67992,17'd67993,17'd67994,17'd67995,17'd67996,17'd67997,17'd0,17'd0
},
'{
17'd0,17'd0,17'd67998,17'd67999,17'd68000,17'd68001,17'd67794,17'd67874,17'd67897,17'd67899,17'd67956,17'd67875,17'd67848,17'd67794,17'd67794,17'd67794,17'd67764,17'd67795,17'd67849,17'd67850,17'd67851,17'd67876,17'd67877,17'd67900,17'd67901,17'd67957,17'd68002,17'd68003,17'd67899,17'd68004,17'd68005,17'd68006,17'd68007,17'd68008,17'd68009,17'd68010,17'd68011,17'd68012,17'd0,17'd0
},
'{
17'd0,17'd0,17'd68013,17'd68014,17'd68015,17'd67765,17'd67794,17'd67874,17'd68016,17'd68017,17'd68018,17'd67875,17'd67794,17'd67794,17'd67794,17'd68019,17'd68001,17'd67765,17'd67849,17'd67921,17'd67851,17'd67876,17'd68020,17'd67900,17'd67901,17'd67957,17'd68021,17'd68022,17'd68023,17'd68024,17'd68025,17'd68026,17'd68027,17'd68028,17'd68029,17'd68030,17'd68031,17'd68032,17'd0,17'd0
},
'{
17'd0,17'd0,17'd68033,17'd68034,17'd68035,17'd67764,17'd68019,17'd67795,17'd68036,17'd68037,17'd67875,17'd67764,17'd67766,17'd67764,17'd67764,17'd68038,17'd68039,17'd68039,17'd67820,17'd68040,17'd68041,17'd68042,17'd68043,17'd68044,17'd68045,17'd68046,17'd68047,17'd68048,17'd68049,17'd68050,17'd68051,17'd68052,17'd68053,17'd68054,17'd68055,17'd68056,17'd68057,17'd68058,17'd0,17'd0
},
'{
17'd0,17'd0,17'd68059,17'd68060,17'd68061,17'd67765,17'd67795,17'd68062,17'd68063,17'd68064,17'd68065,17'd67733,17'd67733,17'd67733,17'd68066,17'd68067,17'd68068,17'd68069,17'd67877,17'd68070,17'd68071,17'd68072,17'd68073,17'd68074,17'd68075,17'd68076,17'd68077,17'd68078,17'd68079,17'd68080,17'd68068,17'd68081,17'd68082,17'd68083,17'd68084,17'd68085,17'd68086,17'd2185,17'd0,17'd0
},
'{
17'd0,17'd0,17'd68087,17'd68088,17'd68089,17'd67765,17'd67764,17'd68090,17'd68091,17'd68092,17'd68093,17'd68093,17'd68093,17'd68093,17'd68093,17'd68094,17'd68095,17'd68095,17'd68096,17'd68097,17'd68098,17'd68099,17'd68100,17'd68101,17'd68102,17'd68103,17'd68104,17'd68105,17'd68106,17'd68107,17'd68108,17'd68109,17'd68110,17'd68111,17'd68112,17'd68113,17'd68114,17'd68115,17'd0,17'd0
},
'{
17'd0,17'd0,17'd68116,17'd68117,17'd68118,17'd68119,17'd68120,17'd68121,17'd68122,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68124,17'd68125,17'd68126,17'd68127,17'd68128,17'd68129,17'd68130,17'd68114,17'd68131,17'd0,17'd0
},
'{
17'd0,17'd0,17'd68132,17'd68133,17'd68134,17'd68135,17'd68136,17'd68137,17'd68138,17'd68139,17'd68140,17'd68140,17'd68141,17'd68141,17'd68142,17'd68140,17'd68140,17'd68142,17'd68141,17'd68141,17'd68143,17'd68144,17'd68145,17'd68146,17'd68147,17'd68148,17'd68149,17'd68150,17'd68151,17'd68152,17'd68153,17'd68154,17'd68155,17'd68156,17'd68157,17'd68158,17'd68159,17'd62262,17'd0,17'd0
},
'{
17'd0,17'd0,17'd68160,17'd68161,17'd68162,17'd68163,17'd68164,17'd68123,17'd68165,17'd68166,17'd68167,17'd68168,17'd68168,17'd68168,17'd68169,17'd68170,17'd68171,17'd68169,17'd68168,17'd68170,17'd68172,17'd68173,17'd68174,17'd68175,17'd68176,17'd68177,17'd68178,17'd68179,17'd68180,17'd68181,17'd68123,17'd68123,17'd68182,17'd68183,17'd68184,17'd68185,17'd68186,17'd68187,17'd0,17'd0
},
'{
17'd0,17'd0,17'd68188,17'd68189,17'd68190,17'd68191,17'd68123,17'd68192,17'd68193,17'd68194,17'd68195,17'd68195,17'd68196,17'd68196,17'd68196,17'd68197,17'd68197,17'd68196,17'd68196,17'd68196,17'd68198,17'd68199,17'd68200,17'd68201,17'd68202,17'd68203,17'd68204,17'd68205,17'd68206,17'd68207,17'd68208,17'd68123,17'd68209,17'd68210,17'd68211,17'd68212,17'd68213,17'd68214,17'd0,17'd0
},
'{
17'd0,17'd0,17'd68215,17'd68216,17'd68217,17'd68218,17'd68219,17'd68220,17'd68221,17'd68222,17'd68223,17'd68224,17'd68225,17'd68226,17'd68227,17'd68227,17'd68228,17'd68226,17'd68227,17'd68228,17'd68229,17'd68230,17'd68231,17'd68232,17'd68233,17'd68234,17'd68235,17'd68236,17'd68237,17'd68238,17'd68239,17'd68240,17'd68241,17'd68242,17'd68243,17'd68244,17'd68186,17'd68245,17'd0,17'd0
},
'{
17'd0,17'd0,17'd68246,17'd68247,17'd68248,17'd68249,17'd68250,17'd68251,17'd68252,17'd68253,17'd68254,17'd68255,17'd68256,17'd68257,17'd68258,17'd68258,17'd68258,17'd68258,17'd68258,17'd68258,17'd68257,17'd68259,17'd68260,17'd68261,17'd68262,17'd68263,17'd68264,17'd68265,17'd68266,17'd68267,17'd68123,17'd68268,17'd68269,17'd68270,17'd68271,17'd68272,17'd68186,17'd68273,17'd0,17'd0
},
'{
17'd0,17'd0,17'd68274,17'd68275,17'd68276,17'd68277,17'd68278,17'd68279,17'd68280,17'd68281,17'd68282,17'd68283,17'd68284,17'd68285,17'd68285,17'd68285,17'd68285,17'd68285,17'd68285,17'd68286,17'd68285,17'd68287,17'd68288,17'd68289,17'd68290,17'd68291,17'd68292,17'd68293,17'd68294,17'd68295,17'd68296,17'd68297,17'd68298,17'd68299,17'd68300,17'd68301,17'd68302,17'd68303,17'd0,17'd0
},
'{
17'd0,17'd0,17'd68304,17'd68305,17'd68306,17'd68307,17'd68308,17'd68309,17'd68310,17'd68311,17'd68312,17'd68313,17'd68314,17'd68315,17'd68315,17'd68315,17'd68315,17'd68315,17'd68315,17'd68315,17'd68316,17'd68317,17'd68318,17'd68319,17'd68320,17'd68321,17'd68322,17'd68323,17'd68324,17'd68325,17'd68326,17'd68327,17'd68328,17'd68329,17'd68330,17'd68331,17'd68332,17'd68333,17'd0,17'd0
},
'{
17'd0,17'd0,17'd68334,17'd68335,17'd68336,17'd68123,17'd68123,17'd68337,17'd68338,17'd68339,17'd68340,17'd68341,17'd68342,17'd68343,17'd68343,17'd68343,17'd68343,17'd68343,17'd68343,17'd68343,17'd68343,17'd68344,17'd68345,17'd68346,17'd68347,17'd68348,17'd68349,17'd68350,17'd68351,17'd68352,17'd68353,17'd68340,17'd68123,17'd68354,17'd68355,17'd68356,17'd65175,17'd68357,17'd0,17'd0
},
'{
17'd0,17'd0,17'd68358,17'd68359,17'd68360,17'd68123,17'd68361,17'd68362,17'd68363,17'd68364,17'd68365,17'd68123,17'd68366,17'd68367,17'd68368,17'd68368,17'd68368,17'd68368,17'd68368,17'd68368,17'd68369,17'd68370,17'd68371,17'd68372,17'd68373,17'd68374,17'd68375,17'd68376,17'd68377,17'd68378,17'd68123,17'd68379,17'd68380,17'd68381,17'd68382,17'd68383,17'd68384,17'd68385,17'd0,17'd0
},
'{
17'd0,17'd68386,17'd68387,17'd68388,17'd68389,17'd68123,17'd68390,17'd68391,17'd68392,17'd68393,17'd68394,17'd68123,17'd68395,17'd68396,17'd68397,17'd68397,17'd68397,17'd68397,17'd68397,17'd68397,17'd68398,17'd68399,17'd68400,17'd68401,17'd68402,17'd68403,17'd68404,17'd68405,17'd68406,17'd68407,17'd68408,17'd68409,17'd68410,17'd68411,17'd68412,17'd68413,17'd68414,17'd68415,17'd0,17'd0
},
'{
17'd0,17'd68416,17'd68417,17'd68418,17'd68419,17'd68123,17'd68420,17'd68421,17'd68422,17'd68423,17'd68424,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68425,17'd68426,17'd68123,17'd68427,17'd68428,17'd68429,17'd68430,17'd68406,17'd68431,17'd68432,17'd68433,17'd0,17'd0
},
'{
17'd0,17'd68434,17'd68435,17'd68436,17'd68437,17'd68123,17'd68438,17'd68439,17'd68440,17'd68441,17'd68442,17'd68443,17'd67972,17'd68444,17'd68444,17'd68445,17'd68446,17'd68447,17'd68448,17'd68449,17'd68450,17'd68451,17'd68452,17'd68453,17'd68454,17'd68455,17'd68456,17'd68457,17'd68458,17'd68340,17'd68459,17'd68460,17'd68461,17'd68462,17'd68463,17'd68464,17'd68465,17'd68466,17'd68467,17'd68468
},
'{
17'd0,17'd68469,17'd68435,17'd68436,17'd68437,17'd68123,17'd68470,17'd68439,17'd68440,17'd68471,17'd68472,17'd68473,17'd68474,17'd68475,17'd68476,17'd68477,17'd68478,17'd68479,17'd68480,17'd68481,17'd68482,17'd68483,17'd68484,17'd68485,17'd68486,17'd68487,17'd68488,17'd68489,17'd68490,17'd68340,17'd68491,17'd68492,17'd68493,17'd68494,17'd68495,17'd68496,17'd68497,17'd68498,17'd68499,17'd68500
},
'{
17'd0,17'd68501,17'd68435,17'd68436,17'd68437,17'd68123,17'd68470,17'd68439,17'd68440,17'd68471,17'd68502,17'd68503,17'd68504,17'd68505,17'd68505,17'd68505,17'd68506,17'd68507,17'd68508,17'd68509,17'd68510,17'd68511,17'd68512,17'd68513,17'd68514,17'd68515,17'd68516,17'd68517,17'd68518,17'd68340,17'd68519,17'd68520,17'd68521,17'd68522,17'd68523,17'd68524,17'd68525,17'd63443,17'd68526,17'd68527
},
'{
17'd0,17'd68434,17'd68435,17'd68528,17'd68437,17'd68123,17'd68470,17'd68439,17'd68440,17'd68471,17'd68529,17'd68530,17'd68531,17'd68532,17'd68532,17'd68532,17'd68533,17'd68534,17'd68535,17'd68536,17'd68537,17'd68538,17'd68539,17'd68540,17'd68541,17'd68542,17'd68543,17'd68544,17'd68545,17'd68546,17'd68547,17'd68548,17'd68549,17'd68550,17'd68551,17'd68552,17'd68553,17'd68554,17'd68555,17'd68556
},
'{
17'd0,17'd68434,17'd68435,17'd68436,17'd68437,17'd68123,17'd68470,17'd68439,17'd68440,17'd68471,17'd68529,17'd68531,17'd68530,17'd68530,17'd68530,17'd68557,17'd68533,17'd68558,17'd68535,17'd68536,17'd68537,17'd68559,17'd68560,17'd68561,17'd68562,17'd68542,17'd68543,17'd68544,17'd68563,17'd68123,17'd68564,17'd68565,17'd68566,17'd68567,17'd68568,17'd68569,17'd68570,17'd68571,17'd68572,17'd68573
},
'{
17'd0,17'd68574,17'd68435,17'd68436,17'd68437,17'd68123,17'd68438,17'd68439,17'd68440,17'd68471,17'd68529,17'd68530,17'd68531,17'd68532,17'd68532,17'd68532,17'd68533,17'd68575,17'd68535,17'd68576,17'd68537,17'd68559,17'd68560,17'd68561,17'd68562,17'd68542,17'd68543,17'd68577,17'd68578,17'd68546,17'd68579,17'd68580,17'd68581,17'd68550,17'd68582,17'd68074,17'd68583,17'd68584,17'd68585,17'd68586
},
'{
17'd0,17'd68587,17'd68435,17'd68436,17'd68437,17'd68123,17'd68438,17'd68439,17'd68440,17'd68471,17'd68588,17'd68589,17'd68589,17'd68590,17'd68532,17'd68531,17'd68591,17'd68592,17'd68535,17'd68576,17'd68537,17'd68593,17'd68560,17'd68561,17'd68594,17'd68595,17'd68596,17'd68597,17'd68598,17'd68599,17'd68600,17'd68601,17'd68602,17'd68603,17'd68604,17'd68605,17'd68606,17'd68607,17'd68608,17'd68500
},
'{
17'd0,17'd68609,17'd68435,17'd68436,17'd68437,17'd68123,17'd68438,17'd68439,17'd68440,17'd68471,17'd68588,17'd68589,17'd68610,17'd68610,17'd68589,17'd68611,17'd68612,17'd68592,17'd68535,17'd68576,17'd68537,17'd68559,17'd68560,17'd68613,17'd68614,17'd68615,17'd68543,17'd68597,17'd68598,17'd68123,17'd68616,17'd68617,17'd68618,17'd68619,17'd68620,17'd68621,17'd68622,17'd68623,17'd68624,17'd68625
},
'{
17'd0,17'd68434,17'd68435,17'd68436,17'd68437,17'd68123,17'd68626,17'd68439,17'd68440,17'd68471,17'd68627,17'd68628,17'd68628,17'd68628,17'd68629,17'd68530,17'd68612,17'd68630,17'd68535,17'd68536,17'd68537,17'd68559,17'd68560,17'd68613,17'd68614,17'd68615,17'd68543,17'd68597,17'd68631,17'd68340,17'd68632,17'd68633,17'd68634,17'd68635,17'd68636,17'd68621,17'd68622,17'd68637,17'd68638,17'd0
},
'{
17'd0,17'd68639,17'd68640,17'd68436,17'd68437,17'd68123,17'd68470,17'd68439,17'd68440,17'd68471,17'd68641,17'd68532,17'd68532,17'd68532,17'd68532,17'd68530,17'd68612,17'd68630,17'd68535,17'd68536,17'd68537,17'd68559,17'd68560,17'd68561,17'd68594,17'd68615,17'd68543,17'd68597,17'd68631,17'd68164,17'd68642,17'd68643,17'd68644,17'd68645,17'd68646,17'd68074,17'd68647,17'd68648,17'd68649,17'd68650
},
'{
17'd0,17'd68651,17'd68652,17'd68653,17'd68654,17'd68123,17'd68438,17'd68439,17'd68440,17'd68471,17'd68529,17'd68530,17'd68531,17'd68532,17'd68532,17'd68531,17'd68655,17'd68575,17'd68535,17'd68536,17'd68537,17'd68656,17'd68560,17'd68561,17'd68562,17'd68542,17'd68543,17'd68657,17'd68631,17'd68658,17'd68659,17'd68660,17'd68661,17'd68662,17'd68663,17'd68664,17'd68665,17'd68666,17'd68667,17'd68668
},
'{
17'd68669,17'd68670,17'd68671,17'd68672,17'd68654,17'd68123,17'd68438,17'd68439,17'd68440,17'd68471,17'd68529,17'd68531,17'd68530,17'd68530,17'd68530,17'd68530,17'd68655,17'd68575,17'd68535,17'd68536,17'd68537,17'd68559,17'd68560,17'd68561,17'd68562,17'd68542,17'd68543,17'd68597,17'd68631,17'd68658,17'd68659,17'd68673,17'd68674,17'd68662,17'd68675,17'd68676,17'd68677,17'd68678,17'd68679,17'd68680
},
'{
17'd68681,17'd68682,17'd67847,17'd68683,17'd68654,17'd68123,17'd68470,17'd68439,17'd68440,17'd68471,17'd68529,17'd68530,17'd68531,17'd68532,17'd68532,17'd68684,17'd68685,17'd68575,17'd68535,17'd68536,17'd68537,17'd68559,17'd68560,17'd68686,17'd68687,17'd68542,17'd68543,17'd68597,17'd68598,17'd68658,17'd68688,17'd68673,17'd68674,17'd68689,17'd68690,17'd68683,17'd68691,17'd68692,17'd68693,17'd68694
},
'{
17'd68695,17'd68696,17'd68697,17'd68683,17'd68654,17'd68123,17'd68470,17'd68439,17'd68440,17'd68471,17'd68529,17'd68530,17'd68531,17'd68532,17'd68590,17'd68589,17'd68591,17'd68575,17'd68535,17'd68536,17'd68537,17'd68593,17'd68560,17'd68561,17'd68698,17'd68595,17'd68543,17'd68577,17'd68699,17'd68700,17'd68701,17'd68702,17'd68703,17'd68645,17'd68704,17'd67794,17'd68705,17'd68706,17'd68707,17'd63871
},
'{
17'd68708,17'd68709,17'd68710,17'd68683,17'd68654,17'd68123,17'd68626,17'd68439,17'd68440,17'd68471,17'd68529,17'd68530,17'd68531,17'd68610,17'd68610,17'd68589,17'd68533,17'd68575,17'd68535,17'd68576,17'd68537,17'd68559,17'd68560,17'd68561,17'd68711,17'd68615,17'd68543,17'd68597,17'd68578,17'd68123,17'd68712,17'd68713,17'd68714,17'd68715,17'd68690,17'd68019,17'd68716,17'd68717,17'd68718,17'd68719
},
'{
17'd68720,17'd68721,17'd68697,17'd68683,17'd68654,17'd68123,17'd68722,17'd68439,17'd68440,17'd68471,17'd68529,17'd68684,17'd68628,17'd68628,17'd68628,17'd68557,17'd68533,17'd68558,17'd68535,17'd68536,17'd68537,17'd68559,17'd68560,17'd68561,17'd68711,17'd68615,17'd68543,17'd68544,17'd68723,17'd68700,17'd68724,17'd68725,17'd68726,17'd68727,17'd68728,17'd67794,17'd68729,17'd68717,17'd68718,17'd68719
},
'{
17'd68730,17'd68731,17'd68697,17'd68683,17'd68654,17'd68123,17'd68470,17'd68439,17'd68440,17'd68471,17'd68529,17'd68530,17'd68531,17'd68532,17'd68532,17'd68532,17'd68533,17'd68558,17'd68535,17'd68536,17'd68537,17'd68559,17'd68560,17'd68561,17'd68711,17'd68615,17'd68543,17'd68577,17'd68578,17'd68123,17'd68732,17'd68733,17'd68714,17'd68645,17'd68728,17'd67794,17'd68729,17'd68717,17'd68718,17'd68719
},
'{
17'd68734,17'd68735,17'd68736,17'd68683,17'd68654,17'd68123,17'd68470,17'd68737,17'd68440,17'd68471,17'd68502,17'd68532,17'd68532,17'd68532,17'd68532,17'd68684,17'd68685,17'd68575,17'd68535,17'd68536,17'd68537,17'd68559,17'd68560,17'd68561,17'd68711,17'd68615,17'd68543,17'd68577,17'd68738,17'd68599,17'd68739,17'd68740,17'd68741,17'd68742,17'd68728,17'd67794,17'd67937,17'd68717,17'd68718,17'd68719
},
'{
17'd68743,17'd68744,17'd68697,17'd68683,17'd68654,17'd68123,17'd68626,17'd68439,17'd68440,17'd68471,17'd68529,17'd68530,17'd68530,17'd68530,17'd68530,17'd68530,17'd68655,17'd68575,17'd68535,17'd68536,17'd68537,17'd68559,17'd68560,17'd68613,17'd68614,17'd68615,17'd68543,17'd68544,17'd68738,17'd68546,17'd68745,17'd68740,17'd68746,17'd68727,17'd68728,17'd67794,17'd67937,17'd68717,17'd68718,17'd68719
},
'{
17'd68747,17'd68748,17'd68697,17'd68683,17'd68654,17'd68123,17'd68470,17'd68439,17'd68440,17'd68471,17'd68502,17'd68532,17'd68532,17'd68532,17'd68532,17'd68531,17'd68685,17'd68575,17'd68749,17'd68536,17'd68537,17'd68559,17'd68539,17'd68613,17'd68614,17'd68595,17'd68750,17'd68751,17'd68578,17'd68546,17'd68752,17'd68740,17'd68746,17'd68645,17'd68728,17'd67794,17'd67937,17'd68717,17'd68718,17'd68719
},
'{
17'd68753,17'd68754,17'd68710,17'd68672,17'd68755,17'd68123,17'd68756,17'd68367,17'd68757,17'd68758,17'd68759,17'd68760,17'd68760,17'd68760,17'd68760,17'd68760,17'd68761,17'd68613,17'd68762,17'd68763,17'd68764,17'd68765,17'd68766,17'd68613,17'd68614,17'd68595,17'd68543,17'd68767,17'd68578,17'd68768,17'd68769,17'd68770,17'd68771,17'd68772,17'd68773,17'd67794,17'd67937,17'd68717,17'd68718,17'd68719
},
'{
17'd68774,17'd68775,17'd68697,17'd68683,17'd68776,17'd68123,17'd68777,17'd68778,17'd68779,17'd68780,17'd68781,17'd68782,17'd68782,17'd68782,17'd68782,17'd68628,17'd68505,17'd68783,17'd68784,17'd68785,17'd68786,17'd68787,17'd68788,17'd68789,17'd68711,17'd68595,17'd68790,17'd68791,17'd68792,17'd68123,17'd68793,17'd68794,17'd68123,17'd68795,17'd68796,17'd67764,17'd67937,17'd68717,17'd68718,17'd68719
},
'{
17'd68797,17'd68798,17'd68697,17'd68683,17'd68799,17'd68800,17'd68801,17'd68802,17'd68803,17'd68804,17'd68805,17'd68806,17'd68806,17'd68806,17'd68806,17'd68807,17'd68808,17'd68809,17'd68810,17'd68811,17'd68812,17'd68813,17'd68814,17'd68815,17'd68711,17'd68816,17'd68817,17'd68818,17'd68819,17'd68820,17'd68821,17'd68822,17'd68823,17'd68824,17'd68825,17'd67794,17'd67937,17'd68717,17'd68718,17'd68719
},
'{
17'd68826,17'd68827,17'd68736,17'd67794,17'd67731,17'd68828,17'd68829,17'd68830,17'd68831,17'd68832,17'd68833,17'd68834,17'd68834,17'd68834,17'd68834,17'd68835,17'd68835,17'd68834,17'd68836,17'd68837,17'd68838,17'd68839,17'd68840,17'd68841,17'd68842,17'd68843,17'd68844,17'd68845,17'd67873,17'd68846,17'd68847,17'd68848,17'd68849,17'd68850,17'd68851,17'd67794,17'd67937,17'd68717,17'd68718,17'd68719
},
'{
17'd68852,17'd68853,17'd67875,17'd67794,17'd67794,17'd68854,17'd68855,17'd67794,17'd67795,17'd67795,17'd67766,17'd67794,17'd67794,17'd67794,17'd67794,17'd67795,17'd67766,17'd67795,17'd68856,17'd67921,17'd67851,17'd67876,17'd68857,17'd67878,17'd67901,17'd68858,17'd67987,17'd68859,17'd67795,17'd67795,17'd67766,17'd67875,17'd68860,17'd68861,17'd67874,17'd67794,17'd68716,17'd68717,17'd68718,17'd68719
},
'{
17'd68862,17'd68863,17'd68697,17'd67794,17'd67794,17'd68864,17'd67794,17'd67794,17'd67794,17'd67794,17'd67794,17'd67794,17'd67794,17'd67794,17'd67794,17'd67794,17'd67764,17'd67795,17'd67849,17'd67921,17'd67851,17'd67876,17'd67877,17'd67900,17'd67901,17'd67880,17'd67987,17'd68859,17'd67794,17'd67794,17'd67794,17'd67875,17'd68860,17'd68865,17'd67874,17'd67794,17'd68716,17'd68717,17'd68718,17'd68719
},
'{
17'd68866,17'd68867,17'd68736,17'd67794,17'd67794,17'd68864,17'd67848,17'd67794,17'd67794,17'd67794,17'd67875,17'd67875,17'd67875,17'd67875,17'd67875,17'd67875,17'd67875,17'd68697,17'd67849,17'd67921,17'd68868,17'd68869,17'd68870,17'd68871,17'd68872,17'd68873,17'd68874,17'd68875,17'd67874,17'd67794,17'd67794,17'd67875,17'd68860,17'd68865,17'd67874,17'd67794,17'd67937,17'd68717,17'd68718,17'd68719
},
'{
17'd68876,17'd68877,17'd68697,17'd67794,17'd67794,17'd68864,17'd67848,17'd67794,17'd67794,17'd68878,17'd67956,17'd68016,17'd68016,17'd68016,17'd68016,17'd68016,17'd67956,17'd68879,17'd68880,17'd68881,17'd68882,17'd68883,17'd68884,17'd68885,17'd68886,17'd68887,17'd68888,17'd68889,17'd68865,17'd67874,17'd67794,17'd67875,17'd68860,17'd68865,17'd67874,17'd67794,17'd67937,17'd68717,17'd68718,17'd68719
},
'{
17'd68890,17'd68891,17'd68697,17'd67794,17'd67794,17'd68864,17'd67848,17'd67794,17'd67794,17'd67955,17'd68023,17'd67971,17'd67971,17'd67971,17'd67971,17'd67971,17'd67971,17'd68023,17'd68880,17'd68892,17'd68893,17'd68894,17'd68895,17'd68896,17'd68897,17'd68898,17'd68899,17'd68900,17'd68901,17'd67875,17'd67794,17'd67875,17'd68860,17'd68865,17'd67874,17'd67794,17'd67937,17'd68717,17'd68718,17'd68719
},
'{
17'd68902,17'd68903,17'd68710,17'd67794,17'd67848,17'd68864,17'd67848,17'd67794,17'd67794,17'd67794,17'd67937,17'd67938,17'd67937,17'd67938,17'd67938,17'd67937,17'd67938,17'd67937,17'd68904,17'd68905,17'd68906,17'd68907,17'd68908,17'd68909,17'd68910,17'd68911,17'd68912,17'd67795,17'd67874,17'd67794,17'd67794,17'd67875,17'd68860,17'd68865,17'd67874,17'd67794,17'd67937,17'd68717,17'd68718,17'd68719
},
'{
17'd68913,17'd68914,17'd68697,17'd67794,17'd67848,17'd68864,17'd67848,17'd67794,17'd67848,17'd67794,17'd67848,17'd68879,17'd68016,17'd68016,17'd68016,17'd68016,17'd68016,17'd67956,17'd68915,17'd68881,17'd68916,17'd68917,17'd68918,17'd68919,17'd68920,17'd68921,17'd68922,17'd67897,17'd67874,17'd67794,17'd67794,17'd67875,17'd68860,17'd68865,17'd67874,17'd67794,17'd67937,17'd68717,17'd68718,17'd68719
},
'{
17'd68923,17'd68924,17'd68697,17'd67794,17'd67848,17'd68925,17'd67848,17'd67794,17'd67848,17'd67794,17'd68926,17'd68023,17'd67971,17'd67971,17'd67971,17'd67971,17'd67971,17'd67971,17'd68927,17'd68928,17'd68929,17'd68930,17'd68931,17'd68932,17'd68933,17'd68934,17'd68935,17'd68936,17'd67874,17'd67794,17'd67794,17'd67875,17'd68860,17'd68865,17'd67874,17'd67794,17'd67937,17'd68717,17'd68718,17'd68719
},
'{
17'd68937,17'd68938,17'd68736,17'd67794,17'd67848,17'd68925,17'd67848,17'd67794,17'd67848,17'd67794,17'd67794,17'd67874,17'd67937,17'd67937,17'd67937,17'd67937,17'd67937,17'd67937,17'd68939,17'd68940,17'd68941,17'd68942,17'd68943,17'd68944,17'd68945,17'd68946,17'd68947,17'd68948,17'd67794,17'd67794,17'd67794,17'd67875,17'd68860,17'd68865,17'd67874,17'd67794,17'd67937,17'd68717,17'd68718,17'd68719
},
'{
17'd68949,17'd68950,17'd67875,17'd67794,17'd67848,17'd68864,17'd67794,17'd67794,17'd67794,17'd67794,17'd67848,17'd67875,17'd68016,17'd67918,17'd67918,17'd67918,17'd67918,17'd67918,17'd68915,17'd68951,17'd68952,17'd68052,17'd68953,17'd68954,17'd68955,17'd68956,17'd68957,17'd68958,17'd67794,17'd67794,17'd67794,17'd67875,17'd68860,17'd68865,17'd67874,17'd67794,17'd67937,17'd68717,17'd68718,17'd68719
},
'{
17'd68959,17'd68960,17'd68710,17'd67794,17'd67794,17'd68864,17'd67794,17'd67794,17'd67794,17'd67794,17'd67794,17'd67874,17'd68900,17'd68900,17'd68900,17'd68900,17'd68900,17'd68925,17'd68915,17'd68961,17'd68962,17'd68963,17'd68964,17'd68965,17'd68966,17'd68967,17'd68968,17'd67794,17'd67794,17'd67794,17'd67794,17'd67875,17'd68860,17'd68865,17'd67874,17'd67794,17'd67937,17'd68717,17'd68718,17'd68719
},
'{
17'd68969,17'd68970,17'd68697,17'd67794,17'd67794,17'd68864,17'd67794,17'd67794,17'd67794,17'd67794,17'd67848,17'd67874,17'd67874,17'd67875,17'd67875,17'd67875,17'd67875,17'd67875,17'd68904,17'd68905,17'd68971,17'd68972,17'd68973,17'd68974,17'd68975,17'd68976,17'd68977,17'd68859,17'd67794,17'd67794,17'd67794,17'd67875,17'd68860,17'd68865,17'd67874,17'd67794,17'd67937,17'd68717,17'd68718,17'd68719
},
'{
17'd68978,17'd68979,17'd68736,17'd67794,17'd67794,17'd68864,17'd67794,17'd67794,17'd67794,17'd67794,17'd67794,17'd67848,17'd67874,17'd68980,17'd68980,17'd68980,17'd68980,17'd68936,17'd68880,17'd68981,17'd68982,17'd68983,17'd68984,17'd68985,17'd68986,17'd68987,17'd68021,17'd68859,17'd67794,17'd67794,17'd67794,17'd67875,17'd68860,17'd68980,17'd67874,17'd67794,17'd67937,17'd68717,17'd68718,17'd68719
},
'{
17'd68988,17'd68989,17'd68697,17'd67794,17'd67794,17'd68864,17'd67794,17'd67794,17'd67794,17'd67794,17'd67794,17'd67848,17'd67875,17'd67920,17'd68925,17'd68925,17'd68925,17'd68925,17'd68880,17'd68990,17'd68991,17'd68992,17'd68993,17'd68994,17'd68995,17'd68996,17'd68021,17'd68859,17'd67794,17'd67794,17'd67794,17'd67875,17'd68860,17'd68980,17'd67874,17'd67794,17'd68997,17'd68717,17'd68718,17'd68719
},
'{
17'd68998,17'd68999,17'd68697,17'd67794,17'd67794,17'd68864,17'd67848,17'd67794,17'd67848,17'd67794,17'd67794,17'd67794,17'd67848,17'd67794,17'd67794,17'd67874,17'd67794,17'd67874,17'd68856,17'd67921,17'd69000,17'd69001,17'd69002,17'd69003,17'd69004,17'd69005,17'd69006,17'd68859,17'd67794,17'd67794,17'd67794,17'd67875,17'd68860,17'd68865,17'd68710,17'd69007,17'd68691,17'd69008,17'd68718,17'd68719
},
'{
17'd69009,17'd69010,17'd68697,17'd67794,17'd67794,17'd68925,17'd67794,17'd67794,17'd67794,17'd67794,17'd67794,17'd67794,17'd67848,17'd68926,17'd67794,17'd67794,17'd67794,17'd67794,17'd67849,17'd67921,17'd67851,17'd69011,17'd69012,17'd69013,17'd69014,17'd69015,17'd69016,17'd68859,17'd67794,17'd67794,17'd67794,17'd67875,17'd69017,17'd68980,17'd68710,17'd69007,17'd69018,17'd69019,17'd68718,17'd68719
},
'{
17'd69020,17'd69021,17'd69022,17'd69023,17'd69024,17'd69025,17'd69026,17'd69027,17'd69026,17'd69027,17'd69026,17'd69027,17'd69026,17'd69027,17'd69027,17'd69027,17'd69026,17'd69026,17'd69028,17'd69029,17'd69030,17'd69031,17'd69032,17'd69033,17'd68911,17'd69034,17'd69035,17'd68697,17'd69027,17'd69026,17'd69027,17'd69022,17'd69036,17'd69037,17'd68418,17'd68773,17'd69038,17'd69039,17'd68718,17'd68719
},
'{
17'd69040,17'd69041,17'd69042,17'd69043,17'd69044,17'd69045,17'd69046,17'd69047,17'd69048,17'd69049,17'd69050,17'd69051,17'd69052,17'd69053,17'd69054,17'd69054,17'd69054,17'd69055,17'd69056,17'd69057,17'd69058,17'd69059,17'd69060,17'd69061,17'd69062,17'd69063,17'd69064,17'd69065,17'd69066,17'd69067,17'd69068,17'd69069,17'd69070,17'd69041,17'd69071,17'd69072,17'd69073,17'd69074,17'd69075,17'd69076
},
'{
17'd69077,17'd69078,17'd69079,17'd69080,17'd69081,17'd69082,17'd69083,17'd69084,17'd69085,17'd69086,17'd69087,17'd69088,17'd69089,17'd69090,17'd69091,17'd69091,17'd69091,17'd69091,17'd69092,17'd69093,17'd69094,17'd69081,17'd69091,17'd69091,17'd69095,17'd69090,17'd69096,17'd69097,17'd69098,17'd69099,17'd69100,17'd69101,17'd69102,17'd69103,17'd69104,17'd69105,17'd69106,17'd69107,17'd69108,17'd69109
},
'{
17'd69110,17'd69111,17'd69112,17'd69113,17'd69114,17'd69115,17'd69112,17'd69116,17'd69117,17'd69118,17'd69119,17'd69120,17'd69121,17'd69122,17'd69123,17'd69124,17'd69122,17'd69122,17'd69122,17'd69122,17'd69122,17'd69123,17'd69124,17'd69122,17'd69122,17'd69125,17'd69126,17'd69127,17'd69118,17'd69128,17'd69129,17'd69130,17'd69131,17'd69132,17'd69133,17'd69115,17'd69134,17'd69135,17'd69136,17'd69137
},
'{
17'd0,17'd69138,17'd69139,17'd69140,17'd69141,17'd69142,17'd69143,17'd69144,17'd69145,17'd69146,17'd69147,17'd69148,17'd69149,17'd69150,17'd69151,17'd69152,17'd69153,17'd69153,17'd69153,17'd69153,17'd69153,17'd69151,17'd69150,17'd69153,17'd69153,17'd69150,17'd69154,17'd69155,17'd69156,17'd69157,17'd69158,17'd69159,17'd69160,17'd69161,17'd69162,17'd69163,17'd69164,17'd69165,17'd69166,17'd0
},
'{
17'd0,17'd69167,17'd69168,17'd69169,17'd69170,17'd69171,17'd69172,17'd69173,17'd68727,17'd68645,17'd68742,17'd69174,17'd69175,17'd69176,17'd69177,17'd69174,17'd69176,17'd69176,17'd69176,17'd69176,17'd69176,17'd69177,17'd69176,17'd69176,17'd69176,17'd69176,17'd69176,17'd69178,17'd69179,17'd68727,17'd69180,17'd69179,17'd68715,17'd69181,17'd69182,17'd69183,17'd69184,17'd69185,17'd69186,17'd0
},
'{
17'd0,17'd0,17'd0,17'd0,17'd69187,17'd69188,17'd69189,17'd69190,17'd69191,17'd51874,17'd51874,17'd51874,17'd51874,17'd51874,17'd48280,17'd69191,17'd51874,17'd51874,17'd51874,17'd51874,17'd69191,17'd48280,17'd51874,17'd51874,17'd51874,17'd51874,17'd51874,17'd69191,17'd48280,17'd51874,17'd69191,17'd69191,17'd51874,17'd51874,17'd69192,17'd69193,17'd69194,17'd69195,17'd0,17'd0
},
'{
17'd0,17'd0,17'd0,17'd0,17'd0,17'd49700,17'd69196,17'd864,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69197,17'd69198,17'd69199,17'd69200,17'd0,17'd0,17'd0
}};
endmodule
