module images/basicbackground(output logic [3:0] rgb[0:639][0:479]);
assign rgb = '{
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd1,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
},
'{
3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4
}};
endmodule
