module basicbackground(output logic [5:0] rgb[0:639][0:479]);
assign rgb = '{
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd15,5'd15,5'd15,5'd15,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
}};
endmodule
