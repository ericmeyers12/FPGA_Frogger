module images/frog3(output logic [17:0] rgb[0:39][0:39]);
assign rgb = '{
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd70854,17'd68123,17'd71295,17'd71304,17'd71305,17'd71306,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd71307,17'd68123,17'd71308,17'd71309,17'd71310,17'd71311,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd71312,17'd71312,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd71313,17'd68123,17'd70857,17'd71177,17'd71245,17'd71274,17'd71314,17'd71308,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71312,17'd71312,17'd70856,17'd68123,17'd68123,17'd71315,17'd71316,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd71312,17'd71312,17'd70862,17'd71306,17'd71317,17'd71312,17'd71296,17'd71318,17'd71319,17'd71320,17'd70893,17'd71226,17'd70946,17'd71225,17'd71321,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd71322,17'd71323,17'd71324,17'd71325,17'd71312,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd71312,17'd68123,17'd71326,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd71327,17'd68123,17'd71133,17'd71328,17'd71329,17'd71330,17'd70946,17'd71331,17'd71332,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71333,17'd71334,17'd71308,17'd71335,17'd71116,17'd71336,17'd68123,17'd71305,17'd71305,17'd71312,17'd71312,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd71337,17'd71338,17'd71339,17'd71340,17'd71341,17'd71342,17'd71343,17'd71344,17'd71312,17'd71345,17'd71329,17'd71346,17'd71347,17'd71348,17'd71349,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71350,17'd71351,17'd70988,17'd71352,17'd71353,17'd71354,17'd71355,17'd68123,17'd68123,17'd71356,17'd71357,17'd71358,17'd71359,17'd68123,17'd68123,17'd68123,17'd68123,17'd71360,17'd71310,17'd49131,17'd71361,17'd71362,17'd71363,17'd71364,17'd71365,17'd71366,17'd71367,17'd71368,17'd39023,17'd71329,17'd71369,17'd71370,17'd71371,17'd71372,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71373,17'd71374,17'd71375,17'd71376,17'd70923,17'd70905,17'd71377,17'd71378,17'd71379,17'd71380,17'd71381,17'd68123,17'd71382,17'd71383,17'd68123,17'd68123,17'd68123,17'd71384,17'd71385,17'd71386,17'd71190,17'd71039,17'd71189,17'd71387,17'd71388,17'd71389,17'd71390,17'd71391,17'd71392,17'd71329,17'd71393,17'd71310,17'd68340,17'd71394,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71395,17'd71396,17'd71397,17'd71398,17'd70905,17'd70923,17'd70906,17'd71399,17'd71400,17'd71401,17'd71402,17'd71403,17'd71404,17'd71405,17'd71312,17'd68123,17'd68123,17'd71406,17'd71407,17'd71408,17'd71409,17'd71410,17'd71411,17'd71412,17'd71413,17'd70922,17'd71414,17'd71415,17'd71416,17'd71417,17'd70877,17'd68123,17'd71418,17'd71419,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71308,17'd71420,17'd71198,17'd70884,17'd71189,17'd71258,17'd70988,17'd71421,17'd71410,17'd71422,17'd71423,17'd71424,17'd71425,17'd68123,17'd70856,17'd71426,17'd71426,17'd23693,17'd71427,17'd71428,17'd46938,17'd71429,17'd71261,17'd71430,17'd71431,17'd71432,17'd71433,17'd71320,17'd71434,17'd71433,17'd71395,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71435,17'd71436,17'd71437,17'd71438,17'd71264,17'd71439,17'd71440,17'd71441,17'd71334,17'd71323,17'd71442,17'd71443,17'd64125,17'd71444,17'd68123,17'd68123,17'd68123,17'd71445,17'd71446,17'd71447,17'd71448,17'd71449,17'd71281,17'd70872,17'd68123,17'd68123,17'd71307,17'd71283,17'd71450,17'd71252,17'd70862,17'd71313,17'd71312,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71306,17'd71451,17'd70872,17'd71318,17'd71452,17'd71453,17'd71454,17'd71455,17'd71456,17'd71333,17'd71457,17'd71458,17'd65027,17'd32726,17'd71459,17'd71460,17'd30322,17'd71461,17'd71462,17'd71463,17'd71464,17'd71465,17'd71219,17'd71411,17'd71466,17'd68123,17'd70862,17'd71426,17'd71467,17'd71468,17'd71283,17'd70854,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd71469,17'd71470,17'd71471,17'd71472,17'd71473,17'd71474,17'd71198,17'd71475,17'd11240,17'd71476,17'd71477,17'd71478,17'd71479,17'd71480,17'd71481,17'd71482,17'd71483,17'd71484,17'd71485,17'd24995,17'd71486,17'd71487,17'd71488,17'd68123,17'd70856,17'd71312,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd71312,17'd71489,17'd71490,17'd71491,17'd71492,17'd71008,17'd70922,17'd71493,17'd71011,17'd71494,17'd71013,17'd71476,17'd71495,17'd71496,17'd71017,17'd71497,17'd71019,17'd71020,17'd71021,17'd71498,17'd71499,17'd71500,17'd71025,17'd71501,17'd71502,17'd68123,17'd71503,17'd71312,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd71312,17'd71504,17'd71505,17'd71506,17'd71507,17'd71508,17'd71509,17'd71036,17'd71037,17'd71510,17'd29466,17'd71039,17'd71040,17'd64726,17'd71042,17'd70978,17'd71511,17'd66641,17'd71074,17'd51878,17'd70955,17'd71512,17'd71513,17'd71514,17'd71515,17'd71516,17'd68123,17'd70856,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd71312,17'd68123,17'd71517,17'd71055,17'd71056,17'd71518,17'd71519,17'd71520,17'd71038,17'd71240,17'd71062,17'd71037,17'd71062,17'd71062,17'd71063,17'd70887,17'd70887,17'd70887,17'd71062,17'd71063,17'd71037,17'd71062,17'd71062,17'd71064,17'd71521,17'd71522,17'd71523,17'd71177,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd71312,17'd68123,17'd71524,17'd71525,17'd71526,17'd61244,17'd66236,17'd71527,17'd71528,17'd71071,17'd71072,17'd20462,17'd71079,17'd71074,17'd70966,17'd71076,17'd38459,17'd70966,17'd71529,17'd66641,17'd71044,17'd71080,17'd71080,17'd71080,17'd71081,17'd71166,17'd71438,17'd71530,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd71312,17'd68123,17'd71531,17'd71086,17'd71532,17'd70887,17'd70887,17'd71088,17'd71059,17'd71089,17'd71533,17'd71059,17'd71090,17'd71534,17'd71088,17'd71061,17'd70887,17'd70887,17'd71092,17'd71091,17'd70906,17'd70906,17'd71092,17'd71039,17'd71094,17'd71535,17'd71536,17'd71537,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd71312,17'd71538,17'd71539,17'd71540,17'd71101,17'd71102,17'd71541,17'd70954,17'd71037,17'd71037,17'd71104,17'd70887,17'd71062,17'd70954,17'd38114,17'd71542,17'd71543,17'd71544,17'd71106,17'd71089,17'd24523,17'd71545,17'd12099,17'd71109,17'd71546,17'd71547,17'd71548,17'd71549,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd71550,17'd71551,17'd71552,17'd71009,17'd71117,17'd71062,17'd71118,17'd71553,17'd71554,17'd71041,17'd71555,17'd71122,17'd71123,17'd71556,17'd71124,17'd71557,17'd71127,17'd71128,17'd71558,17'd71559,17'd71560,17'd71561,17'd71562,17'd68123,17'd70856,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd71312,17'd71563,17'd71564,17'd71565,17'd71566,17'd64822,17'd70952,17'd71567,17'd71568,17'd71569,17'd71570,17'd71571,17'd71572,17'd71146,17'd71573,17'd71148,17'd71574,17'd71575,17'd71576,17'd61648,17'd71577,17'd71578,17'd7684,17'd71579,17'd71548,17'd68123,17'd71312,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd71580,17'd68123,17'd71581,17'd71582,17'd71583,17'd71584,17'd71585,17'd71586,17'd70966,17'd70886,17'd71587,17'd71588,17'd71589,17'd71590,17'd29063,17'd13563,17'd71591,17'd71592,17'd71593,17'd71594,17'd70974,17'd71595,17'd71225,17'd68123,17'd70841,17'd71312,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71432,17'd71596,17'd71597,17'd71598,17'd71451,17'd71599,17'd68123,17'd68123,17'd71600,17'd71601,17'd71602,17'd71223,17'd70921,17'd71395,17'd71603,17'd71604,17'd71605,17'd71606,17'd71607,17'd70898,17'd71608,17'd21423,17'd71609,17'd70924,17'd71530,17'd68123,17'd71317,17'd71310,17'd71610,17'd71195,17'd71611,17'd71612,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71613,17'd70894,17'd71614,17'd71530,17'd70988,17'd71615,17'd56026,17'd71616,17'd71617,17'd71618,17'd71529,17'd71267,17'd71619,17'd68123,17'd71620,17'd71621,17'd71622,17'd71308,17'd68123,17'd71623,17'd71624,17'd9785,17'd71413,17'd71439,17'd71306,17'd68123,17'd71625,17'd71598,17'd71626,17'd71627,17'd71628,17'd71629,17'd71312,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71245,17'd71412,17'd71188,17'd71410,17'd70905,17'd71630,17'd54826,17'd71631,17'd71632,17'd71633,17'd71634,17'd71635,17'd68123,17'd70862,17'd71306,17'd68123,17'd68123,17'd71450,17'd71636,17'd71637,17'd71638,17'd71639,17'd71264,17'd71330,17'd71640,17'd71641,17'd71642,17'd71320,17'd70884,17'd71643,17'd71371,17'd68123,17'd71312,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71644,17'd71645,17'd71646,17'd70868,17'd70887,17'd71092,17'd71647,17'd71648,17'd71649,17'd71650,17'd71651,17'd71652,17'd71426,17'd71450,17'd68123,17'd68123,17'd68123,17'd71653,17'd71603,17'd71654,17'd71655,17'd71116,17'd71375,17'd71266,17'd71219,17'd71656,17'd71657,17'd71658,17'd42322,17'd71659,17'd71660,17'd68123,17'd70856,17'd70862,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71661,17'd71266,17'd70922,17'd71662,17'd71260,17'd70922,17'd71335,17'd71663,17'd71664,17'd71165,17'd71604,17'd68123,17'd70854,17'd68123,17'd68123,17'd68123,17'd68123,17'd71665,17'd71452,17'd71666,17'd71667,17'd71668,17'd71669,17'd71670,17'd71089,17'd71671,17'd71672,17'd71673,17'd42930,17'd71674,17'd71675,17'd71598,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71627,17'd71676,17'd71374,17'd71393,17'd70886,17'd71677,17'd71313,17'd71678,17'd71679,17'd68123,17'd70854,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd71426,17'd71305,17'd71680,17'd71681,17'd71682,17'd71683,17'd71684,17'd71685,17'd71686,17'd71687,17'd71688,17'd71689,17'd71659,17'd71369,17'd71675,17'd70872,17'd71690,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71337,17'd71466,17'd71691,17'd70931,17'd70888,17'd71350,17'd68123,17'd68123,17'd70854,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68340,17'd71307,17'd71692,17'd33280,17'd24864,17'd41917,17'd12413,17'd71693,17'd71694,17'd68123,17'd71695,17'd71696,17'd71697,17'd71347,17'd71432,17'd71698,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd70881,17'd71010,17'd71438,17'd70963,17'd71699,17'd70861,17'd71699,17'd71312,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd71312,17'd68123,17'd70854,17'd68123,17'd68123,17'd68123,17'd71312,17'd68123,17'd19885,17'd68123,17'd71610,17'd71643,17'd71659,17'd71330,17'd71700,17'd71701,17'd71702,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd71373,17'd71315,17'd71626,17'd71648,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd71312,17'd71312,17'd71269,17'd71269,17'd70832,17'd71305,17'd71269,17'd71305,17'd71703,17'd71433,17'd70921,17'd71226,17'd71467,17'd71225,17'd71704,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd71312,17'd68123,17'd70846,17'd70946,17'd71705,17'd71706,17'd70842,17'd71395,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd71312,17'd68123,17'd71707,17'd71663,17'd71708,17'd71691,17'd68123,17'd70856,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd70854,17'd68123,17'd71679,17'd70846,17'd71305,17'd71306,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
}};
endmodule
