module images/numbers(output logic [5:0] rgb[0:239][0:31]);
assign rgb = '{
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd0,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
},
'{
5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14
}};
endmodule
