module lilypad_sprite(output logic [5:0] rgb[0:39][0:39]);
assign rgb = '{
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
}};
endmodule
