nprince@wirelessprvnat-172-17-101-143.near.illinois.edu.14458