module testimage(output logic [17:0] rgb[0:639][0:479]);
assign rgb = '{
'{
17'd0,17'd0,17'd0,17'd0,17'd0,17'd0,17'd0,17'd0,17'd1,17'd1,17'd1,17'd0,17'd2,17'd2,17'd0,17'd3,17'd4,17'd5,17'd6,17'd6,17'd7,17'd6,17'd8,17'd4,17'd9,17'd9,17'd10,17'd11,17'd12,17'd13,17'd2,17'd2,17'd14,17'd14,17'd14,17'd14,17'd15,17'd15,17'd16,17'd17,17'd17,17'd17,17'd17,17'd16,17'd18,17'd18,17'd19,17'd19,17'd18,17'd18,17'd11,17'd11,17'd11,17'd11,17'd20,17'd20,17'd21,17'd21,17'd22,17'd23,17'd23,17'd23,17'd24,17'd24,17'd22,17'd22,17'd23,17'd23,17'd25,17'd25,17'd21,17'd21,17'd26,17'd26,17'd27,17'd27,17'd28,17'd29,17'd30,17'd31,17'd32,17'd33,17'd34,17'd34,17'd35,17'd36,17'd37,17'd38,17'd39,17'd39,17'd39,17'd40,17'd40,17'd40,17'd40,17'd41,17'd42,17'd43,17'd44,17'd44,17'd45,17'd45,17'd46,17'd46,17'd47,17'd48,17'd49,17'd50,17'd51,17'd52,17'd53,17'd54,17'd55,17'd55,17'd56,17'd57,17'd57,17'd57,17'd58,17'd59,17'd60,17'd60,17'd61,17'd61,17'd62,17'd62,17'd63,17'd64,17'd65,17'd66,17'd67,17'd68,17'd69,17'd70,17'd70,17'd69,17'd71,17'd71,17'd72,17'd72,17'd73,17'd73,17'd74,17'd75,17'd76,17'd77,17'd78,17'd79,17'd80,17'd81,17'd82,17'd83,17'd84,17'd85,17'd86,17'd86,17'd86,17'd86,17'd87,17'd88,17'd89,17'd90,17'd91,17'd92,17'd93,17'd94,17'd95,17'd96,17'd97,17'd98,17'd99,17'd100,17'd101,17'd102,17'd103,17'd104,17'd105,17'd106,17'd107,17'd108,17'd109,17'd110,17'd111,17'd112,17'd113,17'd114,17'd115,17'd116,17'd117,17'd118,17'd119,17'd120,17'd121,17'd122,17'd123,17'd124,17'd125,17'd125,17'd126,17'd127,17'd128,17'd128,17'd129,17'd130,17'd130,17'd130,17'd130,17'd130,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd132,17'd134,17'd135,17'd132,17'd131,17'd131,17'd131,17'd130,17'd136,17'd137,17'd138,17'd139,17'd140,17'd141,17'd141,17'd140,17'd142,17'd143,17'd144,17'd145,17'd146,17'd147,17'd148,17'd149,17'd150,17'd151,17'd152,17'd153,17'd154,17'd155,17'd156,17'd157,17'd158,17'd159,17'd160,17'd161,17'd162,17'd163,17'd164,17'd165,17'd166,17'd167,17'd168,17'd169,17'd170,17'd170,17'd169,17'd169,17'd171,17'd172,17'd173,17'd174,17'd175,17'd176,17'd177,17'd178,17'd179,17'd180,17'd181,17'd182,17'd183,17'd184,17'd185,17'd186,17'd187,17'd188,17'd189,17'd190,17'd191,17'd192,17'd193,17'd194,17'd195,17'd195,17'd196,17'd197,17'd198,17'd199,17'd200,17'd201,17'd202,17'd203,17'd204,17'd205,17'd206,17'd206,17'd207,17'd207,17'd208,17'd209,17'd210,17'd211,17'd212,17'd213,17'd214,17'd215,17'd177,17'd216,17'd217,17'd218,17'd219,17'd220,17'd221,17'd222,17'd223,17'd224,17'd225,17'd226,17'd227,17'd228,17'd229,17'd230,17'd231,17'd232,17'd233,17'd233,17'd234,17'd235,17'd236,17'd237,17'd238,17'd239,17'd240,17'd241,17'd241,17'd239,17'd238,17'd242,17'd242,17'd242,17'd242,17'd243,17'd244,17'd245,17'd246,17'd247,17'd248,17'd249,17'd250,17'd251,17'd251,17'd251,17'd180,17'd252,17'd253,17'd253,17'd254,17'd255,17'd256,17'd257,17'd258,17'd258,17'd259,17'd260,17'd258,17'd261,17'd262,17'd256,17'd263,17'd264,17'd265,17'd266,17'd264,17'd267,17'd268,17'd262,17'd262,17'd257,17'd269,17'd270,17'd271,17'd271,17'd272,17'd272,17'd273,17'd274,17'd275,17'd276,17'd277,17'd278,17'd279,17'd280,17'd281,17'd282
},
'{
17'd0,17'd0,17'd0,17'd0,17'd0,17'd0,17'd0,17'd0,17'd1,17'd1,17'd1,17'd0,17'd2,17'd2,17'd1,17'd283,17'd4,17'd5,17'd6,17'd6,17'd6,17'd6,17'd8,17'd4,17'd9,17'd25,17'd10,17'd19,17'd12,17'd13,17'd2,17'd2,17'd14,17'd14,17'd14,17'd14,17'd14,17'd14,17'd17,17'd17,17'd16,17'd16,17'd16,17'd16,17'd18,17'd18,17'd18,17'd18,17'd18,17'd18,17'd11,17'd11,17'd11,17'd11,17'd20,17'd21,17'd21,17'd21,17'd22,17'd23,17'd23,17'd23,17'd284,17'd284,17'd23,17'd23,17'd23,17'd23,17'd25,17'd25,17'd21,17'd21,17'd285,17'd285,17'd286,17'd287,17'd288,17'd289,17'd290,17'd291,17'd292,17'd293,17'd34,17'd294,17'd36,17'd295,17'd37,17'd38,17'd39,17'd39,17'd296,17'd296,17'd39,17'd40,17'd40,17'd297,17'd43,17'd43,17'd44,17'd298,17'd45,17'd45,17'd46,17'd46,17'd299,17'd300,17'd50,17'd51,17'd51,17'd301,17'd301,17'd302,17'd56,17'd56,17'd57,17'd57,17'd57,17'd57,17'd58,17'd59,17'd303,17'd303,17'd61,17'd61,17'd62,17'd62,17'd63,17'd64,17'd304,17'd305,17'd305,17'd68,17'd69,17'd69,17'd69,17'd69,17'd306,17'd307,17'd308,17'd309,17'd310,17'd73,17'd311,17'd312,17'd77,17'd78,17'd313,17'd314,17'd80,17'd315,17'd82,17'd83,17'd316,17'd317,17'd86,17'd318,17'd318,17'd318,17'd319,17'd320,17'd321,17'd322,17'd323,17'd324,17'd325,17'd326,17'd95,17'd96,17'd327,17'd328,17'd329,17'd330,17'd331,17'd332,17'd333,17'd334,17'd335,17'd336,17'd337,17'd338,17'd339,17'd340,17'd341,17'd342,17'd343,17'd344,17'd345,17'd346,17'd347,17'd348,17'd349,17'd350,17'd351,17'd352,17'd353,17'd354,17'd355,17'd355,17'd127,17'd356,17'd128,17'd134,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd132,17'd134,17'd135,17'd135,17'd357,17'd357,17'd357,17'd358,17'd140,17'd359,17'd360,17'd360,17'd361,17'd361,17'd362,17'd363,17'd143,17'd364,17'd365,17'd366,17'd367,17'd368,17'd369,17'd370,17'd371,17'd372,17'd373,17'd374,17'd375,17'd154,17'd376,17'd377,17'd378,17'd379,17'd380,17'd381,17'd382,17'd383,17'd384,17'd385,17'd386,17'd387,17'd388,17'd388,17'd389,17'd390,17'd391,17'd392,17'd393,17'd394,17'd395,17'd396,17'd397,17'd398,17'd177,17'd399,17'd400,17'd401,17'd402,17'd182,17'd403,17'd404,17'd405,17'd406,17'd407,17'd408,17'd409,17'd410,17'd411,17'd412,17'd413,17'd414,17'd415,17'd416,17'd417,17'd418,17'd417,17'd196,17'd419,17'd420,17'd421,17'd422,17'd423,17'd424,17'd425,17'd206,17'd426,17'd426,17'd427,17'd427,17'd428,17'd429,17'd430,17'd431,17'd432,17'd433,17'd434,17'd435,17'd436,17'd437,17'd438,17'd219,17'd221,17'd439,17'd440,17'd441,17'd442,17'd226,17'd443,17'd444,17'd230,17'd445,17'd446,17'd446,17'd443,17'd428,17'd447,17'd448,17'd235,17'd235,17'd236,17'd238,17'd239,17'd449,17'd240,17'd449,17'd450,17'd243,17'd451,17'd451,17'd451,17'd242,17'd244,17'd245,17'd452,17'd453,17'd454,17'd455,17'd251,17'd251,17'd251,17'd213,17'd180,17'd252,17'd253,17'd253,17'd456,17'd255,17'd256,17'd256,17'd261,17'd258,17'd426,17'd260,17'd271,17'd207,17'd256,17'd262,17'd257,17'd457,17'd266,17'd266,17'd263,17'd264,17'd268,17'd257,17'd256,17'd257,17'd269,17'd269,17'd271,17'd271,17'd270,17'd272,17'd273,17'd273,17'd458,17'd275,17'd459,17'd460,17'd461,17'd462,17'd463,17'd464
},
'{
17'd0,17'd0,17'd0,17'd0,17'd0,17'd0,17'd15,17'd15,17'd1,17'd0,17'd0,17'd2,17'd13,17'd12,17'd283,17'd465,17'd8,17'd6,17'd6,17'd6,17'd6,17'd6,17'd4,17'd4,17'd9,17'd25,17'd10,17'd19,17'd12,17'd2,17'd2,17'd466,17'd14,17'd14,17'd14,17'd14,17'd14,17'd14,17'd17,17'd17,17'd16,17'd16,17'd18,17'd18,17'd18,17'd18,17'd18,17'd18,17'd11,17'd11,17'd11,17'd11,17'd11,17'd10,17'd21,17'd21,17'd25,17'd25,17'd23,17'd23,17'd22,17'd22,17'd22,17'd22,17'd24,17'd24,17'd23,17'd23,17'd25,17'd25,17'd25,17'd21,17'd467,17'd467,17'd286,17'd28,17'd29,17'd468,17'd290,17'd469,17'd470,17'd293,17'd33,17'd471,17'd295,17'd472,17'd473,17'd473,17'd38,17'd38,17'd474,17'd474,17'd475,17'd41,17'd297,17'd476,17'd477,17'd44,17'd44,17'd298,17'd45,17'd45,17'd478,17'd478,17'd479,17'd479,17'd51,17'd301,17'd301,17'd302,17'd302,17'd302,17'd57,17'd57,17'd57,17'd57,17'd57,17'd57,17'd480,17'd480,17'd481,17'd482,17'd62,17'd483,17'd483,17'd483,17'd63,17'd64,17'd64,17'd484,17'd484,17'd485,17'd486,17'd486,17'd487,17'd487,17'd487,17'd488,17'd489,17'd489,17'd490,17'd73,17'd491,17'd492,17'd493,17'd494,17'd495,17'd496,17'd80,17'd315,17'd497,17'd498,17'd499,17'd500,17'd318,17'd501,17'd501,17'd501,17'd502,17'd503,17'd504,17'd505,17'd506,17'd507,17'd508,17'd509,17'd510,17'd511,17'd512,17'd513,17'd514,17'd515,17'd516,17'd517,17'd518,17'd519,17'd520,17'd521,17'd522,17'd523,17'd524,17'd525,17'd526,17'd527,17'd528,17'd529,17'd530,17'd531,17'd532,17'd533,17'd534,17'd535,17'd536,17'd537,17'd538,17'd539,17'd540,17'd540,17'd541,17'd542,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd130,17'd130,17'd128,17'd128,17'd358,17'd358,17'd543,17'd544,17'd545,17'd362,17'd546,17'd143,17'd143,17'd547,17'd548,17'd549,17'd550,17'd365,17'd551,17'd552,17'd553,17'd554,17'd555,17'd556,17'd557,17'd558,17'd559,17'd560,17'd561,17'd562,17'd563,17'd564,17'd565,17'd566,17'd567,17'd568,17'd569,17'd570,17'd571,17'd572,17'd573,17'd574,17'd575,17'd576,17'd577,17'd578,17'd579,17'd580,17'd581,17'd582,17'd583,17'd584,17'd585,17'd586,17'd587,17'd588,17'd589,17'd590,17'd591,17'd592,17'd593,17'd430,17'd594,17'd594,17'd595,17'd596,17'd597,17'd426,17'd191,17'd192,17'd598,17'd415,17'd198,17'd197,17'd417,17'd599,17'd599,17'd418,17'd417,17'd600,17'd194,17'd601,17'd602,17'd603,17'd604,17'd605,17'd606,17'd206,17'd260,17'd260,17'd607,17'd608,17'd609,17'd610,17'd611,17'd612,17'd613,17'd614,17'd434,17'd615,17'd616,17'd617,17'd618,17'd619,17'd620,17'd455,17'd621,17'd622,17'd428,17'd623,17'd227,17'd446,17'd624,17'd625,17'd626,17'd627,17'd447,17'd447,17'd628,17'd629,17'd630,17'd630,17'd630,17'd237,17'd631,17'd632,17'd631,17'd237,17'd451,17'd451,17'd451,17'd451,17'd622,17'd633,17'd245,17'd634,17'd635,17'd636,17'd637,17'd637,17'd213,17'd638,17'd639,17'd182,17'd181,17'd253,17'd456,17'd460,17'd255,17'd255,17'd256,17'd257,17'd640,17'd270,17'd641,17'd642,17'd207,17'd257,17'd257,17'd268,17'd268,17'd257,17'd256,17'd262,17'd257,17'd268,17'd257,17'd256,17'd261,17'd258,17'd207,17'd271,17'd271,17'd642,17'd643,17'd644,17'd645,17'd273,17'd646,17'd255,17'd253,17'd647,17'd648,17'd649
},
'{
17'd0,17'd0,17'd0,17'd0,17'd0,17'd0,17'd15,17'd15,17'd0,17'd0,17'd2,17'd2,17'd13,17'd12,17'd650,17'd651,17'd8,17'd6,17'd6,17'd6,17'd6,17'd4,17'd4,17'd25,17'd25,17'd10,17'd19,17'd18,17'd2,17'd2,17'd2,17'd2,17'd14,17'd14,17'd14,17'd14,17'd14,17'd14,17'd17,17'd17,17'd16,17'd16,17'd18,17'd18,17'd18,17'd18,17'd19,17'd19,17'd11,17'd11,17'd11,17'd11,17'd10,17'd10,17'd25,17'd25,17'd25,17'd25,17'd23,17'd22,17'd22,17'd22,17'd22,17'd22,17'd24,17'd24,17'd23,17'd23,17'd25,17'd25,17'd25,17'd25,17'd467,17'd286,17'd652,17'd653,17'd468,17'd30,17'd654,17'd655,17'd470,17'd33,17'd656,17'd657,17'd658,17'd472,17'd659,17'd659,17'd660,17'd660,17'd474,17'd474,17'd475,17'd41,17'd297,17'd661,17'd477,17'd44,17'd44,17'd298,17'd45,17'd45,17'd478,17'd662,17'd479,17'd663,17'd301,17'd302,17'd54,17'd54,17'd664,17'd665,17'd666,17'd666,17'd666,17'd57,17'd57,17'd57,17'd667,17'd667,17'd481,17'd482,17'd62,17'd483,17'd483,17'd483,17'd63,17'd668,17'd668,17'd668,17'd484,17'd669,17'd670,17'd670,17'd488,17'd488,17'd671,17'd672,17'd489,17'd308,17'd73,17'd673,17'd491,17'd674,17'd313,17'd314,17'd314,17'd80,17'd675,17'd315,17'd498,17'd676,17'd677,17'd678,17'd679,17'd680,17'd681,17'd681,17'd682,17'd683,17'd684,17'd685,17'd686,17'd687,17'd687,17'd687,17'd688,17'd689,17'd690,17'd691,17'd692,17'd693,17'd694,17'd695,17'd696,17'd697,17'd698,17'd699,17'd700,17'd701,17'd702,17'd703,17'd704,17'd705,17'd706,17'd707,17'd708,17'd709,17'd710,17'd711,17'd712,17'd713,17'd714,17'd715,17'd716,17'd717,17'd718,17'd719,17'd542,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd720,17'd721,17'd722,17'd722,17'd723,17'd724,17'd725,17'd726,17'd727,17'd728,17'd729,17'd730,17'd729,17'd731,17'd732,17'd733,17'd734,17'd367,17'd367,17'd735,17'd736,17'd737,17'd737,17'd738,17'd739,17'd740,17'd741,17'd742,17'd743,17'd371,17'd744,17'd745,17'd746,17'd747,17'd748,17'd749,17'd750,17'd751,17'd752,17'd753,17'd754,17'd755,17'd756,17'd757,17'd758,17'd759,17'd760,17'd761,17'd762,17'd763,17'd764,17'd765,17'd766,17'd767,17'd768,17'd769,17'd770,17'd591,17'd592,17'd611,17'd430,17'd442,17'd594,17'd771,17'd188,17'd772,17'd258,17'd773,17'd774,17'd775,17'd193,17'd414,17'd776,17'd197,17'd196,17'd417,17'd418,17'd418,17'd418,17'd418,17'd777,17'd778,17'd779,17'd780,17'd602,17'd192,17'd781,17'd605,17'd260,17'd260,17'd427,17'd607,17'd782,17'd783,17'd234,17'd622,17'd784,17'd454,17'd785,17'd786,17'd787,17'd788,17'd436,17'd789,17'd790,17'd791,17'd454,17'd792,17'd793,17'd794,17'd626,17'd231,17'd625,17'd625,17'd625,17'd626,17'd795,17'd447,17'd447,17'd628,17'd796,17'd448,17'd448,17'd630,17'd237,17'd797,17'd797,17'd797,17'd243,17'd242,17'd798,17'd798,17'd799,17'd622,17'd244,17'd633,17'd800,17'd621,17'd636,17'd432,17'd638,17'd638,17'd639,17'd182,17'd182,17'd181,17'd254,17'd456,17'd255,17'd801,17'd256,17'd257,17'd269,17'd270,17'd642,17'd641,17'd641,17'd642,17'd268,17'd257,17'd646,17'd268,17'd262,17'd802,17'd262,17'd257,17'd257,17'd262,17'd261,17'd258,17'd207,17'd271,17'd642,17'd259,17'd644,17'd644,17'd803,17'd644,17'd273,17'd262,17'd804,17'd805,17'd279,17'd612
},
'{
17'd12,17'd12,17'd0,17'd0,17'd15,17'd15,17'd15,17'd15,17'd15,17'd14,17'd2,17'd2,17'd12,17'd806,17'd651,17'd807,17'd8,17'd6,17'd6,17'd6,17'd4,17'd4,17'd23,17'd25,17'd20,17'd11,17'd12,17'd12,17'd2,17'd2,17'd14,17'd14,17'd14,17'd14,17'd14,17'd14,17'd14,17'd14,17'd17,17'd17,17'd16,17'd16,17'd18,17'd18,17'd18,17'd19,17'd19,17'd19,17'd11,17'd11,17'd11,17'd10,17'd10,17'd808,17'd25,17'd25,17'd21,17'd21,17'd22,17'd22,17'd23,17'd23,17'd23,17'd23,17'd24,17'd24,17'd23,17'd23,17'd25,17'd25,17'd808,17'd808,17'd27,17'd27,17'd652,17'd653,17'd289,17'd809,17'd654,17'd655,17'd32,17'd656,17'd657,17'd810,17'd658,17'd811,17'd36,17'd812,17'd813,17'd814,17'd296,17'd296,17'd41,17'd815,17'd816,17'd816,17'd817,17'd663,17'd818,17'd819,17'd819,17'd818,17'd818,17'd663,17'd301,17'd302,17'd302,17'd820,17'd820,17'd821,17'd822,17'd823,17'd824,17'd824,17'd825,17'd825,17'd826,17'd826,17'd667,17'd827,17'd828,17'd829,17'd830,17'd830,17'd831,17'd831,17'd832,17'd832,17'd833,17'd834,17'd835,17'd835,17'd836,17'd836,17'd837,17'd837,17'd672,17'd488,17'd838,17'd839,17'd840,17'd841,17'd842,17'd843,17'd844,17'd845,17'd846,17'd80,17'd847,17'd675,17'd848,17'd849,17'd850,17'd851,17'd852,17'd853,17'd854,17'd855,17'd855,17'd856,17'd857,17'd858,17'd859,17'd859,17'd860,17'd861,17'd862,17'd863,17'd864,17'd865,17'd866,17'd867,17'd868,17'd869,17'd870,17'd871,17'd872,17'd873,17'd874,17'd875,17'd876,17'd877,17'd878,17'd879,17'd880,17'd881,17'd882,17'd883,17'd884,17'd885,17'd886,17'd887,17'd715,17'd718,17'd718,17'd888,17'd888,17'd889,17'd542,17'd133,17'd133,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd130,17'd130,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd130,17'd130,17'd128,17'd720,17'd721,17'd890,17'd363,17'd891,17'd892,17'd893,17'd894,17'd895,17'd896,17'd897,17'd898,17'd898,17'd898,17'd899,17'd900,17'd901,17'd902,17'd903,17'd904,17'd905,17'd906,17'd907,17'd908,17'd909,17'd910,17'd911,17'd912,17'd913,17'd914,17'd915,17'd916,17'd917,17'd918,17'd919,17'd920,17'd921,17'd922,17'd923,17'd756,17'd924,17'd925,17'd926,17'd927,17'd928,17'd929,17'd930,17'd930,17'd455,17'd455,17'd931,17'd932,17'd932,17'd933,17'd181,17'd934,17'd405,17'd610,17'd188,17'd608,17'd935,17'd641,17'd458,17'd645,17'd936,17'd937,17'd938,17'd939,17'd940,17'd941,17'd942,17'd943,17'd944,17'd945,17'd945,17'd599,17'd946,17'd947,17'd948,17'd949,17'd950,17'd951,17'd598,17'd952,17'd605,17'd644,17'd259,17'd259,17'd953,17'd954,17'd443,17'd782,17'd234,17'd244,17'd955,17'd956,17'd614,17'd434,17'd615,17'd957,17'd464,17'd958,17'd249,17'd635,17'd634,17'd622,17'd782,17'd626,17'd227,17'd446,17'd625,17'd625,17'd446,17'd443,17'd232,17'd447,17'd447,17'd447,17'd959,17'd959,17'd796,17'd960,17'd236,17'd797,17'd797,17'd236,17'd235,17'd448,17'd234,17'd793,17'd961,17'd244,17'd784,17'd962,17'd621,17'd635,17'd592,17'd592,17'd963,17'd964,17'd182,17'd182,17'd965,17'd804,17'd456,17'd966,17'd967,17'd263,17'd968,17'd968,17'd272,17'd273,17'd274,17'd274,17'd272,17'd269,17'd271,17'd271,17'd257,17'd802,17'd969,17'd459,17'd266,17'd459,17'd262,17'd256,17'd207,17'd271,17'd259,17'd970,17'd803,17'd605,17'd971,17'd972,17'd973,17'd640,17'd974,17'd967,17'd975,17'd976
},
'{
17'd12,17'd12,17'd0,17'd0,17'd15,17'd15,17'd15,17'd15,17'd14,17'd14,17'd2,17'd12,17'd806,17'd465,17'd977,17'd978,17'd6,17'd6,17'd6,17'd4,17'd4,17'd25,17'd25,17'd10,17'd11,17'd19,17'd12,17'd2,17'd2,17'd2,17'd14,17'd14,17'd14,17'd14,17'd14,17'd14,17'd14,17'd14,17'd17,17'd17,17'd16,17'd16,17'd18,17'd18,17'd18,17'd19,17'd19,17'd979,17'd11,17'd11,17'd10,17'd10,17'd808,17'd808,17'd25,17'd25,17'd25,17'd25,17'd23,17'd23,17'd23,17'd23,17'd23,17'd23,17'd24,17'd24,17'd23,17'd23,17'd25,17'd25,17'd808,17'd10,17'd980,17'd652,17'd28,17'd288,17'd981,17'd31,17'd982,17'd32,17'd983,17'd984,17'd984,17'd657,17'd811,17'd471,17'd35,17'd35,17'd985,17'd986,17'd296,17'd41,17'd815,17'd815,17'd815,17'd987,17'd663,17'd663,17'd818,17'd818,17'd818,17'd663,17'd663,17'd988,17'd54,17'd665,17'd665,17'd821,17'd822,17'd989,17'd990,17'd990,17'd991,17'd824,17'd824,17'd824,17'd992,17'd992,17'd827,17'd827,17'd828,17'd829,17'd993,17'd830,17'd994,17'd994,17'd995,17'd996,17'd997,17'd997,17'd998,17'd998,17'd836,17'd999,17'd837,17'd837,17'd307,17'd307,17'd1000,17'd839,17'd840,17'd842,17'd843,17'd1001,17'd1002,17'd845,17'd846,17'd1003,17'd1004,17'd1005,17'd1006,17'd1007,17'd1008,17'd1009,17'd1010,17'd1011,17'd1012,17'd1013,17'd1014,17'd1015,17'd1016,17'd1017,17'd1018,17'd1019,17'd1020,17'd1021,17'd1022,17'd1023,17'd1024,17'd1025,17'd1026,17'd1027,17'd1028,17'd1029,17'd1030,17'd1031,17'd1032,17'd1033,17'd1034,17'd1035,17'd1036,17'd1037,17'd1038,17'd1039,17'd1040,17'd1041,17'd1042,17'd711,17'd712,17'd885,17'd1043,17'd715,17'd1044,17'd718,17'd718,17'd889,17'd889,17'd1045,17'd1045,17'd1045,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd130,17'd130,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd128,17'd720,17'd720,17'd721,17'd721,17'd1046,17'd1047,17'd1048,17'd892,17'd1049,17'd1050,17'd1051,17'd1052,17'd1053,17'd1054,17'd1055,17'd1056,17'd1057,17'd1057,17'd1058,17'd1059,17'd1060,17'd1061,17'd1062,17'd1063,17'd1064,17'd1065,17'd1066,17'd1067,17'd1068,17'd1069,17'd1070,17'd1071,17'd1072,17'd1073,17'd1074,17'd1075,17'd1076,17'd1077,17'd1078,17'd1079,17'd1080,17'd1081,17'd1082,17'd1083,17'd1084,17'd1085,17'd1086,17'd1087,17'd1088,17'd1089,17'd1090,17'd1091,17'd1092,17'd1093,17'd1094,17'd1095,17'd404,17'd1096,17'd801,17'd408,17'd1097,17'd209,17'd207,17'd642,17'd644,17'd803,17'd1098,17'd1099,17'd598,17'd1100,17'd1101,17'd1102,17'd1103,17'd1104,17'd943,17'd944,17'd945,17'd1105,17'd945,17'd1106,17'd1106,17'd1107,17'd1108,17'd1109,17'd1110,17'd780,17'd602,17'd191,17'd1111,17'd425,17'd1112,17'd1112,17'd1113,17'd1113,17'd231,17'd1114,17'd959,17'd799,17'd1115,17'd455,17'd614,17'd1116,17'd786,17'd1117,17'd1117,17'd1118,17'd249,17'd963,17'd593,17'd429,17'd794,17'd623,17'd446,17'd228,17'd1119,17'd228,17'd446,17'd227,17'd443,17'd795,17'd447,17'd959,17'd447,17'd1120,17'd628,17'd1121,17'd236,17'd237,17'd237,17'd630,17'd448,17'd1122,17'd1122,17'd793,17'd961,17'd242,17'd784,17'd800,17'd962,17'd963,17'd592,17'd963,17'd964,17'd182,17'd182,17'd1123,17'd965,17'd804,17'd456,17'd801,17'd967,17'd256,17'd968,17'd273,17'd274,17'd273,17'd273,17'd273,17'd273,17'd271,17'd271,17'd207,17'd256,17'd265,17'd265,17'd265,17'd265,17'd262,17'd256,17'd207,17'd271,17'd259,17'd970,17'd605,17'd781,17'd424,17'd204,17'd1098,17'd1124,17'd1125,17'd257,17'd1126,17'd460
},
'{
17'd12,17'd12,17'd1,17'd1,17'd15,17'd15,17'd15,17'd14,17'd1127,17'd14,17'd0,17'd3,17'd465,17'd977,17'd978,17'd978,17'd6,17'd6,17'd4,17'd4,17'd23,17'd25,17'd21,17'd10,17'd10,17'd19,17'd12,17'd2,17'd2,17'd14,17'd14,17'd14,17'd1127,17'd1127,17'd1127,17'd14,17'd17,17'd17,17'd16,17'd16,17'd16,17'd16,17'd18,17'd18,17'd18,17'd19,17'd19,17'd19,17'd1128,17'd11,17'd10,17'd808,17'd25,17'd25,17'd25,17'd21,17'd25,17'd25,17'd25,17'd25,17'd23,17'd23,17'd23,17'd23,17'd24,17'd24,17'd4,17'd4,17'd25,17'd10,17'd27,17'd27,17'd652,17'd652,17'd652,17'd29,17'd809,17'd1129,17'd982,17'd1130,17'd983,17'd1130,17'd656,17'd656,17'd656,17'd656,17'd294,17'd35,17'd659,17'd986,17'd39,17'd40,17'd1131,17'd1132,17'd987,17'd987,17'd663,17'd663,17'd663,17'd663,17'd302,17'd54,17'd54,17'd665,17'd1133,17'd822,17'd822,17'd990,17'd990,17'd1134,17'd1135,17'd1135,17'd1136,17'd1137,17'd1138,17'd1138,17'd1139,17'd1139,17'd1140,17'd1140,17'd1141,17'd1142,17'd1143,17'd1143,17'd1144,17'd1144,17'd1144,17'd1145,17'd1146,17'd1147,17'd998,17'd998,17'd836,17'd1148,17'd670,17'd487,17'd70,17'd70,17'd839,17'd1149,17'd1150,17'd1151,17'd1152,17'd1152,17'd844,17'd845,17'd1153,17'd1153,17'd1154,17'd1155,17'd1156,17'd1157,17'd1158,17'd1159,17'd1160,17'd1161,17'd1162,17'd1163,17'd1164,17'd1165,17'd1166,17'd1167,17'd1168,17'd1169,17'd1170,17'd1171,17'd1172,17'd1173,17'd1174,17'd1175,17'd1176,17'd1177,17'd1178,17'd1179,17'd1180,17'd1181,17'd1182,17'd1183,17'd1184,17'd1185,17'd1186,17'd1187,17'd1188,17'd1189,17'd1190,17'd709,17'd1191,17'd1192,17'd1193,17'd1194,17'd537,17'd713,17'd715,17'd1195,17'd1196,17'd1196,17'd541,17'd1197,17'd1197,17'd134,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd129,17'd141,17'd141,17'd141,17'd140,17'd1198,17'd545,17'd1199,17'd1200,17'd1201,17'd1202,17'd1203,17'd1204,17'd904,17'd1205,17'd1206,17'd1207,17'd1208,17'd1209,17'd1210,17'd1211,17'd1212,17'd1213,17'd1211,17'd1214,17'd1215,17'd1216,17'd1217,17'd1218,17'd1219,17'd1220,17'd1221,17'd1222,17'd1223,17'd1224,17'd1225,17'd1226,17'd1227,17'd1228,17'd1229,17'd1230,17'd1231,17'd1232,17'd922,17'd1233,17'd1234,17'd1235,17'd1236,17'd1237,17'd1238,17'd1089,17'd225,17'd1239,17'd1240,17'd607,17'd1241,17'd801,17'd1242,17'd641,17'd1243,17'd643,17'd206,17'd644,17'd803,17'd971,17'd971,17'd1244,17'd1245,17'd1246,17'd602,17'd414,17'd1247,17'd1103,17'd199,17'd197,17'd944,17'd945,17'd945,17'd1105,17'd1248,17'd1249,17'd1250,17'd1251,17'd1252,17'd1108,17'd948,17'd1110,17'd1253,17'd603,17'd424,17'd775,17'd1254,17'd1255,17'd1255,17'd1256,17'd953,17'd233,17'd429,17'd1257,17'd442,17'd964,17'd251,17'd249,17'd433,17'd1258,17'd1259,17'd214,17'd213,17'd462,17'd1092,17'd1122,17'd623,17'd446,17'd1260,17'd228,17'd1261,17'd1262,17'd1263,17'd954,17'd443,17'd443,17'd795,17'd795,17'd795,17'd795,17'd1264,17'd959,17'd960,17'd1265,17'd1265,17'd960,17'd234,17'd1122,17'd234,17'd793,17'd451,17'd242,17'd238,17'd1115,17'd212,17'd453,17'd212,17'd634,17'd181,17'd181,17'd181,17'd182,17'd1123,17'd965,17'd456,17'd1126,17'd1266,17'd1267,17'd1268,17'd1269,17'd273,17'd273,17'd803,17'd645,17'd644,17'd272,17'd270,17'd968,17'd266,17'd265,17'd1270,17'd1271,17'd459,17'd266,17'd257,17'd268,17'd271,17'd970,17'd605,17'd781,17'd424,17'd204,17'd1272,17'd971,17'd1273,17'd968,17'd266,17'd1274
},
'{
17'd12,17'd3,17'd1,17'd1,17'd15,17'd15,17'd14,17'd14,17'd1127,17'd2,17'd12,17'd1275,17'd977,17'd807,17'd978,17'd978,17'd6,17'd6,17'd4,17'd4,17'd25,17'd10,17'd10,17'd979,17'd979,17'd1276,17'd1,17'd0,17'd14,17'd1127,17'd1127,17'd1127,17'd1127,17'd1127,17'd1127,17'd1127,17'd17,17'd16,17'd16,17'd16,17'd1277,17'd16,17'd18,17'd18,17'd18,17'd18,17'd19,17'd19,17'd1128,17'd11,17'd10,17'd808,17'd25,17'd25,17'd21,17'd21,17'd9,17'd9,17'd25,17'd25,17'd23,17'd23,17'd23,17'd23,17'd24,17'd23,17'd4,17'd9,17'd808,17'd10,17'd980,17'd1278,17'd28,17'd652,17'd289,17'd30,17'd1129,17'd982,17'd292,17'd292,17'd1130,17'd32,17'd293,17'd293,17'd293,17'd33,17'd294,17'd36,17'd473,17'd1279,17'd40,17'd40,17'd41,17'd1132,17'd1280,17'd987,17'd817,17'd663,17'd663,17'd817,17'd54,17'd820,17'd665,17'd821,17'd823,17'd990,17'd990,17'd1281,17'd1281,17'd1282,17'd1283,17'd1283,17'd1136,17'd1136,17'd1284,17'd1138,17'd1285,17'd1139,17'd1140,17'd1286,17'd1141,17'd1141,17'd1287,17'd1287,17'd1288,17'd1288,17'd1288,17'd1144,17'd1146,17'd1289,17'd998,17'd1290,17'd1148,17'd488,17'd487,17'd307,17'd1291,17'd1000,17'd1149,17'd841,17'd1151,17'd1292,17'd1292,17'd1293,17'd1002,17'd1002,17'd1294,17'd1294,17'd1295,17'd1296,17'd1297,17'd1298,17'd1299,17'd1299,17'd1300,17'd1301,17'd1302,17'd1303,17'd1304,17'd1167,17'd1305,17'd1306,17'd1307,17'd1308,17'd1309,17'd1310,17'd1311,17'd1312,17'd1313,17'd1314,17'd1315,17'd1316,17'd1317,17'd1318,17'd1319,17'd1320,17'd1321,17'd1322,17'd1323,17'd1324,17'd1325,17'd1326,17'd1327,17'd1328,17'd1329,17'd1330,17'd1331,17'd1332,17'd1333,17'd1334,17'd1335,17'd1336,17'd538,17'd1195,17'd1195,17'd1196,17'd541,17'd356,17'd1197,17'd1197,17'd1197,17'd134,17'd130,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd130,17'd136,17'd136,17'd136,17'd136,17'd1337,17'd1338,17'd1339,17'd1340,17'd1201,17'd1341,17'd1342,17'd1343,17'd1344,17'd1345,17'd1346,17'd1347,17'd1348,17'd1349,17'd1213,17'd1350,17'd1351,17'd1352,17'd1353,17'd1353,17'd1354,17'd1355,17'd1356,17'd1357,17'd1358,17'd1359,17'd1360,17'd1361,17'd1362,17'd1363,17'd1364,17'd1365,17'd1366,17'd1367,17'd1368,17'd1369,17'd1370,17'd1371,17'd1372,17'd1373,17'd1374,17'd1375,17'd1234,17'd1376,17'd1377,17'd1378,17'd1379,17'd783,17'd953,17'd1380,17'd409,17'd641,17'd260,17'd643,17'd605,17'd424,17'd1272,17'd1381,17'd1381,17'd1244,17'd1381,17'd1382,17'd422,17'd1246,17'd1383,17'd779,17'd941,17'd941,17'd198,17'd198,17'd942,17'd944,17'd945,17'd1105,17'd1384,17'd1385,17'd1386,17'd1387,17'd1388,17'd1389,17'd1390,17'd1391,17'd1392,17'd1393,17'd1099,17'd1272,17'd1394,17'd1254,17'd1395,17'd1396,17'd427,17'd953,17'd794,17'd609,17'd622,17'd244,17'd634,17'd592,17'd432,17'd1397,17'd214,17'd1398,17'd589,17'd638,17'd431,17'd799,17'd627,17'd227,17'd1399,17'd1400,17'd1401,17'd1401,17'd1263,17'd1263,17'd443,17'd443,17'd1402,17'd1402,17'd795,17'd795,17'd795,17'd795,17'd628,17'd1121,17'd1265,17'd1265,17'd793,17'd1122,17'd1122,17'd234,17'd448,17'd451,17'd242,17'd238,17'd452,17'd453,17'd212,17'd593,17'd253,17'd461,17'd461,17'd182,17'd1403,17'd1404,17'd804,17'd966,17'd263,17'd1405,17'd1406,17'd1407,17'd273,17'd458,17'd645,17'd803,17'd803,17'd644,17'd272,17'd272,17'd268,17'd459,17'd969,17'd1270,17'd265,17'd459,17'd266,17'd268,17'd646,17'd259,17'd605,17'd781,17'd423,17'd1408,17'd603,17'd1409,17'd1410,17'd1411,17'd1407,17'd257
},
'{
17'd0,17'd1,17'd1412,17'd1,17'd15,17'd1127,17'd1127,17'd14,17'd0,17'd1,17'd283,17'd651,17'd1413,17'd8,17'd6,17'd6,17'd4,17'd4,17'd4,17'd23,17'd21,17'd10,17'd1275,17'd283,17'd283,17'd1,17'd2,17'd1127,17'd1127,17'd1127,17'd1127,17'd1127,17'd1414,17'd1415,17'd1415,17'd1414,17'd1416,17'd16,17'd16,17'd17,17'd18,17'd18,17'd18,17'd19,17'd19,17'd18,17'd18,17'd18,17'd808,17'd808,17'd808,17'd808,17'd25,17'd25,17'd25,17'd25,17'd25,17'd25,17'd25,17'd25,17'd23,17'd23,17'd23,17'd4,17'd23,17'd4,17'd23,17'd21,17'd1128,17'd1128,17'd28,17'd287,17'd652,17'd653,17'd468,17'd468,17'd290,17'd291,17'd982,17'd32,17'd470,17'd292,17'd292,17'd32,17'd33,17'd656,17'd811,17'd811,17'd1417,17'd1418,17'd38,17'd474,17'd475,17'd41,17'd815,17'd816,17'd1419,17'd1420,17'd820,17'd820,17'd665,17'd822,17'd823,17'd990,17'd1421,17'd1281,17'd1135,17'd1283,17'd1283,17'd1422,17'd1423,17'd1283,17'd1424,17'd1424,17'd1424,17'd1424,17'd1285,17'd1285,17'd1425,17'd1426,17'd1427,17'd1427,17'd1428,17'd1428,17'd1288,17'd1288,17'd1144,17'd1144,17'd998,17'd998,17'd998,17'd836,17'd837,17'd487,17'd307,17'd1000,17'd839,17'd1149,17'd1429,17'd1150,17'd1430,17'd1292,17'd843,17'd78,17'd494,17'd1431,17'd1432,17'd1433,17'd1434,17'd1435,17'd1436,17'd1437,17'd1438,17'd1439,17'd1440,17'd1441,17'd1442,17'd1443,17'd1305,17'd1444,17'd1445,17'd1446,17'd1447,17'd1448,17'd1449,17'd1450,17'd1451,17'd1452,17'd1453,17'd1454,17'd1455,17'd1456,17'd1457,17'd1458,17'd1459,17'd1460,17'd1461,17'd1322,17'd1462,17'd1463,17'd1464,17'd1465,17'd1466,17'd1467,17'd1468,17'd1469,17'd1470,17'd1471,17'd1472,17'd1473,17'd1474,17'd1475,17'd536,17'd1476,17'd1477,17'd1478,17'd1478,17'd1479,17'd1196,17'd1196,17'd1480,17'd1481,17'd133,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd358,17'd543,17'd358,17'd1482,17'd1483,17'd363,17'd546,17'd143,17'd366,17'd365,17'd551,17'd552,17'd1484,17'd1485,17'd1343,17'd1486,17'd1487,17'd1488,17'd561,17'd1489,17'd1490,17'd1491,17'd1492,17'd1493,17'd1494,17'd1495,17'd1496,17'd1497,17'd1498,17'd1499,17'd1500,17'd1501,17'd1502,17'd1503,17'd1504,17'd1505,17'd1506,17'd1507,17'd1508,17'd1509,17'd1510,17'd1511,17'd1512,17'd1513,17'd1514,17'd1515,17'd1516,17'd1517,17'd1518,17'd1519,17'd1520,17'd1521,17'd1522,17'd1523,17'd1524,17'd800,17'd793,17'd607,17'd410,17'd645,17'd1111,17'd1394,17'd1525,17'd203,17'd1526,17'd420,17'd1527,17'd1528,17'd1528,17'd420,17'd1529,17'd415,17'd415,17'd415,17'd194,17'd778,17'd417,17'd196,17'd197,17'd196,17'd1530,17'd1531,17'd1532,17'd1533,17'd1251,17'd1534,17'd1534,17'd1534,17'd1535,17'd1535,17'd1536,17'd949,17'd780,17'd602,17'd952,17'd1537,17'd1538,17'd425,17'd259,17'd259,17'd607,17'd1539,17'd783,17'd783,17'd210,17'd1540,17'd635,17'd637,17'd1541,17'd613,17'd1542,17'd1543,17'd612,17'd430,17'd609,17'd443,17'd1260,17'd228,17'd1401,17'd1401,17'd1263,17'd1262,17'd625,17'd227,17'd1544,17'd227,17'd446,17'd227,17'd795,17'd795,17'd1402,17'd795,17'd959,17'd1545,17'd1545,17'd1546,17'd447,17'd226,17'd448,17'd448,17'd793,17'd622,17'd633,17'd1540,17'd453,17'd1547,17'd593,17'd611,17'd253,17'd461,17'd253,17'd402,17'd1548,17'd804,17'd459,17'd263,17'd968,17'd968,17'd270,17'd274,17'd803,17'd644,17'd645,17'd803,17'd273,17'd272,17'd935,17'd264,17'd459,17'd969,17'd1270,17'd1126,17'd1274,17'd265,17'd646,17'd641,17'd644,17'd605,17'd1272,17'd1272,17'd1381,17'd1549,17'd1550,17'd1551,17'd1273,17'd1552
},
'{
17'd1,17'd1,17'd1412,17'd1,17'd14,17'd1127,17'd14,17'd14,17'd1,17'd283,17'd465,17'd977,17'd8,17'd8,17'd6,17'd6,17'd4,17'd4,17'd23,17'd25,17'd10,17'd10,17'd283,17'd1412,17'd1412,17'd15,17'd14,17'd1127,17'd1127,17'd1127,17'd1127,17'd1127,17'd1414,17'd1415,17'd1415,17'd1415,17'd17,17'd16,17'd16,17'd16,17'd18,17'd18,17'd18,17'd18,17'd19,17'd19,17'd19,17'd19,17'd10,17'd10,17'd10,17'd10,17'd21,17'd21,17'd21,17'd21,17'd25,17'd25,17'd25,17'd25,17'd23,17'd23,17'd23,17'd23,17'd4,17'd23,17'd21,17'd20,17'd10,17'd10,17'd28,17'd652,17'd652,17'd653,17'd468,17'd290,17'd1129,17'd1129,17'd982,17'd292,17'd292,17'd470,17'd470,17'd292,17'd33,17'd984,17'd811,17'd472,17'd1553,17'd37,17'd660,17'd296,17'd41,17'd1131,17'd816,17'd1419,17'd1554,17'd1555,17'd821,17'd821,17'd822,17'd990,17'd990,17'd1281,17'd1556,17'd1557,17'd1283,17'd1558,17'd1422,17'd1422,17'd1423,17'd1559,17'd1424,17'd1424,17'd1424,17'd1424,17'd1285,17'd1285,17'd1560,17'd1425,17'd1561,17'd1427,17'd1428,17'd1428,17'd1288,17'd1144,17'd1144,17'd1144,17'd998,17'd998,17'd836,17'd837,17'd488,17'd487,17'd1000,17'd839,17'd1149,17'd840,17'd841,17'd842,17'd843,17'd843,17'd1562,17'd77,17'd1563,17'd1564,17'd1565,17'd1566,17'd1567,17'd1568,17'd1569,17'd1570,17'd1571,17'd1572,17'd1573,17'd1574,17'd1575,17'd1576,17'd1577,17'd1578,17'd1579,17'd1580,17'd1581,17'd1582,17'd1583,17'd1584,17'd1585,17'd1586,17'd1587,17'd1588,17'd1589,17'd1590,17'd1591,17'd1592,17'd1593,17'd1594,17'd1595,17'd1596,17'd1597,17'd1598,17'd1599,17'd1600,17'd1601,17'd1602,17'd1603,17'd1604,17'd1605,17'd1606,17'd1607,17'd1608,17'd1609,17'd534,17'd1610,17'd1611,17'd1612,17'd1477,17'd1613,17'd1613,17'd719,17'd719,17'd1480,17'd1480,17'd133,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd358,17'd543,17'd726,17'd1614,17'd1615,17'd1616,17'd1617,17'd1618,17'd1619,17'd1620,17'd1621,17'd1622,17'd899,17'd1623,17'd1624,17'd1625,17'd1626,17'd1627,17'd1628,17'd1629,17'd1630,17'd1631,17'd1632,17'd1633,17'd1355,17'd1634,17'd1635,17'd1636,17'd1637,17'd1638,17'd1639,17'd1640,17'd1641,17'd1642,17'd1643,17'd1644,17'd1645,17'd1646,17'd1647,17'd1648,17'd1649,17'd1650,17'd1651,17'd1652,17'd1653,17'd1654,17'd1655,17'd1656,17'd1657,17'd1658,17'd1659,17'd1660,17'd1661,17'd1662,17'd1663,17'd1664,17'd1665,17'd451,17'd607,17'd1666,17'd1667,17'd1668,17'd193,17'd1669,17'd1103,17'd199,17'd1670,17'd1670,17'd198,17'd198,17'd941,17'd1671,17'd1672,17'd194,17'd194,17'd194,17'd417,17'd417,17'd417,17'd418,17'd1673,17'd1673,17'd1532,17'd1531,17'd1251,17'd1674,17'd1534,17'd1534,17'd1675,17'd1535,17'd1388,17'd1389,17'd1676,17'd1677,17'd1099,17'd1272,17'd605,17'd425,17'd259,17'd970,17'd1678,17'd1679,17'd607,17'd443,17'd232,17'd233,17'd245,17'd962,17'd441,17'd1541,17'd770,17'd1543,17'd638,17'd611,17'd210,17'd428,17'd227,17'd446,17'd1263,17'd1262,17'd1262,17'd1680,17'd624,17'd446,17'd227,17'd227,17'd227,17'd227,17'd1402,17'd1402,17'd1402,17'd795,17'd447,17'd959,17'd1546,17'd959,17'd447,17'd447,17'd796,17'd448,17'd234,17'd793,17'd1681,17'd245,17'd1540,17'd212,17'd634,17'd212,17'd1682,17'd461,17'd461,17'd181,17'd639,17'd1683,17'd804,17'd459,17'd1406,17'd968,17'd270,17'd272,17'd644,17'd803,17'd645,17'd803,17'd274,17'd273,17'd641,17'd646,17'd257,17'd459,17'd1684,17'd1271,17'd1270,17'd1270,17'd263,17'd935,17'd803,17'd1111,17'd1685,17'd1272,17'd1381,17'd1245,17'd1686,17'd1410,17'd1687,17'd1273
},
'{
17'd1,17'd1,17'd1,17'd0,17'd2,17'd2,17'd2,17'd0,17'd283,17'd650,17'd808,17'd9,17'd8,17'd8,17'd6,17'd6,17'd4,17'd23,17'd25,17'd25,17'd10,17'd10,17'd283,17'd1412,17'd1,17'd15,17'd1127,17'd1688,17'd1688,17'd1688,17'd1689,17'd1689,17'd1414,17'd1414,17'd17,17'd17,17'd16,17'd16,17'd16,17'd1277,17'd12,17'd12,17'd12,17'd12,17'd3,17'd3,17'd3,17'd3,17'd10,17'd10,17'd10,17'd10,17'd10,17'd10,17'd21,17'd21,17'd25,17'd25,17'd23,17'd23,17'd23,17'd23,17'd23,17'd23,17'd1690,17'd1691,17'd285,17'd285,17'd286,17'd287,17'd28,17'd652,17'd289,17'd468,17'd1692,17'd1692,17'd290,17'd1129,17'd1693,17'd1693,17'd470,17'd470,17'd470,17'd292,17'd656,17'd657,17'd811,17'd295,17'd1694,17'd1553,17'd660,17'd38,17'd1695,17'd1696,17'd1697,17'd1697,17'd1698,17'd1699,17'd1699,17'd1700,17'd1134,17'd1281,17'd1281,17'd1282,17'd1701,17'd1702,17'd1422,17'd1422,17'd1422,17'd1422,17'd1423,17'd1703,17'd1704,17'd1424,17'd1705,17'd1706,17'd1707,17'd1707,17'd1708,17'd1708,17'd1561,17'd1561,17'd1428,17'd1428,17'd1428,17'd1287,17'd1144,17'd1144,17'd1709,17'd1710,17'd669,17'd670,17'd487,17'd69,17'd839,17'd839,17'd840,17'd840,17'd841,17'd491,17'd492,17'd312,17'd76,17'd1711,17'd1712,17'd1713,17'd1714,17'd1715,17'd1716,17'd1717,17'd1717,17'd1718,17'd1718,17'd1719,17'd1720,17'd1721,17'd1722,17'd1723,17'd1724,17'd1725,17'd1726,17'd1727,17'd1728,17'd1729,17'd1730,17'd1731,17'd1732,17'd1733,17'd1734,17'd1735,17'd1736,17'd1737,17'd1738,17'd1739,17'd1740,17'd1741,17'd1742,17'd1743,17'd1744,17'd1745,17'd1746,17'd1747,17'd1748,17'd1749,17'd1750,17'd1751,17'd1752,17'd1753,17'd1754,17'd1755,17'd1756,17'd1757,17'd1333,17'd1758,17'd537,17'd1336,17'd1477,17'd1477,17'd1478,17'd1478,17'd541,17'd541,17'd133,17'd133,17'd133,17'd133,17'd131,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd135,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd132,17'd132,17'd134,17'd1759,17'd358,17'd543,17'd544,17'd1760,17'd1048,17'd547,17'd1761,17'd1762,17'd1763,17'd1764,17'd1765,17'd1766,17'd899,17'd1767,17'd1768,17'd1769,17'd1770,17'd1771,17'd1772,17'd1773,17'd1774,17'd1775,17'd1776,17'd1777,17'd1778,17'd1779,17'd1780,17'd1781,17'd1782,17'd1783,17'd1784,17'd1785,17'd1786,17'd1787,17'd1788,17'd1788,17'd1789,17'd1790,17'd1791,17'd1792,17'd1793,17'd1794,17'd1795,17'd1795,17'd1796,17'd1797,17'd1798,17'd1799,17'd1800,17'd1801,17'd1802,17'd1803,17'd1804,17'd1805,17'd1806,17'd1807,17'd1808,17'd1809,17'd630,17'd232,17'd1680,17'd1810,17'd412,17'd413,17'd776,17'd197,17'd1811,17'd1811,17'd1811,17'd1812,17'd196,17'd417,17'd777,17'd777,17'd418,17'd417,17'd418,17'd599,17'd1530,17'd1530,17'd1673,17'd1813,17'd1814,17'd1815,17'd1251,17'd1674,17'd1675,17'd1675,17'd1535,17'd1535,17'd1816,17'd1817,17'd1818,17'd1819,17'd1820,17'd1821,17'd1098,17'd1410,17'd643,17'd644,17'd970,17'd259,17'd260,17'd427,17'd427,17'd782,17'd1257,17'd442,17'd1092,17'd1822,17'd638,17'd251,17'd592,17'd634,17'd244,17'd234,17'd627,17'd623,17'd954,17'd1262,17'd1823,17'd1823,17'd1261,17'd1261,17'd228,17'd1399,17'd227,17'd446,17'd1824,17'd1825,17'd1402,17'd795,17'd795,17'd795,17'd1264,17'd1264,17'd1264,17'd447,17'd959,17'd959,17'd959,17'd234,17'd793,17'd244,17'd633,17'd245,17'd1540,17'd453,17'd634,17'd611,17'd431,17'd933,17'd431,17'd1826,17'd965,17'd1684,17'd459,17'd257,17'd269,17'd269,17'd643,17'd803,17'd803,17'd803,17'd645,17'd458,17'd274,17'd1268,17'd1407,17'd1267,17'd1271,17'd1270,17'd1270,17'd1270,17'd265,17'd268,17'd274,17'd645,17'd1685,17'd1685,17'd1381,17'd1381,17'd1549,17'd1827,17'd1828,17'd1829
},
'{
17'd1,17'd1,17'd0,17'd2,17'd2,17'd2,17'd0,17'd3,17'd650,17'd465,17'd9,17'd1413,17'd8,17'd8,17'd5,17'd5,17'd23,17'd23,17'd25,17'd21,17'd10,17'd979,17'd1,17'd1830,17'd15,17'd14,17'd1688,17'd1831,17'd1688,17'd1688,17'd1689,17'd1689,17'd1415,17'd1414,17'd1416,17'd16,17'd1277,17'd16,17'd16,17'd1277,17'd12,17'd12,17'd12,17'd12,17'd3,17'd3,17'd283,17'd283,17'd11,17'd11,17'd10,17'd10,17'd10,17'd10,17'd21,17'd21,17'd25,17'd25,17'd23,17'd23,17'd4,17'd4,17'd23,17'd23,17'd1832,17'd467,17'd467,17'd1833,17'd28,17'd652,17'd653,17'd652,17'd289,17'd468,17'd468,17'd468,17'd30,17'd31,17'd1693,17'd1693,17'd1834,17'd470,17'd32,17'd656,17'd984,17'd471,17'd36,17'd985,17'd1553,17'd37,17'd38,17'd1835,17'd1695,17'd1699,17'd1699,17'd1836,17'd1836,17'd1700,17'd1837,17'd1838,17'd1557,17'd1557,17'd1557,17'd1839,17'd1840,17'd1702,17'd1422,17'd1422,17'd1422,17'd1423,17'd1423,17'd1559,17'd1841,17'd1841,17'd1706,17'd1706,17'd1707,17'd1707,17'd1842,17'd1842,17'd1561,17'd1561,17'd1428,17'd1428,17'd1287,17'd1287,17'd1144,17'd1144,17'd1709,17'd1843,17'd837,17'd486,17'd69,17'd70,17'd839,17'd839,17'd840,17'd673,17'd491,17'd1844,17'd1845,17'd1846,17'd1712,17'd1847,17'd1848,17'd1849,17'd1850,17'd1851,17'd1852,17'd1853,17'd1854,17'd1855,17'd1856,17'd1857,17'd1858,17'd1859,17'd1860,17'd1861,17'd1862,17'd1863,17'd1864,17'd1865,17'd1866,17'd1867,17'd1868,17'd1869,17'd1870,17'd1871,17'd1872,17'd1873,17'd1874,17'd1875,17'd1876,17'd1877,17'd1878,17'd1879,17'd1880,17'd1881,17'd1882,17'd1883,17'd1884,17'd1885,17'd1886,17'd1887,17'd1888,17'd1889,17'd1602,17'd1890,17'd1891,17'd1892,17'd1893,17'd1894,17'd710,17'd1895,17'd535,17'd1334,17'd1335,17'd537,17'd1336,17'd1477,17'd538,17'd1478,17'd1195,17'd541,17'd719,17'd719,17'd133,17'd133,17'd541,17'd541,17'd1481,17'd1481,17'd1481,17'd133,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd134,17'd358,17'd358,17'd1482,17'd1482,17'd545,17'd362,17'd546,17'd1896,17'd1761,17'd1897,17'd1050,17'd1898,17'd1899,17'd1900,17'd1901,17'd1902,17'd1903,17'd1904,17'd1905,17'd1906,17'd1907,17'd1908,17'd1909,17'd1910,17'd1911,17'd1912,17'd1913,17'd1914,17'd1915,17'd1916,17'd1917,17'd1918,17'd1792,17'd1919,17'd1919,17'd1920,17'd1921,17'd1922,17'd1923,17'd1924,17'd1925,17'd1926,17'd1927,17'd1928,17'd1929,17'd1930,17'd1931,17'd1932,17'd1933,17'd1934,17'd1935,17'd1936,17'd1937,17'd1938,17'd1939,17'd1940,17'd1941,17'd1808,17'd1942,17'd1943,17'd1944,17'd1945,17'd1810,17'd1946,17'd1383,17'd1672,17'd417,17'd1947,17'd1948,17'd1947,17'd945,17'd1105,17'd1949,17'd1950,17'd1384,17'd599,17'd599,17'd946,17'd1951,17'd1951,17'd1951,17'd1951,17'd1952,17'd1815,17'd1251,17'd1388,17'd1535,17'd1535,17'd1535,17'd1535,17'd1817,17'd1816,17'd1953,17'd1954,17'd1819,17'd1820,17'd1955,17'd1409,17'd605,17'd425,17'd1112,17'd1956,17'd1112,17'd1112,17'd1256,17'd427,17'd1957,17'd1958,17'd1959,17'd1960,17'd933,17'd964,17'd963,17'd963,17'd1092,17'd1961,17'd1239,17'd1239,17'd1240,17'd1962,17'd1823,17'd1396,17'd1261,17'd445,17'd1119,17'd1260,17'd227,17'd446,17'd1824,17'd1825,17'd1402,17'd1402,17'd1402,17'd1402,17'd1402,17'd795,17'd1264,17'd1264,17'd447,17'd959,17'd959,17'd959,17'd959,17'd793,17'd961,17'd244,17'd245,17'd452,17'd634,17'd593,17'd963,17'd964,17'd431,17'd431,17'd804,17'd277,17'd969,17'd459,17'd257,17'd640,17'd206,17'd803,17'd803,17'd645,17'd1963,17'd1963,17'd274,17'd273,17'd272,17'd1407,17'd263,17'd265,17'd265,17'd969,17'd1964,17'd256,17'd273,17'd273,17'd1410,17'd1685,17'd1381,17'd1381,17'd1549,17'd1965,17'd1685,17'd1966
},
'{
17'd1830,17'd15,17'd14,17'd14,17'd2,17'd0,17'd3,17'd283,17'd651,17'd977,17'd9,17'd8,17'd4,17'd4,17'd4,17'd23,17'd23,17'd23,17'd21,17'd21,17'd1275,17'd283,17'd1,17'd15,17'd14,17'd1689,17'd1688,17'd1831,17'd1688,17'd1688,17'd1689,17'd1967,17'd1415,17'd1416,17'd17,17'd16,17'd1277,17'd16,17'd16,17'd1277,17'd12,17'd12,17'd12,17'd12,17'd3,17'd3,17'd1275,17'd1275,17'd11,17'd11,17'd11,17'd10,17'd10,17'd10,17'd21,17'd25,17'd25,17'd25,17'd23,17'd23,17'd4,17'd4,17'd23,17'd23,17'd26,17'd285,17'd467,17'd286,17'd652,17'd653,17'd468,17'd289,17'd468,17'd468,17'd289,17'd29,17'd981,17'd981,17'd654,17'd31,17'd1693,17'd292,17'd1130,17'd656,17'd656,17'd34,17'd1968,17'd1553,17'd1969,17'd38,17'd1970,17'd1970,17'd1970,17'd1700,17'd1700,17'd1837,17'd1838,17'd1838,17'd1971,17'd1972,17'd1972,17'd1973,17'd1974,17'd1974,17'd1975,17'd1974,17'd1976,17'd1977,17'd1423,17'd1423,17'd1283,17'd1559,17'd1841,17'd1706,17'd1706,17'd1706,17'd1978,17'd1978,17'd1842,17'd1842,17'd1561,17'd1561,17'd1979,17'd1428,17'd1428,17'd1287,17'd1287,17'd1144,17'd995,17'd1980,17'd485,17'd1981,17'd69,17'd70,17'd839,17'd839,17'd1982,17'd1983,17'd1984,17'd1985,17'd1986,17'd1986,17'd1987,17'd1988,17'd1989,17'd1990,17'd1991,17'd1992,17'd1993,17'd1994,17'd1995,17'd1996,17'd1997,17'd1998,17'd1999,17'd2000,17'd2001,17'd2002,17'd2003,17'd2004,17'd2005,17'd2006,17'd2007,17'd2008,17'd2009,17'd2010,17'd2011,17'd2012,17'd2013,17'd1872,17'd2014,17'd2015,17'd2016,17'd2017,17'd2018,17'd2019,17'd2020,17'd2021,17'd2022,17'd2023,17'd2024,17'd2025,17'd2026,17'd2027,17'd2028,17'd1888,17'd1600,17'd2029,17'd2030,17'd2031,17'd1891,17'd2032,17'd2033,17'd2034,17'd1756,17'd1757,17'd2035,17'd1192,17'd1332,17'd1193,17'd2036,17'd1334,17'd1194,17'd536,17'd713,17'd713,17'd2037,17'd538,17'd714,17'd1336,17'd2038,17'd1195,17'd2039,17'd2039,17'd2040,17'd1481,17'd1481,17'd1481,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd128,17'd128,17'd1046,17'd2041,17'd1760,17'd2042,17'd2043,17'd2044,17'd2045,17'd2046,17'd1766,17'd2047,17'd2048,17'd2049,17'd2050,17'd2051,17'd2052,17'd2053,17'd2054,17'd2055,17'd2056,17'd2057,17'd2058,17'd2059,17'd2060,17'd2061,17'd2062,17'd2063,17'd2064,17'd2065,17'd2066,17'd2067,17'd2067,17'd2068,17'd2069,17'd2070,17'd2071,17'd2071,17'd2072,17'd2073,17'd2074,17'd2075,17'd2076,17'd2077,17'd2077,17'd2078,17'd2079,17'd2080,17'd2081,17'd2082,17'd2083,17'd2084,17'd2085,17'd2086,17'd2087,17'd2088,17'd2089,17'd2090,17'd2091,17'd2092,17'd2093,17'd2094,17'd2095,17'd2096,17'd2097,17'd2098,17'd777,17'd946,17'd1248,17'd1248,17'd2099,17'd2099,17'd2100,17'd2101,17'd1948,17'd2102,17'd2103,17'd2104,17'd2104,17'd2104,17'd1532,17'd1531,17'd1249,17'd1249,17'd1252,17'd1388,17'd1535,17'd2105,17'd2105,17'd2105,17'd2105,17'd1954,17'd1954,17'd2106,17'd1954,17'd2107,17'd1820,17'd1253,17'd1099,17'd1098,17'd605,17'd425,17'd1396,17'd1666,17'd1666,17'd954,17'd1240,17'd2108,17'd2108,17'd1957,17'd1961,17'd442,17'd431,17'd964,17'd431,17'd2109,17'd2110,17'd2111,17'd2112,17'd1678,17'd1962,17'd1263,17'd1261,17'd445,17'd1119,17'd1260,17'd1399,17'd1260,17'd446,17'd227,17'd446,17'd446,17'd626,17'd623,17'd623,17'd623,17'd443,17'd443,17'd232,17'd232,17'd2113,17'd959,17'd959,17'd234,17'd793,17'd961,17'd633,17'd633,17'd1115,17'd800,17'd792,17'd2114,17'd635,17'd933,17'd456,17'd804,17'd2115,17'd265,17'd256,17'd257,17'd270,17'd273,17'd644,17'd645,17'd1963,17'd1963,17'd803,17'd644,17'd643,17'd272,17'd1268,17'd1405,17'd266,17'd459,17'd1964,17'd459,17'd1268,17'd273,17'd1828,17'd971,17'd1244,17'd1381,17'd2116,17'd2117,17'd603,17'd972
},
'{
17'd15,17'd15,17'd14,17'd14,17'd2,17'd1,17'd283,17'd465,17'd977,17'd977,17'd4,17'd4,17'd4,17'd4,17'd23,17'd23,17'd23,17'd22,17'd21,17'd10,17'd283,17'd1,17'd15,17'd14,17'd1689,17'd1688,17'd1831,17'd1831,17'd1688,17'd1689,17'd1689,17'd1967,17'd1414,17'd1416,17'd17,17'd16,17'd1277,17'd16,17'd16,17'd16,17'd12,17'd12,17'd12,17'd3,17'd3,17'd3,17'd806,17'd806,17'd11,17'd11,17'd11,17'd10,17'd10,17'd808,17'd25,17'd25,17'd25,17'd25,17'd23,17'd23,17'd4,17'd4,17'd23,17'd22,17'd467,17'd26,17'd980,17'd980,17'd652,17'd652,17'd289,17'd468,17'd289,17'd289,17'd29,17'd288,17'd2118,17'd981,17'd31,17'd1129,17'd982,17'd32,17'd656,17'd33,17'd2119,17'd2120,17'd1694,17'd1969,17'd660,17'd660,17'd1700,17'd1700,17'd1700,17'd1837,17'd1837,17'd1838,17'd2121,17'd1972,17'd1972,17'd2122,17'd2122,17'd2122,17'd1974,17'd1974,17'd1975,17'd1974,17'd1977,17'd1977,17'd1423,17'd1423,17'd1283,17'd1283,17'd2123,17'd1706,17'd1706,17'd1706,17'd1707,17'd1707,17'd1842,17'd1842,17'd1561,17'd1561,17'd1979,17'd1428,17'd1428,17'd1287,17'd1287,17'd1144,17'd832,17'd1980,17'd485,17'd1981,17'd69,17'd70,17'd839,17'd72,17'd2124,17'd2125,17'd2126,17'd2127,17'd2128,17'd2129,17'd2129,17'd2130,17'd2131,17'd2132,17'd2133,17'd2134,17'd2135,17'd2136,17'd2137,17'd2138,17'd2139,17'd2140,17'd2141,17'd2001,17'd2142,17'd2143,17'd2144,17'd2145,17'd2146,17'd2147,17'd2148,17'd2149,17'd2150,17'd2151,17'd2152,17'd2153,17'd2013,17'd2154,17'd2155,17'd2156,17'd2157,17'd2158,17'd2159,17'd2159,17'd2160,17'd2160,17'd2161,17'd2162,17'd2163,17'd2164,17'd2165,17'd2166,17'd2167,17'd2168,17'd2169,17'd2170,17'd2029,17'd2171,17'd2172,17'd2173,17'd2174,17'd1754,17'd2175,17'd2176,17'd2177,17'd2178,17'd2179,17'd2180,17'd2181,17'd2182,17'd2182,17'd2183,17'd1757,17'd2184,17'd2184,17'd2184,17'd1193,17'd2185,17'd1194,17'd2186,17'd1336,17'd539,17'd1613,17'd2040,17'd1480,17'd1481,17'd133,17'd133,17'd132,17'd132,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd129,17'd358,17'd543,17'd544,17'd1483,17'd2187,17'd1615,17'd727,17'd2188,17'd2189,17'd2190,17'd2191,17'd2192,17'd2193,17'd2194,17'd2195,17'd2196,17'd2197,17'd2198,17'd2199,17'd2200,17'd2201,17'd2202,17'd2203,17'd2204,17'd2205,17'd2206,17'd2207,17'd2208,17'd2209,17'd2210,17'd2211,17'd2212,17'd2212,17'd2213,17'd2214,17'd2215,17'd2216,17'd2217,17'd2218,17'd2219,17'd2220,17'd2221,17'd2222,17'd2223,17'd2224,17'd2225,17'd2226,17'd2227,17'd2228,17'd2229,17'd2230,17'd2231,17'd2232,17'd2233,17'd2234,17'd2235,17'd2236,17'd2237,17'd2238,17'd2239,17'd2095,17'd2240,17'd1946,17'd779,17'd777,17'd1248,17'd1248,17'd2241,17'd2242,17'd2243,17'd2244,17'd2245,17'd2102,17'd2104,17'd2246,17'd2246,17'd2246,17'd1532,17'd1532,17'd1250,17'd1250,17'd1252,17'd1388,17'd2106,17'd2105,17'd2105,17'd2105,17'd2105,17'd2247,17'd2248,17'd2106,17'd2106,17'd2106,17'd1819,17'd1677,17'd951,17'd602,17'd1668,17'd604,17'd1396,17'd1666,17'd1666,17'd970,17'd953,17'd953,17'd2249,17'd794,17'd2250,17'd1959,17'd442,17'd933,17'd2251,17'd2252,17'd2253,17'd2254,17'd2111,17'd1678,17'd1962,17'd1262,17'd1261,17'd1261,17'd228,17'd1260,17'd1260,17'd1260,17'd227,17'd231,17'd446,17'd446,17'd626,17'd623,17'd623,17'd623,17'd626,17'd626,17'd623,17'd443,17'd1264,17'd1264,17'd447,17'd447,17'd234,17'd793,17'd961,17'd622,17'd450,17'd1115,17'd784,17'd792,17'd454,17'd962,17'd403,17'd456,17'd2255,17'd595,17'd262,17'd256,17'd269,17'd270,17'd644,17'd803,17'd645,17'd645,17'd803,17'd644,17'd643,17'd643,17'd272,17'd968,17'd257,17'd256,17'd802,17'd262,17'd1407,17'd273,17'd1828,17'd971,17'd2256,17'd1381,17'd1245,17'd2116,17'd603,17'd1408
},
'{
17'd1967,17'd1967,17'd14,17'd14,17'd0,17'd3,17'd465,17'd651,17'd977,17'd977,17'd4,17'd4,17'd4,17'd23,17'd23,17'd23,17'd23,17'd22,17'd21,17'd21,17'd1275,17'd3,17'd2,17'd1127,17'd1688,17'd1831,17'd1831,17'd1688,17'd1688,17'd1689,17'd1689,17'd1127,17'd1416,17'd17,17'd16,17'd16,17'd16,17'd16,17'd0,17'd2,17'd12,17'd12,17'd3,17'd3,17'd3,17'd3,17'd806,17'd806,17'd19,17'd19,17'd11,17'd10,17'd10,17'd808,17'd25,17'd25,17'd25,17'd25,17'd22,17'd23,17'd4,17'd4,17'd24,17'd22,17'd285,17'd26,17'd980,17'd1278,17'd652,17'd28,17'd29,17'd29,17'd652,17'd652,17'd28,17'd28,17'd29,17'd289,17'd2257,17'd2258,17'd2259,17'd2259,17'd292,17'd293,17'd2260,17'd2261,17'd1553,17'd660,17'd1837,17'd1837,17'd1837,17'd1837,17'd1838,17'd1971,17'd1971,17'd2121,17'd2260,17'd2262,17'd2263,17'd2264,17'd2264,17'd2263,17'd2265,17'd2265,17'd2265,17'd2266,17'd1976,17'd1976,17'd1422,17'd1422,17'd1558,17'd2267,17'd2268,17'd2268,17'd1706,17'd1706,17'd1707,17'd1707,17'd1842,17'd1561,17'd1561,17'd1561,17'd1979,17'd1979,17'd1428,17'd1428,17'd1287,17'd1145,17'd832,17'd484,17'd1981,17'd1981,17'd69,17'd69,17'd308,17'd308,17'd2269,17'd2270,17'd2271,17'd2272,17'd2273,17'd2274,17'd2274,17'd2275,17'd2276,17'd2277,17'd2278,17'd2279,17'd2280,17'd2281,17'd2282,17'd2283,17'd2284,17'd2285,17'd2286,17'd2287,17'd2288,17'd2289,17'd2290,17'd2291,17'd2292,17'd2293,17'd2294,17'd2295,17'd2296,17'd2297,17'd2298,17'd2299,17'd2300,17'd2301,17'd2302,17'd2303,17'd2304,17'd2305,17'd2305,17'd2306,17'd2307,17'd2308,17'd2161,17'd2309,17'd2310,17'd2311,17'd2312,17'd2026,17'd2313,17'd2314,17'd2315,17'd2316,17'd2317,17'd2318,17'd1601,17'd2319,17'd2320,17'd2321,17'd2031,17'd2322,17'd2323,17'd2324,17'd2324,17'd2325,17'd2326,17'd2327,17'd1189,17'd2328,17'd2329,17'd2330,17'd2331,17'd2332,17'd2333,17'd2334,17'd2335,17'd2336,17'd2337,17'd2338,17'd2339,17'd1612,17'd2340,17'd1479,17'd541,17'd541,17'd1481,17'd1481,17'd134,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd128,17'd129,17'd129,17'd358,17'd1482,17'd1483,17'd548,17'd2341,17'd2342,17'd2343,17'd2344,17'd2345,17'd2346,17'd2193,17'd2347,17'd2348,17'd2349,17'd2350,17'd2351,17'd2352,17'd2353,17'd2354,17'd2355,17'd2356,17'd2357,17'd2358,17'd2359,17'd2360,17'd2361,17'd2362,17'd2363,17'd2364,17'd2365,17'd2366,17'd2367,17'd2368,17'd2369,17'd2370,17'd2371,17'd2220,17'd2372,17'd2373,17'd2374,17'd2375,17'd2375,17'd2376,17'd2377,17'd2378,17'd2379,17'd2380,17'd2381,17'd2382,17'd2383,17'd2384,17'd2385,17'd2386,17'd2387,17'd2388,17'd2389,17'd2390,17'd2391,17'd2392,17'd2393,17'd2394,17'd1950,17'd1105,17'd2099,17'd2395,17'd2396,17'd2396,17'd2397,17'd2397,17'd2398,17'd2399,17'd2400,17'd2400,17'd2400,17'd2246,17'd1250,17'd1250,17'd1252,17'd1389,17'd1953,17'd2401,17'd2402,17'd2403,17'd2404,17'd2405,17'd2405,17'd2105,17'd2105,17'd2406,17'd1818,17'd2407,17'd2408,17'd1383,17'd2409,17'd1668,17'd411,17'd605,17'd970,17'd970,17'd1962,17'd1962,17'd1962,17'd626,17'd2410,17'd2411,17'd2412,17'd2109,17'd224,17'd2413,17'd2414,17'd2415,17'd2416,17'd1239,17'd1380,17'd2417,17'd1261,17'd1401,17'd228,17'd228,17'd228,17'd1260,17'd227,17'd231,17'd227,17'd227,17'd446,17'd446,17'd446,17'd446,17'd626,17'd626,17'd2249,17'd623,17'd443,17'd232,17'd447,17'd447,17'd447,17'd234,17'd448,17'd242,17'd243,17'd238,17'd2418,17'd1115,17'd2419,17'd636,17'd2420,17'd1094,17'd801,17'd255,17'd262,17'd262,17'd1406,17'd968,17'd273,17'd274,17'd645,17'd645,17'd1111,17'd605,17'd425,17'd643,17'd643,17'd272,17'd207,17'd257,17'd257,17'd256,17'd268,17'd273,17'd1828,17'd1828,17'd971,17'd952,17'd598,17'd193,17'd193,17'd193
},
'{
17'd14,17'd14,17'd14,17'd2,17'd12,17'd283,17'd465,17'd977,17'd977,17'd2421,17'd4,17'd4,17'd4,17'd23,17'd23,17'd22,17'd23,17'd22,17'd21,17'd10,17'd283,17'd1,17'd1967,17'd1689,17'd2422,17'd1831,17'd1831,17'd1688,17'd1689,17'd1689,17'd1689,17'd1689,17'd1414,17'd17,17'd16,17'd17,17'd16,17'd1277,17'd0,17'd466,17'd12,17'd12,17'd3,17'd3,17'd3,17'd3,17'd2423,17'd2423,17'd19,17'd19,17'd11,17'd10,17'd808,17'd808,17'd25,17'd9,17'd25,17'd25,17'd22,17'd23,17'd4,17'd4,17'd23,17'd22,17'd26,17'd26,17'd27,17'd980,17'd1278,17'd652,17'd28,17'd2424,17'd28,17'd28,17'd652,17'd29,17'd289,17'd30,17'd2425,17'd2426,17'd982,17'd470,17'd2427,17'd34,17'd2428,17'd2429,17'd1553,17'd1694,17'd1838,17'd1838,17'd1838,17'd1838,17'd2121,17'd1972,17'd2122,17'd2122,17'd2430,17'd2430,17'd2264,17'd2264,17'd2264,17'd2263,17'd2265,17'd2266,17'd2266,17'd2266,17'd2431,17'd2431,17'd2432,17'd2432,17'd2433,17'd2267,17'd2434,17'd2268,17'd1706,17'd1707,17'd1707,17'd2435,17'd1708,17'd1561,17'd1561,17'd1561,17'd1561,17'd2436,17'd2436,17'd2437,17'd2438,17'd994,17'd668,17'd2439,17'd486,17'd487,17'd487,17'd487,17'd309,17'd2440,17'd2441,17'd2442,17'd2443,17'd2444,17'd2445,17'd2446,17'd2447,17'd2448,17'd2449,17'd2450,17'd2451,17'd2280,17'd2452,17'd2453,17'd2454,17'd2455,17'd2456,17'd2457,17'd2458,17'd2459,17'd2289,17'd2460,17'd2461,17'd2462,17'd2463,17'd2464,17'd2465,17'd2466,17'd2467,17'd2467,17'd2298,17'd2299,17'd2468,17'd2468,17'd2469,17'd2470,17'd2471,17'd2472,17'd2473,17'd2474,17'd2475,17'd2476,17'd2477,17'd2478,17'd2479,17'd2480,17'd2481,17'd2482,17'd2483,17'd1745,17'd2484,17'd2485,17'd2486,17'd2487,17'd2488,17'd2489,17'd2490,17'd2491,17'd2492,17'd2493,17'd2494,17'd2495,17'd2496,17'd2497,17'd2497,17'd2498,17'd2499,17'd2500,17'd2501,17'd2502,17'd2326,17'd2503,17'd2504,17'd2505,17'd2505,17'd2506,17'd2507,17'd2508,17'd2509,17'd2510,17'd1611,17'd2511,17'd2340,17'd540,17'd1480,17'd1480,17'd1481,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd128,17'd130,17'd130,17'd130,17'd129,17'd543,17'd141,17'd1337,17'd142,17'd546,17'd1896,17'd2512,17'd2513,17'd2514,17'd2515,17'd2516,17'd2517,17'd2518,17'd2519,17'd2520,17'd2521,17'd2522,17'd2523,17'd2524,17'd2525,17'd2526,17'd2527,17'd2075,17'd2528,17'd2529,17'd2530,17'd2531,17'd2532,17'd2533,17'd2534,17'd2535,17'd2535,17'd2536,17'd2366,17'd2537,17'd2538,17'd2539,17'd2540,17'd2541,17'd2542,17'd2543,17'd2544,17'd2543,17'd2545,17'd2546,17'd2547,17'd2548,17'd2549,17'd2550,17'd2551,17'd2552,17'd2553,17'd2554,17'd2555,17'd2556,17'd2557,17'd2558,17'd2559,17'd412,17'd779,17'd2560,17'd2101,17'd2561,17'd2562,17'd2563,17'd2564,17'd2565,17'd2398,17'd2398,17'd2566,17'd2567,17'd2567,17'd2568,17'd1250,17'd1250,17'd1390,17'd1252,17'd1388,17'd1818,17'd2401,17'd2105,17'd2569,17'd2570,17'd2569,17'd2569,17'd2247,17'd2571,17'd2572,17'd2573,17'd2574,17'd2408,17'd2575,17'd412,17'd2576,17'd2577,17'd411,17'd605,17'd1667,17'd2417,17'd1680,17'd1962,17'd2578,17'd2579,17'd2580,17'd2110,17'd2581,17'd2252,17'd2582,17'd2583,17'd2584,17'd1239,17'd2578,17'd2585,17'd1680,17'd230,17'd1260,17'd1119,17'd2586,17'd228,17'd227,17'd227,17'd231,17'd227,17'd446,17'd625,17'd625,17'd625,17'd625,17'd446,17'd624,17'd2249,17'd443,17'd232,17'd1264,17'd2587,17'd447,17'd447,17'd448,17'd235,17'd451,17'd242,17'd450,17'd784,17'd784,17'd2114,17'd246,17'd1094,17'd2588,17'd967,17'd408,17'd802,17'd256,17'd1406,17'd273,17'd273,17'd803,17'd645,17'd1111,17'd1111,17'd605,17'd425,17'd643,17'd644,17'd271,17'd207,17'd268,17'd256,17'd256,17'd272,17'd274,17'd1687,17'd972,17'd952,17'd598,17'd598,17'd414,17'd2589
},
'{
17'd2590,17'd2590,17'd2,17'd12,17'd283,17'd465,17'd977,17'd2591,17'd23,17'd5,17'd5,17'd5,17'd23,17'd23,17'd2591,17'd2591,17'd21,17'd21,17'd21,17'd10,17'd1,17'd1967,17'd2592,17'd2593,17'd2592,17'd2422,17'd2594,17'd2595,17'd1416,17'd1415,17'd2596,17'd2597,17'd1414,17'd1415,17'd16,17'd16,17'd16,17'd16,17'd12,17'd12,17'd3,17'd3,17'd3,17'd3,17'd12,17'd12,17'd3,17'd3,17'd11,17'd11,17'd11,17'd10,17'd21,17'd25,17'd23,17'd23,17'd23,17'd4,17'd4,17'd4,17'd25,17'd21,17'd21,17'd21,17'd20,17'd20,17'd2598,17'd20,17'd26,17'd286,17'd286,17'd286,17'd980,17'd28,17'd28,17'd29,17'd1692,17'd2599,17'd290,17'd31,17'd1834,17'd2427,17'd33,17'd471,17'd2261,17'd2261,17'd2261,17'd2261,17'd2121,17'd2121,17'd2600,17'd1973,17'd2263,17'd2264,17'd2264,17'd2264,17'd2601,17'd2601,17'd2601,17'd2602,17'd2602,17'd2602,17'd2602,17'd2603,17'd2604,17'd2604,17'd2605,17'd2606,17'd2607,17'd2607,17'd2267,17'd2608,17'd2268,17'd1978,17'd1707,17'd2435,17'd2435,17'd2609,17'd2609,17'd2435,17'd2435,17'd2610,17'd2611,17'd2436,17'd2612,17'd994,17'd832,17'd668,17'd2613,17'd2614,17'd2615,17'd2616,17'd2616,17'd2617,17'd2618,17'd2619,17'd2620,17'd2621,17'd2622,17'd2623,17'd2624,17'd2625,17'd2626,17'd2627,17'd2628,17'd2629,17'd2630,17'd2631,17'd2632,17'd2633,17'd2634,17'd2635,17'd2636,17'd2637,17'd2638,17'd2639,17'd2640,17'd2641,17'd2642,17'd2643,17'd2644,17'd2645,17'd2646,17'd2647,17'd2648,17'd2649,17'd2650,17'd2651,17'd2652,17'd2653,17'd2654,17'd2655,17'd2656,17'd2656,17'd2657,17'd2468,17'd2658,17'd2659,17'd2476,17'd2478,17'd2660,17'd2661,17'd2662,17'd2663,17'd2664,17'd2665,17'd2666,17'd1745,17'd2667,17'd2668,17'd2028,17'd2669,17'd2670,17'd2671,17'd2672,17'd2673,17'd2674,17'd2675,17'd2676,17'd2677,17'd2678,17'd2679,17'd2680,17'd2681,17'd2682,17'd2683,17'd2684,17'd2685,17'd2686,17'd2687,17'd2688,17'd2689,17'd2690,17'd2691,17'd2692,17'd2693,17'd2694,17'd2695,17'd2696,17'd2697,17'd538,17'd539,17'd2039,17'd1480,17'd542,17'd542,17'd542,17'd133,17'd133,17'd133,17'd132,17'd132,17'd135,17'd135,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd135,17'd132,17'd132,17'd134,17'd134,17'd130,17'd358,17'd358,17'd130,17'd130,17'd543,17'd129,17'd2698,17'd2699,17'd2700,17'd2701,17'd2702,17'd2703,17'd2704,17'd2705,17'd2706,17'd2707,17'd2708,17'd2709,17'd2710,17'd2711,17'd2712,17'd2713,17'd2714,17'd2715,17'd2716,17'd2717,17'd2718,17'd2719,17'd2720,17'd2720,17'd2721,17'd2722,17'd2723,17'd2724,17'd2724,17'd2725,17'd2543,17'd2542,17'd2726,17'd2726,17'd2727,17'd2727,17'd2542,17'd2728,17'd2729,17'd2730,17'd2731,17'd2731,17'd2732,17'd2733,17'd2734,17'd2735,17'd2554,17'd2736,17'd2737,17'd2738,17'd629,17'd2739,17'd2740,17'd413,17'd2394,17'd2741,17'd2742,17'd2743,17'd2744,17'd2745,17'd2746,17'd2747,17'd2568,17'd2568,17'd2748,17'd2749,17'd2750,17'd2751,17'd1386,17'd2752,17'd1387,17'd1388,17'd1816,17'd2753,17'd2754,17'd2755,17'd2756,17'd2757,17'd2756,17'd2758,17'd2759,17'd2760,17'd2402,17'd2761,17'd1677,17'd602,17'd2762,17'd2763,17'd1382,17'd1393,17'd191,17'd2764,17'd2765,17'd1962,17'd1240,17'd2766,17'd2767,17'd2768,17'd2769,17'd2412,17'd2581,17'd2581,17'd2770,17'd2771,17'd2772,17'd2773,17'd2774,17'd2775,17'd1962,17'd1263,17'd1262,17'd1680,17'd625,17'd227,17'd2776,17'd1399,17'd1260,17'd228,17'd228,17'd228,17'd228,17'd625,17'd2777,17'd2777,17'd624,17'd626,17'd443,17'd232,17'd447,17'd2587,17'd1122,17'd1122,17'd1122,17'd234,17'd961,17'd244,17'd633,17'd633,17'd211,17'd1094,17'd610,17'd967,17'd2778,17'd256,17'd256,17'd257,17'd272,17'd272,17'd644,17'd645,17'd411,17'd411,17'd605,17'd425,17'd2779,17'd270,17'd1268,17'd1268,17'd1407,17'd968,17'd269,17'd269,17'd274,17'd803,17'd971,17'd1685,17'd1244,17'd1381,17'd422,17'd1527
},
'{
17'd2780,17'd2780,17'd12,17'd3,17'd1275,17'd465,17'd2591,17'd2591,17'd23,17'd5,17'd5,17'd5,17'd23,17'd23,17'd2591,17'd2591,17'd21,17'd21,17'd10,17'd979,17'd15,17'd2781,17'd2782,17'd2783,17'd2782,17'd2784,17'd2594,17'd2595,17'd1416,17'd1415,17'd2596,17'd2596,17'd1415,17'd1415,17'd16,17'd16,17'd16,17'd16,17'd12,17'd3,17'd3,17'd3,17'd3,17'd3,17'd12,17'd12,17'd3,17'd3,17'd11,17'd11,17'd10,17'd10,17'd21,17'd25,17'd23,17'd23,17'd4,17'd4,17'd4,17'd4,17'd25,17'd21,17'd21,17'd21,17'd21,17'd20,17'd20,17'd21,17'd285,17'd467,17'd467,17'd285,17'd27,17'd28,17'd29,17'd289,17'd30,17'd1129,17'd1129,17'd1693,17'd470,17'd293,17'd294,17'd471,17'd2261,17'd2261,17'd2261,17'd2261,17'd1973,17'd2600,17'd2785,17'd2785,17'd2602,17'd2601,17'd2601,17'd2601,17'd2601,17'd2601,17'd2602,17'd2602,17'd2602,17'd2602,17'd2601,17'd2601,17'd2604,17'd2604,17'd2605,17'd2606,17'd2607,17'd2607,17'd2608,17'd2608,17'd2786,17'd1978,17'd1707,17'd2435,17'd2435,17'd2609,17'd2609,17'd2435,17'd2435,17'd2610,17'd2787,17'd2788,17'd2789,17'd2790,17'd2791,17'd484,17'd996,17'd1290,17'd2792,17'd2792,17'd2793,17'd2794,17'd2795,17'd2796,17'd2797,17'd2798,17'd2799,17'd2800,17'd2801,17'd2626,17'd2802,17'd2628,17'd2803,17'd2804,17'd2805,17'd2806,17'd2807,17'd2808,17'd2809,17'd2810,17'd2811,17'd2812,17'd2813,17'd2814,17'd2815,17'd2816,17'd2817,17'd2818,17'd2819,17'd2646,17'd2820,17'd2821,17'd2648,17'd2822,17'd2822,17'd2822,17'd2823,17'd2824,17'd2824,17'd2824,17'd2824,17'd2825,17'd2826,17'd2827,17'd2302,17'd2659,17'd2828,17'd2829,17'd2021,17'd2830,17'd2831,17'd2832,17'd2833,17'd2834,17'd2664,17'd2665,17'd2835,17'd2836,17'd2837,17'd2838,17'd2838,17'd2839,17'd2840,17'd2841,17'd2842,17'd2843,17'd2844,17'd2676,17'd2845,17'd2846,17'd2847,17'd2495,17'd2848,17'd2849,17'd2501,17'd2850,17'd2851,17'd2852,17'd2853,17'd1754,17'd2854,17'd2855,17'd2334,17'd2335,17'd2336,17'd2856,17'd2857,17'd2696,17'd2858,17'd2859,17'd1478,17'd2039,17'd719,17'd542,17'd542,17'd542,17'd542,17'd1197,17'd1197,17'd1197,17'd132,17'd132,17'd132,17'd132,17'd133,17'd1197,17'd1197,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd2698,17'd2860,17'd2861,17'd2862,17'd2863,17'd2864,17'd2865,17'd2866,17'd2867,17'd2868,17'd2869,17'd2870,17'd2871,17'd2872,17'd2873,17'd2874,17'd2875,17'd2876,17'd2877,17'd2878,17'd2879,17'd2880,17'd2881,17'd2882,17'd2883,17'd2884,17'd2885,17'd2886,17'd2887,17'd2887,17'd2888,17'd2889,17'd2723,17'd2724,17'd2536,17'd2890,17'd2891,17'd2892,17'd2892,17'd2890,17'd2542,17'd2893,17'd2894,17'd2895,17'd2896,17'd2896,17'd2897,17'd2898,17'd2899,17'd2900,17'd2901,17'd2902,17'd2903,17'd2904,17'd630,17'd2739,17'd2905,17'd2097,17'd2906,17'd2907,17'd2908,17'd2909,17'd2746,17'd2910,17'd2910,17'd2911,17'd2911,17'd2912,17'd2912,17'd2913,17'd2914,17'd2752,17'd1386,17'd1386,17'd1386,17'd1534,17'd2915,17'd2754,17'd2755,17'd2756,17'd2756,17'd2916,17'd2917,17'd2918,17'd2919,17'd2403,17'd2402,17'd1819,17'd1677,17'd780,17'd601,17'd415,17'd2920,17'd2921,17'd2922,17'd2775,17'd2765,17'd2923,17'd2924,17'd2773,17'd2925,17'd2926,17'd2927,17'd2770,17'd2928,17'd2770,17'd2771,17'd2929,17'd2580,17'd2930,17'd2585,17'd2765,17'd1962,17'd1262,17'd1262,17'd625,17'd446,17'd1399,17'd1399,17'd1260,17'd1260,17'd228,17'd1119,17'd1119,17'd1119,17'd2586,17'd2586,17'd2586,17'd624,17'd446,17'd623,17'd795,17'd447,17'd447,17'd226,17'd226,17'd1122,17'd234,17'd961,17'd1681,17'd1681,17'd2931,17'd1094,17'd610,17'd1096,17'd2778,17'd2778,17'd257,17'd257,17'd270,17'd272,17'd644,17'd645,17'd411,17'd1111,17'd1111,17'd605,17'd206,17'd270,17'd1268,17'd1268,17'd1268,17'd1407,17'd270,17'd270,17'd274,17'd803,17'd971,17'd1685,17'd1244,17'd1381,17'd2932,17'd1527
},
'{
17'd0,17'd0,17'd3,17'd283,17'd650,17'd465,17'd25,17'd25,17'd4,17'd4,17'd5,17'd5,17'd23,17'd23,17'd2933,17'd1275,17'd10,17'd10,17'd979,17'd1277,17'd1689,17'd2422,17'd2593,17'd2934,17'd2935,17'd2422,17'd1688,17'd1127,17'd1414,17'd1414,17'd2596,17'd2936,17'd1415,17'd17,17'd16,17'd16,17'd16,17'd16,17'd3,17'd3,17'd3,17'd3,17'd12,17'd12,17'd13,17'd12,17'd12,17'd3,17'd10,17'd10,17'd10,17'd10,17'd21,17'd25,17'd23,17'd23,17'd5,17'd5,17'd4,17'd23,17'd22,17'd22,17'd20,17'd21,17'd21,17'd21,17'd21,17'd25,17'd467,17'd2937,17'd467,17'd467,17'd286,17'd980,17'd2938,17'd468,17'd809,17'd654,17'd31,17'd469,17'd292,17'd32,17'd656,17'd656,17'd2939,17'd2939,17'd2939,17'd2939,17'd2263,17'd2785,17'd2602,17'd2601,17'd2940,17'd2941,17'd2942,17'd2943,17'd2944,17'd2944,17'd2602,17'd2602,17'd2602,17'd2601,17'd2945,17'd2945,17'd2945,17'd2946,17'd2605,17'd2947,17'd2948,17'd2607,17'd2608,17'd2608,17'd2608,17'd2786,17'd2786,17'd2435,17'd2435,17'd2435,17'd1842,17'd1842,17'd1708,17'd1708,17'd2949,17'd1141,17'd993,17'd1145,17'd996,17'd669,17'd2950,17'd835,17'd2951,17'd2951,17'd2952,17'd2953,17'd2954,17'd2954,17'd2955,17'd2956,17'd2957,17'd2958,17'd2959,17'd2960,17'd2961,17'd2629,17'd2962,17'd2963,17'd2964,17'd2965,17'd2966,17'd2967,17'd2968,17'd2969,17'd2970,17'd2971,17'd2972,17'd2973,17'd2974,17'd2643,17'd2975,17'd2976,17'd2977,17'd2464,17'd2978,17'd2979,17'd2980,17'd2981,17'd2982,17'd2983,17'd2984,17'd2985,17'd2986,17'd2987,17'd2988,17'd2989,17'd2990,17'd2991,17'd2992,17'd2993,17'd2994,17'd2995,17'd2996,17'd2997,17'd2020,17'd2830,17'd2998,17'd2999,17'd3000,17'd3001,17'd3002,17'd3003,17'd1884,17'd3004,17'd3005,17'd3006,17'd3007,17'd3008,17'd2672,17'd2674,17'd1749,17'd3009,17'd3010,17'd3011,17'd3012,17'd3013,17'd3014,17'd3015,17'd3016,17'd3017,17'd3018,17'd3019,17'd1892,17'd2175,17'd3020,17'd2180,17'd3021,17'd1757,17'd3022,17'd3023,17'd3024,17'd712,17'd2858,17'd2859,17'd1478,17'd1613,17'd1480,17'd1480,17'd1480,17'd541,17'd541,17'd541,17'd1196,17'd1196,17'd719,17'd542,17'd133,17'd1197,17'd134,17'd134,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd3025,17'd3025,17'd3025,17'd1759,17'd135,17'd2861,17'd2862,17'd3026,17'd3027,17'd3028,17'd3029,17'd3030,17'd3031,17'd3032,17'd3033,17'd3034,17'd3035,17'd3036,17'd3037,17'd3038,17'd3039,17'd3040,17'd3041,17'd3042,17'd3043,17'd3044,17'd3045,17'd3046,17'd3047,17'd3048,17'd3049,17'd3050,17'd3051,17'd3052,17'd3053,17'd3053,17'd3051,17'd2885,17'd2720,17'd3054,17'd3055,17'd2534,17'd2536,17'd3056,17'd3056,17'd3057,17'd3058,17'd3059,17'd3060,17'd3061,17'd3062,17'd3063,17'd3064,17'd3065,17'd3062,17'd2894,17'd3066,17'd3067,17'd3068,17'd3069,17'd3070,17'd3071,17'd3072,17'd1810,17'd3073,17'd3074,17'd3075,17'd3076,17'd2748,17'd3077,17'd3078,17'd3078,17'd3078,17'd3077,17'd3079,17'd3080,17'd3081,17'd3081,17'd1387,17'd1674,17'd1251,17'd1534,17'd1535,17'd2754,17'd2569,17'd3082,17'd3082,17'd3083,17'd3083,17'd3083,17'd3083,17'd3083,17'd2756,17'd3084,17'd3085,17'd3086,17'd2762,17'd3086,17'd3086,17'd3087,17'd3088,17'd3089,17'd3090,17'd2923,17'd2923,17'd3091,17'd3092,17'd3093,17'd2926,17'd2929,17'd2770,17'd2770,17'd2110,17'd2771,17'd3094,17'd2773,17'd3095,17'd3096,17'd3097,17'd1962,17'd953,17'd1262,17'd1680,17'd230,17'd3098,17'd1399,17'd1260,17'd228,17'd1119,17'd1119,17'd1119,17'd3099,17'd2586,17'd2586,17'd2777,17'd2777,17'd2249,17'd443,17'd428,17'd2587,17'd2587,17'd2587,17'd2587,17'd447,17'd959,17'd1546,17'd961,17'd1681,17'd961,17'd429,17'd3100,17'd2778,17'd2778,17'd257,17'd257,17'd269,17'd270,17'd644,17'd645,17'd645,17'd645,17'd1111,17'd645,17'd273,17'd270,17'd270,17'd272,17'd273,17'd272,17'd272,17'd272,17'd274,17'd274,17'd1410,17'd1685,17'd1244,17'd1381,17'd422,17'd1246
},
'{
17'd0,17'd1,17'd283,17'd283,17'd650,17'd465,17'd25,17'd25,17'd4,17'd4,17'd5,17'd4,17'd23,17'd25,17'd1275,17'd1275,17'd10,17'd979,17'd1277,17'd1415,17'd2422,17'd3101,17'd3101,17'd2934,17'd2935,17'd2422,17'd1689,17'd1127,17'd1414,17'd2257,17'd2596,17'd1415,17'd16,17'd16,17'd16,17'd16,17'd16,17'd16,17'd3,17'd3,17'd3,17'd12,17'd12,17'd13,17'd13,17'd12,17'd12,17'd3,17'd10,17'd10,17'd10,17'd808,17'd25,17'd25,17'd23,17'd23,17'd5,17'd5,17'd23,17'd23,17'd22,17'd22,17'd21,17'd21,17'd25,17'd25,17'd9,17'd9,17'd2937,17'd467,17'd285,17'd286,17'd27,17'd652,17'd289,17'd809,17'd3102,17'd654,17'd1693,17'd982,17'd32,17'd32,17'd33,17'd33,17'd2260,17'd2260,17'd2939,17'd3103,17'd2264,17'd2601,17'd2601,17'd3104,17'd2941,17'd2941,17'd2941,17'd2940,17'd2944,17'd2944,17'd2944,17'd2601,17'd2601,17'd3105,17'd3106,17'd3106,17'd2945,17'd2946,17'd2947,17'd2431,17'd3107,17'd3107,17'd2608,17'd2608,17'd2608,17'd2608,17'd2608,17'd2786,17'd1978,17'd2435,17'd1842,17'd1842,17'd1708,17'd3108,17'd2949,17'd1141,17'd1143,17'd1145,17'd1710,17'd998,17'd2950,17'd997,17'd1147,17'd3109,17'd3110,17'd3111,17'd3111,17'd3112,17'd2956,17'd3113,17'd3114,17'd3115,17'd3116,17'd2451,17'd3117,17'd2804,17'd3118,17'd3119,17'd3120,17'd3121,17'd3122,17'd3123,17'd3124,17'd3125,17'd3126,17'd3127,17'd3128,17'd3129,17'd3130,17'd3131,17'd3132,17'd2976,17'd2976,17'd3133,17'd3133,17'd3133,17'd3134,17'd3135,17'd2984,17'd3136,17'd3137,17'd3138,17'd3139,17'd3140,17'd3141,17'd3142,17'd3143,17'd3144,17'd3145,17'd3146,17'd3147,17'd2994,17'd2157,17'd2158,17'd2017,17'd2018,17'd2022,17'd2023,17'd3148,17'd3149,17'd3150,17'd3151,17'd3152,17'd1884,17'd3153,17'd3154,17'd3155,17'd3156,17'd3157,17'd3158,17'd1750,17'd3159,17'd2319,17'd3160,17'd3161,17'd3014,17'd3015,17'd3162,17'd1189,17'd1189,17'd3018,17'd2174,17'd1754,17'd3163,17'd2854,17'd3164,17'd3021,17'd1757,17'd3023,17'd3165,17'd3166,17'd2186,17'd713,17'd2037,17'd2037,17'd1478,17'd1479,17'd1196,17'd1196,17'd541,17'd540,17'd1195,17'd1195,17'd1195,17'd3167,17'd1044,17'd719,17'd1197,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd133,17'd133,17'd133,17'd133,17'd133,17'd132,17'd3168,17'd3169,17'd3170,17'd3171,17'd3172,17'd3173,17'd3174,17'd3175,17'd3176,17'd3177,17'd3178,17'd3179,17'd3180,17'd3181,17'd3182,17'd3183,17'd3184,17'd3185,17'd3186,17'd3187,17'd3188,17'd3189,17'd3190,17'd3191,17'd3192,17'd3193,17'd3194,17'd3195,17'd3196,17'd3197,17'd3198,17'd3199,17'd3200,17'd3201,17'd3201,17'd3202,17'd3203,17'd3204,17'd3205,17'd3206,17'd3207,17'd3207,17'd3208,17'd2535,17'd2535,17'd3209,17'd3210,17'd3211,17'd3212,17'd3213,17'd3214,17'd3215,17'd3216,17'd3216,17'd3217,17'd3218,17'd3219,17'd3220,17'd3221,17'd3222,17'd1825,17'd2392,17'd2098,17'd3223,17'd3224,17'd3225,17'd3226,17'd3078,17'd3227,17'd3227,17'd3228,17'd3078,17'd3229,17'd3229,17'd3229,17'd3229,17'd3230,17'd3231,17'd1534,17'd1389,17'd1535,17'd2404,17'd2405,17'd3082,17'd3083,17'd3083,17'd3232,17'd3232,17'd3233,17'd3083,17'd3232,17'd3083,17'd3234,17'd1392,17'd3086,17'd3235,17'd3236,17'd3237,17'd3238,17'd3239,17'd2774,17'd3240,17'd3240,17'd3091,17'd3241,17'd3242,17'd3243,17'd2771,17'd2770,17'd2412,17'd2771,17'd2580,17'd3244,17'd2930,17'd3096,17'd3095,17'd3245,17'd953,17'd1263,17'd1680,17'd1401,17'd230,17'd1399,17'd1260,17'd228,17'd2586,17'd2586,17'd1119,17'd3246,17'd3246,17'd3246,17'd3247,17'd3247,17'd2777,17'd446,17'd443,17'd795,17'd447,17'd2587,17'd2587,17'd3248,17'd2587,17'd447,17'd1546,17'd1546,17'd793,17'd429,17'd3100,17'd609,17'd608,17'd608,17'd257,17'd207,17'd270,17'd644,17'd803,17'd645,17'd645,17'd411,17'd1963,17'd803,17'd272,17'd269,17'd272,17'd273,17'd272,17'd272,17'd273,17'd273,17'd803,17'd971,17'd971,17'd1244,17'd1381,17'd422,17'd1246
},
'{
17'd1,17'd1,17'd283,17'd650,17'd808,17'd808,17'd25,17'd25,17'd4,17'd4,17'd4,17'd23,17'd23,17'd25,17'd10,17'd979,17'd19,17'd1277,17'd3249,17'd3250,17'd3101,17'd3251,17'd3251,17'd3101,17'd3252,17'd3250,17'd2781,17'd1689,17'd2597,17'd2597,17'd2257,17'd1415,17'd16,17'd16,17'd17,17'd17,17'd0,17'd0,17'd3,17'd3,17'd12,17'd12,17'd13,17'd13,17'd13,17'd12,17'd18,17'd19,17'd10,17'd10,17'd21,17'd25,17'd23,17'd4,17'd5,17'd5,17'd5,17'd24,17'd24,17'd24,17'd23,17'd23,17'd23,17'd23,17'd9,17'd9,17'd9,17'd9,17'd467,17'd285,17'd27,17'd27,17'd980,17'd652,17'd29,17'd29,17'd981,17'd31,17'd982,17'd2259,17'd2259,17'd2259,17'd3253,17'd3253,17'd2262,17'd2262,17'd2262,17'd3253,17'd2942,17'd2941,17'd2941,17'd3254,17'd3255,17'd3255,17'd3254,17'd3256,17'd3257,17'd3256,17'd3104,17'd3105,17'd3258,17'd3259,17'd2945,17'd2945,17'd2606,17'd2431,17'd2948,17'd3260,17'd3261,17'd3261,17'd2608,17'd2608,17'd3107,17'd3107,17'd2267,17'd2268,17'd1978,17'd1707,17'd2610,17'd3262,17'd1427,17'd1427,17'd3263,17'd3263,17'd3264,17'd1146,17'd1146,17'd3265,17'd1146,17'd3266,17'd3267,17'd3268,17'd3269,17'd3270,17'd3271,17'd3272,17'd2800,17'd2958,17'd3273,17'd3274,17'd3275,17'd3276,17'd3277,17'd3278,17'd3279,17'd3280,17'd3281,17'd3282,17'd3283,17'd3284,17'd3285,17'd3286,17'd3287,17'd3288,17'd3289,17'd3290,17'd3291,17'd3292,17'd3132,17'd3293,17'd3293,17'd2984,17'd2984,17'd3294,17'd3295,17'd3296,17'd3297,17'd3298,17'd3299,17'd3300,17'd3300,17'd3301,17'd3302,17'd3303,17'd3304,17'd3305,17'd3306,17'd3307,17'd3145,17'd3146,17'd3308,17'd2303,17'd3309,17'd3310,17'd3311,17'd3312,17'd3313,17'd3314,17'd3315,17'd3316,17'd3317,17'd1884,17'd3318,17'd3319,17'd3320,17'd2676,17'd1600,17'd3321,17'd3322,17'd3323,17'd3324,17'd3161,17'd1890,17'd3325,17'd3326,17'd3327,17'd2325,17'd2325,17'd3328,17'd3329,17'd3330,17'd3331,17'd1755,17'd3164,17'd2182,17'd1331,17'd1757,17'd883,17'd3023,17'd1193,17'd712,17'd536,17'd1612,17'd3332,17'd3333,17'd3333,17'd3334,17'd1478,17'd2037,17'd2037,17'd3335,17'd3335,17'd3336,17'd3337,17'd719,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd134,17'd3168,17'd3338,17'd3339,17'd3340,17'd3341,17'd3342,17'd3343,17'd3344,17'd3345,17'd3346,17'd3347,17'd3348,17'd3349,17'd3350,17'd3351,17'd3352,17'd3353,17'd3354,17'd3355,17'd3356,17'd3357,17'd3358,17'd3359,17'd3360,17'd3361,17'd3362,17'd3363,17'd3364,17'd3365,17'd3366,17'd3367,17'd3368,17'd3369,17'd3370,17'd3371,17'd3372,17'd3373,17'd3374,17'd3375,17'd3206,17'd3376,17'd3206,17'd3206,17'd3205,17'd2886,17'd3377,17'd3208,17'd2535,17'd3378,17'd3379,17'd3380,17'd3381,17'd3381,17'd3382,17'd3383,17'd3384,17'd3385,17'd3386,17'd3387,17'd3388,17'd3389,17'd3390,17'd1825,17'd3391,17'd2098,17'd3392,17'd3393,17'd3394,17'd3395,17'd3396,17'd3397,17'd3398,17'd3399,17'd3399,17'd3400,17'd3401,17'd3401,17'd3402,17'd3403,17'd1817,17'd1389,17'd1535,17'd2753,17'd2247,17'd3404,17'd3082,17'd3082,17'd3405,17'd3406,17'd3407,17'd3407,17'd3407,17'd3408,17'd3405,17'd3409,17'd3410,17'd3235,17'd3411,17'd3411,17'd3412,17'd3413,17'd3414,17'd3415,17'd2923,17'd3092,17'd3416,17'd2926,17'd3417,17'd3418,17'd2412,17'd2770,17'd3419,17'd2771,17'd2580,17'd3244,17'd3420,17'd3421,17'd3422,17'd2739,17'd1263,17'd1262,17'd1401,17'd230,17'd230,17'd230,17'd228,17'd1119,17'd2586,17'd2586,17'd3423,17'd3424,17'd3425,17'd3423,17'd3423,17'd3247,17'd1119,17'd446,17'd3426,17'd1264,17'd1264,17'd795,17'd1402,17'd1402,17'd795,17'd447,17'd447,17'd959,17'd959,17'd233,17'd428,17'd607,17'd1539,17'd258,17'd258,17'd207,17'd643,17'd644,17'd803,17'd645,17'd973,17'd1550,17'd1410,17'd1124,17'd269,17'd270,17'd272,17'd272,17'd272,17'd273,17'd644,17'd803,17'd971,17'd971,17'd1272,17'd952,17'd422,17'd422
},
'{
17'd1,17'd1412,17'd650,17'd650,17'd808,17'd808,17'd25,17'd25,17'd4,17'd4,17'd23,17'd23,17'd25,17'd808,17'd979,17'd979,17'd16,17'd2936,17'd3250,17'd2935,17'd3427,17'd3428,17'd3101,17'd2935,17'd2422,17'd3250,17'd2781,17'd3250,17'd3429,17'd2258,17'd2257,17'd1414,17'd16,17'd16,17'd17,17'd16,17'd0,17'd0,17'd12,17'd12,17'd13,17'd13,17'd3430,17'd13,17'd13,17'd12,17'd19,17'd19,17'd10,17'd10,17'd21,17'd25,17'd23,17'd4,17'd5,17'd6,17'd5,17'd24,17'd24,17'd24,17'd23,17'd4,17'd4,17'd4,17'd9,17'd9,17'd9,17'd25,17'd285,17'd26,17'd980,17'd980,17'd652,17'd28,17'd288,17'd2118,17'd654,17'd1129,17'd982,17'd982,17'd982,17'd982,17'd2940,17'd2943,17'd2943,17'd3253,17'd2943,17'd2940,17'd3431,17'd3254,17'd3254,17'd3255,17'd3255,17'd3255,17'd3254,17'd3254,17'd3432,17'd3433,17'd3434,17'd3435,17'd3258,17'd3259,17'd2945,17'd2946,17'd2431,17'd2431,17'd2948,17'd3260,17'd3261,17'd3261,17'd2608,17'd2608,17'd3107,17'd1422,17'd2267,17'd2268,17'd1978,17'd2610,17'd2611,17'd2611,17'd1427,17'd1427,17'd1427,17'd1427,17'd3436,17'd3437,17'd3438,17'd3438,17'd3439,17'd3440,17'd3441,17'd3442,17'd3443,17'd3444,17'd3445,17'd3446,17'd3447,17'd3448,17'd3449,17'd3275,17'd3450,17'd3118,17'd3451,17'd3452,17'd3453,17'd3454,17'd3455,17'd3456,17'd3457,17'd3458,17'd3459,17'd3460,17'd3461,17'd3462,17'd3463,17'd3464,17'd3465,17'd3466,17'd3467,17'd3295,17'd3295,17'd3468,17'd3469,17'd3470,17'd3470,17'd3471,17'd3472,17'd3473,17'd3474,17'd3475,17'd3475,17'd3476,17'd3477,17'd3478,17'd3479,17'd3480,17'd3481,17'd3482,17'd3483,17'd3484,17'd3485,17'd3486,17'd3487,17'd3488,17'd3489,17'd3312,17'd2162,17'd3490,17'd3491,17'd3492,17'd3493,17'd3494,17'd3495,17'd3496,17'd3497,17'd2488,17'd1750,17'd3498,17'd3499,17'd3500,17'd3501,17'd2500,17'd3502,17'd3503,17'd3504,17'd1604,17'd3505,17'd2326,17'd2503,17'd3506,17'd3507,17'd3508,17'd2690,17'd2033,17'd3509,17'd3510,17'd2183,17'd1757,17'd3022,17'd711,17'd2338,17'd712,17'd536,17'd1476,17'd1476,17'd1476,17'd1476,17'd1612,17'd2859,17'd2859,17'd3511,17'd3336,17'd3337,17'd1196,17'd542,17'd133,17'd133,17'd132,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd133,17'd132,17'd135,17'd2698,17'd2860,17'd3512,17'd3513,17'd3514,17'd3515,17'd3516,17'd3517,17'd3518,17'd3519,17'd3520,17'd3521,17'd3522,17'd3523,17'd3524,17'd3525,17'd3526,17'd3527,17'd3528,17'd3529,17'd3530,17'd3531,17'd3532,17'd3533,17'd3534,17'd3535,17'd3536,17'd3537,17'd3538,17'd3539,17'd3540,17'd3541,17'd3542,17'd3543,17'd3544,17'd3545,17'd3546,17'd3547,17'd3548,17'd3549,17'd3550,17'd3551,17'd3552,17'd3553,17'd3554,17'd3554,17'd3552,17'd3555,17'd3556,17'd3557,17'd3558,17'd3559,17'd3560,17'd3560,17'd3561,17'd3562,17'd3563,17'd3384,17'd3384,17'd3564,17'd3565,17'd3566,17'd3567,17'd3568,17'd3569,17'd1825,17'd2392,17'd3570,17'd3392,17'd3571,17'd3394,17'd3572,17'd3573,17'd3574,17'd3574,17'd3574,17'd3398,17'd3400,17'd3400,17'd3402,17'd3575,17'd3403,17'd1817,17'd1535,17'd1535,17'd2105,17'd2247,17'd3082,17'd3082,17'd3405,17'd3406,17'd3576,17'd3577,17'd3578,17'd3408,17'd3408,17'd3405,17'd3579,17'd3580,17'd3581,17'd3582,17'd3237,17'd3583,17'd3413,17'd3584,17'd3585,17'd3586,17'd3095,17'd3241,17'd3417,17'd3243,17'd2929,17'd2770,17'd3587,17'd3419,17'd2929,17'd3588,17'd2580,17'd3589,17'd3421,17'd3590,17'd1680,17'd1262,17'd1261,17'd1401,17'd230,17'd230,17'd1260,17'd228,17'd2586,17'd3246,17'd3425,17'd3425,17'd3425,17'd3425,17'd3423,17'd3423,17'd2586,17'd2586,17'd3591,17'd1825,17'd3426,17'd795,17'd795,17'd1402,17'd1402,17'd1402,17'd2587,17'd447,17'd447,17'd447,17'd428,17'd782,17'd607,17'd1539,17'd207,17'd207,17'd2779,17'd643,17'd803,17'd645,17'd973,17'd973,17'd973,17'd1828,17'd272,17'd270,17'd270,17'd272,17'd272,17'd272,17'd644,17'd803,17'd971,17'd971,17'd1272,17'd952,17'd1382,17'd422
},
'{
17'd283,17'd283,17'd650,17'd650,17'd10,17'd808,17'd25,17'd4,17'd5,17'd5,17'd23,17'd23,17'd25,17'd808,17'd283,17'd1412,17'd14,17'd2781,17'd2935,17'd3427,17'd3592,17'd3427,17'd3101,17'd3252,17'd1831,17'd3250,17'd3250,17'd2784,17'd3593,17'd3429,17'd2596,17'd1415,17'd16,17'd17,17'd17,17'd16,17'd0,17'd0,17'd0,17'd2,17'd2,17'd466,17'd466,17'd2,17'd12,17'd3,17'd19,17'd19,17'd10,17'd10,17'd21,17'd25,17'd23,17'd4,17'd5,17'd5,17'd3594,17'd3594,17'd24,17'd5,17'd5,17'd5,17'd4,17'd4,17'd25,17'd25,17'd25,17'd21,17'd26,17'd26,17'd27,17'd27,17'd28,17'd28,17'd288,17'd289,17'd30,17'd1129,17'd1129,17'd1129,17'd3256,17'd3254,17'd3254,17'd2940,17'd2940,17'd2940,17'd2941,17'd3255,17'd3255,17'd3595,17'd3433,17'd3433,17'd3595,17'd3595,17'd3433,17'd3433,17'd3595,17'd3595,17'd3434,17'd3435,17'd3258,17'd3596,17'd1975,17'd1974,17'd2431,17'd2431,17'd2607,17'd2607,17'd3597,17'd3261,17'd2608,17'd3261,17'd2948,17'd2948,17'd3597,17'd2608,17'd3598,17'd3599,17'd1425,17'd2949,17'd2949,17'd2949,17'd3108,17'd1708,17'd3600,17'd3601,17'd3602,17'd3602,17'd3603,17'd3604,17'd3442,17'd3443,17'd3605,17'd3606,17'd3607,17'd3608,17'd3609,17'd3610,17'd2628,17'd3276,17'd3611,17'd3612,17'd3613,17'd3281,17'd3614,17'd3615,17'd3616,17'd3617,17'd3618,17'd3619,17'd3460,17'd3620,17'd3621,17'd3622,17'd3464,17'd3623,17'd3465,17'd3624,17'd3296,17'd3625,17'd3470,17'd3471,17'd3471,17'd3472,17'd3626,17'd3627,17'd3628,17'd3629,17'd3630,17'd3631,17'd3632,17'd3633,17'd3634,17'd3477,17'd3635,17'd3636,17'd2466,17'd3481,17'd3637,17'd3638,17'd2300,17'd3486,17'd3639,17'd3309,17'd3640,17'd2017,17'd2021,17'd2998,17'd3641,17'd2663,17'd3642,17'd3643,17'd3495,17'd3644,17'd3496,17'd2487,17'd3645,17'd3646,17'd3498,17'd3647,17'd3648,17'd3649,17'd2320,17'd1752,17'd2321,17'd3650,17'd3325,17'd3326,17'd2325,17'd3651,17'd3018,17'd3652,17'd3163,17'd3653,17'd3164,17'd3654,17'd3655,17'd2183,17'd3656,17'd883,17'd884,17'd535,17'd1475,17'd1758,17'd1334,17'd1334,17'd1475,17'd1475,17'd3657,17'd1612,17'd2340,17'd3658,17'd541,17'd1481,17'd1481,17'd1481,17'd133,17'd1197,17'd1197,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd1197,17'd133,17'd132,17'd132,17'd131,17'd357,17'd2862,17'd3659,17'd3028,17'd3660,17'd3661,17'd3662,17'd3663,17'd3664,17'd3665,17'd3666,17'd3667,17'd3668,17'd3669,17'd3670,17'd3671,17'd3672,17'd3673,17'd3674,17'd3675,17'd3676,17'd3677,17'd3678,17'd3679,17'd3680,17'd3681,17'd3682,17'd3683,17'd3684,17'd3685,17'd3686,17'd3687,17'd3688,17'd3688,17'd3689,17'd3690,17'd3691,17'd3692,17'd3369,17'd3548,17'd3549,17'd3693,17'd3694,17'd3695,17'd3696,17'd3696,17'd3696,17'd3697,17'd3554,17'd3552,17'd3698,17'd3699,17'd3700,17'd3701,17'd3560,17'd3702,17'd3703,17'd3704,17'd3705,17'd3706,17'd3707,17'd3708,17'd3709,17'd3710,17'd3568,17'd3711,17'd3072,17'd1810,17'd3712,17'd3713,17'd3714,17'd3715,17'd3716,17'd3399,17'd3398,17'd3717,17'd3717,17'd3398,17'd3399,17'd3402,17'd3575,17'd3718,17'd3402,17'd3403,17'd3230,17'd2753,17'd3719,17'd3082,17'd3082,17'd3720,17'd3721,17'd3576,17'd3722,17'd3723,17'd3724,17'd3724,17'd3725,17'd3726,17'd3727,17'd3728,17'd3729,17'd3730,17'd3582,17'd3731,17'd3732,17'd3238,17'd3733,17'd3734,17'd3735,17'd3736,17'd2926,17'd3737,17'd2771,17'd3738,17'd3738,17'd3739,17'd3739,17'd2929,17'd3740,17'd3096,17'd3741,17'd3742,17'd2417,17'd3743,17'd3743,17'd1401,17'd230,17'd1399,17'd1260,17'd1119,17'd3247,17'd3391,17'd3744,17'd3425,17'd3425,17'd3423,17'd3423,17'd3423,17'd3247,17'd1119,17'd625,17'd1824,17'd3426,17'd795,17'd795,17'd3072,17'd3745,17'd3248,17'd2587,17'd2587,17'd2587,17'd782,17'd782,17'd607,17'd607,17'd207,17'd207,17'd3746,17'd206,17'd644,17'd1963,17'd973,17'd973,17'd1550,17'd973,17'd1828,17'd3747,17'd269,17'd272,17'd273,17'd272,17'd803,17'd803,17'd971,17'd971,17'd1272,17'd952,17'd1245,17'd2116
},
'{
17'd283,17'd283,17'd650,17'd283,17'd10,17'd21,17'd23,17'd4,17'd5,17'd5,17'd23,17'd25,17'd808,17'd3748,17'd283,17'd3749,17'd3750,17'd2592,17'd3751,17'd3592,17'd3592,17'd3427,17'd2935,17'd2422,17'd1831,17'd2422,17'd2784,17'd2935,17'd3593,17'd3752,17'd2596,17'd1415,17'd16,17'd17,17'd17,17'd16,17'd0,17'd0,17'd0,17'd2,17'd466,17'd466,17'd466,17'd2,17'd12,17'd3,17'd19,17'd19,17'd10,17'd10,17'd25,17'd25,17'd23,17'd23,17'd5,17'd5,17'd3753,17'd3594,17'd5,17'd5,17'd5,17'd5,17'd4,17'd23,17'd25,17'd25,17'd25,17'd21,17'd26,17'd26,17'd27,17'd286,17'd287,17'd28,17'd289,17'd468,17'd290,17'd1129,17'd1129,17'd31,17'd3256,17'd3254,17'd3254,17'd3256,17'd3256,17'd3254,17'd3255,17'd3754,17'd3755,17'd3595,17'd3433,17'd3433,17'd3433,17'd3595,17'd3433,17'd3433,17'd3755,17'd3755,17'd3756,17'd3435,17'd3105,17'd2264,17'd1975,17'd1974,17'd2431,17'd2431,17'd2607,17'd2607,17'd3597,17'd3597,17'd3757,17'd3261,17'd3597,17'd3597,17'd3757,17'd2268,17'd1707,17'd1560,17'd1425,17'd1141,17'd1141,17'd1425,17'd1708,17'd2435,17'd2609,17'd3758,17'd3759,17'd3759,17'd3760,17'd3761,17'd3762,17'd3763,17'd3764,17'd2800,17'd3765,17'd3766,17'd3767,17'd3768,17'd3769,17'd3770,17'd3771,17'd3772,17'd3773,17'd3455,17'd3774,17'd3775,17'd3617,17'd3776,17'd3459,17'd3460,17'd3777,17'd3778,17'd3779,17'd3464,17'd3623,17'd3623,17'd3138,17'd3138,17'd3471,17'd3780,17'd3781,17'd3627,17'd3473,17'd3473,17'd3782,17'd3783,17'd3784,17'd3785,17'd3786,17'd3785,17'd3631,17'd3787,17'd3788,17'd3789,17'd3790,17'd3791,17'd2465,17'd2467,17'd3637,17'd3638,17'd2300,17'd3308,17'd2303,17'd2828,17'd3792,17'd3793,17'd3794,17'd2999,17'd3001,17'd3795,17'd2665,17'd3796,17'd1747,17'd3797,17'd3798,17'd2169,17'd2488,17'd3799,17'd3321,17'd2029,17'd3159,17'd1602,17'd2171,17'd3160,17'd3800,17'd3801,17'd3801,17'd3802,17'd3503,17'd2850,17'd3803,17'd3804,17'd3805,17'd3806,17'd3807,17'd3808,17'd3809,17'd3810,17'd1756,17'd1757,17'd3022,17'd3022,17'd711,17'd2337,17'd884,17'd711,17'd1610,17'd535,17'd2339,17'd3333,17'd1479,17'd2040,17'd1481,17'd1481,17'd1481,17'd1481,17'd1197,17'd1197,17'd542,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd132,17'd132,17'd357,17'd3811,17'd3812,17'd3813,17'd3814,17'd3815,17'd3816,17'd3817,17'd3818,17'd3819,17'd3820,17'd3821,17'd3822,17'd3823,17'd3824,17'd3825,17'd3826,17'd3827,17'd3828,17'd3829,17'd3830,17'd3831,17'd3832,17'd3833,17'd3834,17'd3835,17'd3836,17'd3837,17'd3838,17'd3839,17'd3840,17'd3841,17'd3842,17'd3843,17'd3844,17'd3845,17'd3846,17'd3847,17'd3848,17'd3849,17'd3850,17'd3851,17'd3852,17'd3853,17'd3854,17'd3855,17'd3856,17'd3857,17'd3857,17'd3858,17'd3859,17'd3860,17'd3861,17'd3862,17'd3863,17'd3864,17'd3865,17'd3702,17'd3866,17'd3867,17'd3868,17'd3869,17'd3869,17'd3870,17'd3871,17'd3872,17'd3872,17'd3873,17'd3874,17'd1824,17'd3391,17'd3875,17'd3713,17'd3714,17'd1953,17'd3876,17'd3401,17'd3401,17'd3717,17'd3877,17'd3574,17'd3575,17'd3575,17'd3878,17'd3878,17'd3402,17'd3879,17'd2753,17'd2915,17'd3082,17'd3082,17'd3720,17'd3721,17'd3722,17'd3880,17'd3881,17'd3725,17'd3724,17'd3725,17'd3882,17'd3883,17'd3884,17'd3728,17'd3581,17'd3885,17'd3886,17'd3887,17'd3888,17'd3413,17'd3889,17'd3586,17'd2767,17'd2926,17'd3417,17'd3737,17'd3739,17'd3419,17'd3890,17'd3891,17'd3892,17'd2772,17'd3416,17'd3893,17'd3894,17'd2559,17'd1823,17'd3743,17'd1261,17'd230,17'd1399,17'd1399,17'd1119,17'd3247,17'd3895,17'd3744,17'd3896,17'd3896,17'd3423,17'd3423,17'd3423,17'd3897,17'd3247,17'd2586,17'd3898,17'd1825,17'd1264,17'd1264,17'd3072,17'd3745,17'd3248,17'd3248,17'd3248,17'd2587,17'd782,17'd782,17'd607,17'd1679,17'd607,17'd258,17'd3899,17'd2779,17'd644,17'd1963,17'd973,17'd1410,17'd1550,17'd3900,17'd1410,17'd1829,17'd269,17'd273,17'd274,17'd272,17'd803,17'd803,17'd971,17'd971,17'd1272,17'd1272,17'd1245,17'd2116
},
'{
17'd806,17'd1275,17'd1275,17'd1275,17'd25,17'd25,17'd23,17'd24,17'd24,17'd24,17'd23,17'd9,17'd651,17'd283,17'd2,17'd1688,17'd2784,17'd3901,17'd3902,17'd3902,17'd3903,17'd3904,17'd2935,17'd3252,17'd2422,17'd2422,17'd2935,17'd2593,17'd3593,17'd3752,17'd1414,17'd17,17'd3905,17'd18,17'd0,17'd1,17'd1,17'd0,17'd2,17'd466,17'd2595,17'd2595,17'd466,17'd466,17'd3905,17'd18,17'd979,17'd979,17'd10,17'd21,17'd25,17'd25,17'd23,17'd4,17'd5,17'd5,17'd3594,17'd3594,17'd5,17'd6,17'd6,17'd6,17'd4,17'd23,17'd9,17'd25,17'd21,17'd20,17'd3906,17'd26,17'd286,17'd1833,17'd652,17'd652,17'd289,17'd468,17'd30,17'd30,17'd30,17'd30,17'd3433,17'd3433,17'd3433,17'd3433,17'd3595,17'd3755,17'd3907,17'd3907,17'd3908,17'd3908,17'd3909,17'd3909,17'd3908,17'd3908,17'd3755,17'd3755,17'd3910,17'd3910,17'd3434,17'd3104,17'd2604,17'd2946,17'd2606,17'd2606,17'd3911,17'd2948,17'd2948,17'd2948,17'd3912,17'd3912,17'd3913,17'd3913,17'd3913,17'd3914,17'd3915,17'd3598,17'd3916,17'd3108,17'd1425,17'd1425,17'd1560,17'd1707,17'd3917,17'd3918,17'd3919,17'd3920,17'd3921,17'd3922,17'd3923,17'd3924,17'd3925,17'd3926,17'd3927,17'd2625,17'd3928,17'd3929,17'd3768,17'd3930,17'd3931,17'd3932,17'd3933,17'd3934,17'd3935,17'd3936,17'd3937,17'd3938,17'd3939,17'd3940,17'd3941,17'd3942,17'd3943,17'd3944,17'd3944,17'd3945,17'd3945,17'd3945,17'd3945,17'd3946,17'd3946,17'd3473,17'd3947,17'd3948,17'd3949,17'd3950,17'd3950,17'd3951,17'd3951,17'd3952,17'd3953,17'd3954,17'd3955,17'd3632,17'd3956,17'd3957,17'd3302,17'd3958,17'd3959,17'd3960,17'd3638,17'd3961,17'd2301,17'd2302,17'd2303,17'd3962,17'd3963,17'd3964,17'd2998,17'd3641,17'd3965,17'd3966,17'd3967,17'd3968,17'd3969,17'd2486,17'd3970,17'd3971,17'd3972,17'd3972,17'd3973,17'd3973,17'd3974,17'd3975,17'd3976,17'd2679,17'd3977,17'd3978,17'd3978,17'd3979,17'd3980,17'd3981,17'd3982,17'd3983,17'd3984,17'd3985,17'd3986,17'd3987,17'd3988,17'd3989,17'd3990,17'd3991,17'd3992,17'd3993,17'd1894,17'd1756,17'd3994,17'd2184,17'd884,17'd1334,17'd537,17'd1477,17'd1613,17'd3995,17'd356,17'd356,17'd356,17'd356,17'd719,17'd719,17'd719,17'd719,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd2698,17'd131,17'd3996,17'd3170,17'd3997,17'd3998,17'd3999,17'd4000,17'd4001,17'd4002,17'd4003,17'd4004,17'd4005,17'd4006,17'd4007,17'd4008,17'd4009,17'd4010,17'd4011,17'd4012,17'd4013,17'd4014,17'd4015,17'd4016,17'd4017,17'd4018,17'd4019,17'd4020,17'd4021,17'd4022,17'd4023,17'd4024,17'd4025,17'd4026,17'd4027,17'd4028,17'd4029,17'd4030,17'd4031,17'd4032,17'd4033,17'd4034,17'd4035,17'd4036,17'd4037,17'd4038,17'd4039,17'd4040,17'd4041,17'd4042,17'd4043,17'd4044,17'd4045,17'd4046,17'd4047,17'd4048,17'd3860,17'd4049,17'd4050,17'd4051,17'd4052,17'd3866,17'd4053,17'd4054,17'd4055,17'd4056,17'd3709,17'd4057,17'd4057,17'd4058,17'd2390,17'd4059,17'd1260,17'd2096,17'd4060,17'd4061,17'd2407,17'd2750,17'd3081,17'd3399,17'd3398,17'd3398,17'd3574,17'd4062,17'd4062,17'd4063,17'd4064,17'd4065,17'd4066,17'd1817,17'd3719,17'd4067,17'd4068,17'd4069,17'd4070,17'd4071,17'd3576,17'd3576,17'd3722,17'd3724,17'd3725,17'd4072,17'd4073,17'd3232,17'd3884,17'd3728,17'd3728,17'd4074,17'd4075,17'd3886,17'd4076,17'd4077,17'd4078,17'd3241,17'd3736,17'd4079,17'd4079,17'd4080,17'd3739,17'd4081,17'd4081,17'd4082,17'd4083,17'd2768,17'd3241,17'd3734,17'd3894,17'd4084,17'd1823,17'd1401,17'd445,17'd1401,17'd3098,17'd1399,17'd1119,17'd4085,17'd4085,17'd3391,17'd3391,17'd4085,17'd4085,17'd3423,17'd3423,17'd2096,17'd2096,17'd2777,17'd625,17'd443,17'd232,17'd795,17'd3072,17'd1402,17'd3072,17'd3072,17'd1402,17'd623,17'd443,17'd443,17'd427,17'd954,17'd259,17'd260,17'd3899,17'd2779,17'd803,17'd1963,17'd1963,17'd1098,17'd1098,17'd973,17'd1687,17'd206,17'd643,17'd273,17'd273,17'd644,17'd803,17'd971,17'd971,17'd1272,17'd1272,17'd1245,17'd2116
},
'{
17'd806,17'd1275,17'd1275,17'd465,17'd25,17'd25,17'd23,17'd24,17'd24,17'd23,17'd23,17'd25,17'd650,17'd1,17'd14,17'd3250,17'd2934,17'd4086,17'd4087,17'd4087,17'd3903,17'd4088,17'd2935,17'd2935,17'd2935,17'd2935,17'd2593,17'd2593,17'd3593,17'd3752,17'd1415,17'd17,17'd4089,17'd3905,17'd0,17'd1,17'd0,17'd2,17'd466,17'd466,17'd466,17'd466,17'd466,17'd2,17'd18,17'd18,17'd19,17'd10,17'd21,17'd21,17'd25,17'd25,17'd23,17'd4,17'd5,17'd5,17'd3594,17'd3594,17'd5,17'd6,17'd6,17'd6,17'd4,17'd23,17'd25,17'd21,17'd20,17'd20,17'd285,17'd285,17'd286,17'd286,17'd652,17'd653,17'd289,17'd289,17'd809,17'd30,17'd30,17'd30,17'd3433,17'd3433,17'd3595,17'd3755,17'd3755,17'd3907,17'd3755,17'd3755,17'd3908,17'd3908,17'd4090,17'd4090,17'd3908,17'd4091,17'd3755,17'd3755,17'd3910,17'd3434,17'd3104,17'd3105,17'd2946,17'd2946,17'd2606,17'd2606,17'd2948,17'd2948,17'd2948,17'd2948,17'd3912,17'd4092,17'd3913,17'd3913,17'd4093,17'd3915,17'd3598,17'd3598,17'd3916,17'd1708,17'd2610,17'd1707,17'd4094,17'd2786,17'd4095,17'd4096,17'd4097,17'd3922,17'd3923,17'd4098,17'd4099,17'd4100,17'd4101,17'd4102,17'd4103,17'd4104,17'd4105,17'd4106,17'd4107,17'd4108,17'd4109,17'd4110,17'd4111,17'd4112,17'd4113,17'd4114,17'd3938,17'd4115,17'd4116,17'd3941,17'd4117,17'd4118,17'd4119,17'd4120,17'd4121,17'd4121,17'd3945,17'd3946,17'd3946,17'd3627,17'd3627,17'd3628,17'd4122,17'd4123,17'd4124,17'd4125,17'd4126,17'd4126,17'd4127,17'd3952,17'd3953,17'd3954,17'd4123,17'd4128,17'd3947,17'd3301,17'd3141,17'd4129,17'd2990,17'd4130,17'd3961,17'd2301,17'd2302,17'd2659,17'd2305,17'd4131,17'd3964,17'd2163,17'd3491,17'd4132,17'd4133,17'd4134,17'd4135,17'd2840,17'd4136,17'd3969,17'd4137,17'd2671,17'd4138,17'd4138,17'd4139,17'd2676,17'd4140,17'd4140,17'd4141,17'd4142,17'd4143,17'd4144,17'd4145,17'd4146,17'd4147,17'd4148,17'd4149,17'd4150,17'd4151,17'd4152,17'd4153,17'd4154,17'd4154,17'd4155,17'd4156,17'd4157,17'd4158,17'd3992,17'd4159,17'd4160,17'd4161,17'd2694,17'd4162,17'd2338,17'd536,17'd1477,17'd1613,17'd3995,17'd1196,17'd1196,17'd4163,17'd4163,17'd3025,17'd3025,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd4164,17'd4165,17'd4166,17'd4167,17'd4168,17'd4169,17'd4170,17'd4171,17'd4172,17'd4173,17'd4174,17'd4175,17'd4176,17'd4177,17'd4178,17'd4179,17'd4180,17'd4181,17'd4182,17'd4183,17'd4184,17'd4185,17'd4186,17'd4187,17'd4188,17'd4189,17'd4190,17'd4191,17'd4192,17'd4193,17'd4194,17'd4194,17'd4195,17'd4196,17'd4197,17'd4198,17'd4199,17'd4200,17'd4201,17'd4202,17'd4203,17'd4204,17'd4205,17'd4206,17'd4207,17'd4208,17'd4209,17'd4210,17'd4211,17'd4212,17'd4213,17'd4214,17'd4215,17'd4216,17'd4217,17'd4218,17'd4219,17'd4220,17'd3698,17'd4221,17'd4222,17'd3702,17'd4223,17'd4224,17'd4225,17'd3567,17'd4226,17'd4057,17'd4057,17'd4227,17'd4228,17'd3426,17'd4229,17'd3247,17'd3712,17'd4230,17'd4231,17'd2751,17'd3876,17'd3400,17'd3398,17'd3574,17'd4232,17'd4232,17'd4063,17'd4063,17'd4232,17'd4233,17'd3575,17'd3403,17'd3719,17'd4067,17'd3082,17'd4069,17'd3406,17'd3576,17'd3576,17'd3576,17'd3881,17'd3724,17'd4072,17'd4073,17'd4234,17'd3083,17'd3884,17'd3729,17'd3885,17'd3885,17'd3887,17'd3886,17'd4235,17'd4236,17'd4237,17'd4238,17'd3589,17'd3243,17'd3740,17'd4080,17'd3891,17'd4239,17'd4082,17'd4240,17'd3740,17'd2926,17'd4238,17'd3734,17'd4241,17'd4084,17'd1680,17'd1261,17'd1261,17'd230,17'd1260,17'd228,17'd3895,17'd3391,17'd4085,17'd4085,17'd4085,17'd3391,17'd3897,17'd3897,17'd2096,17'd2096,17'd3247,17'd624,17'd446,17'd443,17'd795,17'd795,17'd1402,17'd3072,17'd3072,17'd3072,17'd626,17'd623,17'd443,17'd443,17'd954,17'd954,17'd260,17'd426,17'd426,17'd644,17'd645,17'd645,17'd1685,17'd1098,17'd973,17'd1687,17'd643,17'd643,17'd273,17'd273,17'd644,17'd803,17'd971,17'd971,17'd1272,17'd1272,17'd1245,17'd2116
},
'{
17'd1275,17'd806,17'd1275,17'd465,17'd977,17'd977,17'd4,17'd23,17'd2421,17'd4242,17'd2591,17'd1275,17'd1,17'd15,17'd1688,17'd2935,17'd4243,17'd4087,17'd4087,17'd4087,17'd4244,17'd4088,17'd4245,17'd4246,17'd2935,17'd2934,17'd2934,17'd2593,17'd2592,17'd1689,17'd1415,17'd17,17'd466,17'd2,17'd0,17'd0,17'd14,17'd1127,17'd1127,17'd4247,17'd466,17'd2,17'd2,17'd0,17'd18,17'd19,17'd11,17'd11,17'd25,17'd25,17'd23,17'd23,17'd24,17'd5,17'd3594,17'd3753,17'd3753,17'd3753,17'd5,17'd5,17'd5,17'd5,17'd23,17'd22,17'd21,17'd20,17'd20,17'd21,17'd1833,17'd1833,17'd286,17'd980,17'd653,17'd653,17'd289,17'd289,17'd289,17'd289,17'd468,17'd1692,17'd3908,17'd3908,17'd289,17'd29,17'd29,17'd29,17'd289,17'd468,17'd653,17'd653,17'd4248,17'd4248,17'd4091,17'd4091,17'd3755,17'd3755,17'd3434,17'd4249,17'd4250,17'd4251,17'd2604,17'd2946,17'd2605,17'd2605,17'd4252,17'd4252,17'd4253,17'd4253,17'd4092,17'd4254,17'd4254,17'd4255,17'd3914,17'd4256,17'd4257,17'd4257,17'd4258,17'd4095,17'd4259,17'd4259,17'd4259,17'd3915,17'd4260,17'd4261,17'd4262,17'd4263,17'd4098,17'd4264,17'd4265,17'd4266,17'd4267,17'd4268,17'd4269,17'd4270,17'd4271,17'd4272,17'd4273,17'd4109,17'd4274,17'd4275,17'd4276,17'd4277,17'd4278,17'd4279,17'd4280,17'd4281,17'd4282,17'd4283,17'd4117,17'd4284,17'd4119,17'd4285,17'd4286,17'd4287,17'd3779,17'd4288,17'd4289,17'd4122,17'd4290,17'd3950,17'd4291,17'd4291,17'd4291,17'd4291,17'd4291,17'd4291,17'd4127,17'd4127,17'd4292,17'd3954,17'd3955,17'd4293,17'd3475,17'd4294,17'd4295,17'd4296,17'd4297,17'd4298,17'd4299,17'd4300,17'd4301,17'd2659,17'd4302,17'd4303,17'd3964,17'd2479,17'd4304,17'd2834,17'd2665,17'd2166,17'd4305,17'd4306,17'd4307,17'd4307,17'd4308,17'd4308,17'd4309,17'd4310,17'd4311,17'd4312,17'd4313,17'd4140,17'd2846,17'd4314,17'd4315,17'd4316,17'd4317,17'd4318,17'd3802,17'd4319,17'd4320,17'd4321,17'd4322,17'd4323,17'd4324,17'd4325,17'd4326,17'd3993,17'd4327,17'd4328,17'd4329,17'd4330,17'd4331,17'd4332,17'd4333,17'd4334,17'd2338,17'd1194,17'd2186,17'd713,17'd713,17'd2037,17'd3511,17'd3337,17'd4335,17'd4163,17'd3025,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd135,17'd4336,17'd4337,17'd4338,17'd4339,17'd4340,17'd4341,17'd4342,17'd4343,17'd4344,17'd4345,17'd4346,17'd4347,17'd4348,17'd4349,17'd4350,17'd4351,17'd4352,17'd4353,17'd4354,17'd4015,17'd4355,17'd4016,17'd4356,17'd4357,17'd4358,17'd4359,17'd4360,17'd4361,17'd4362,17'd4363,17'd4364,17'd4363,17'd4365,17'd4366,17'd4367,17'd4368,17'd4369,17'd4370,17'd4370,17'd4371,17'd4371,17'd4372,17'd4373,17'd4374,17'd4375,17'd4375,17'd4376,17'd4377,17'd4378,17'd4379,17'd4380,17'd4381,17'd4382,17'd4383,17'd4384,17'd4385,17'd4386,17'd4387,17'd3856,17'd4388,17'd4389,17'd4390,17'd4391,17'd4392,17'd3562,17'd4393,17'd4394,17'd3567,17'd4057,17'd4395,17'd4396,17'd4397,17'd4398,17'd4399,17'd4400,17'd4085,17'd4401,17'd4402,17'd2407,17'd2750,17'd3876,17'd3397,17'd4403,17'd4404,17'd4232,17'd4405,17'd4406,17'd4062,17'd4407,17'd4062,17'd3575,17'd3719,17'd3719,17'd4408,17'd4067,17'd4409,17'd3720,17'd3405,17'd4410,17'd4410,17'd3406,17'd4411,17'd4412,17'd4413,17'd4234,17'd3083,17'd3884,17'd3728,17'd3729,17'd4074,17'd4414,17'd3727,17'd3732,17'd4415,17'd4416,17'd4238,17'd3736,17'd3243,17'd4417,17'd4418,17'd4419,17'd3892,17'd4240,17'd4080,17'd3736,17'd4238,17'd4420,17'd4421,17'd4241,17'd2775,17'd1680,17'd1261,17'd1261,17'd1401,17'd3098,17'd1401,17'd445,17'd1810,17'd4422,17'd4085,17'd4085,17'd4085,17'd4423,17'd3897,17'd2096,17'd2096,17'd4424,17'd624,17'd446,17'd231,17'd1544,17'd1402,17'd1402,17'd3072,17'd3072,17'd3072,17'd3072,17'd623,17'd443,17'd427,17'd954,17'd954,17'd260,17'd426,17'd259,17'd644,17'd803,17'd1685,17'd1098,17'd1550,17'd1410,17'd644,17'd643,17'd643,17'd643,17'd644,17'd803,17'd971,17'd1685,17'd1244,17'd1244,17'd1382,17'd422
},
'{
17'd1275,17'd806,17'd1275,17'd465,17'd651,17'd807,17'd9,17'd23,17'd978,17'd977,17'd1275,17'd3,17'd15,17'd1689,17'd2422,17'd2934,17'd4425,17'd4426,17'd4087,17'd4427,17'd3903,17'd4428,17'd4088,17'd4088,17'd3751,17'd2934,17'd2934,17'd2935,17'd3250,17'd1967,17'd1415,17'd17,17'd2,17'd0,17'd0,17'd0,17'd1127,17'd1127,17'd1127,17'd1127,17'd2,17'd2,17'd2,17'd0,17'd19,17'd19,17'd11,17'd11,17'd25,17'd25,17'd23,17'd23,17'd24,17'd5,17'd3753,17'd3753,17'd3753,17'd3753,17'd6,17'd5,17'd5,17'd24,17'd23,17'd22,17'd20,17'd20,17'd21,17'd25,17'd4429,17'd1833,17'd27,17'd1278,17'd653,17'd653,17'd289,17'd289,17'd289,17'd289,17'd468,17'd468,17'd4091,17'd4091,17'd289,17'd29,17'd29,17'd29,17'd289,17'd468,17'd653,17'd653,17'd4430,17'd4430,17'd4431,17'd4091,17'd3755,17'd3255,17'd4249,17'd3104,17'd4251,17'd2604,17'd2604,17'd2946,17'd2605,17'd2605,17'd4252,17'd4253,17'd4253,17'd4432,17'd4254,17'd4254,17'd4254,17'd3913,17'd4433,17'd4434,17'd4257,17'd4257,17'd4095,17'd4260,17'd4435,17'd4435,17'd4433,17'd4436,17'd4437,17'd4438,17'd4439,17'd4098,17'd4099,17'd4265,17'd4266,17'd4440,17'd4441,17'd4442,17'd4443,17'd4444,17'd4445,17'd4446,17'd4447,17'd4448,17'd4449,17'd4450,17'd4451,17'd4452,17'd4453,17'd4454,17'd4455,17'd4456,17'd4283,17'd4457,17'd4458,17'd4459,17'd4287,17'd4287,17'd4460,17'd4460,17'd4461,17'd4462,17'd4122,17'd3950,17'd4463,17'd4126,17'd4464,17'd4464,17'd4291,17'd4291,17'd4291,17'd4291,17'd3952,17'd4292,17'd4292,17'd4123,17'd4293,17'd3474,17'd4465,17'd4466,17'd4467,17'd2981,17'd4468,17'd2827,17'd4469,17'd2470,17'd2658,17'd2305,17'd2161,17'd4470,17'd4471,17'd4472,17'd4473,17'd4474,17'd2165,17'd2026,17'd1885,17'd1885,17'd4475,17'd4476,17'd4477,17'd4478,17'd4479,17'd3319,17'd4480,17'd4481,17'd4482,17'd4483,17'd4484,17'd4485,17'd4486,17'd4487,17'd2685,17'd4488,17'd4320,17'd4321,17'd4322,17'd3988,17'd2504,17'd2689,17'd4159,17'd4489,17'd4490,17'd4490,17'd4491,17'd4492,17'd4493,17'd2184,17'd711,17'd3024,17'd2338,17'd712,17'd1194,17'd2186,17'd4494,17'd4494,17'd2697,17'd2858,17'd4495,17'd3336,17'd1196,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd3169,17'd4496,17'd4497,17'd4498,17'd4499,17'd4500,17'd4501,17'd4502,17'd4503,17'd4504,17'd4505,17'd4506,17'd4507,17'd4508,17'd4509,17'd4352,17'd4510,17'd4511,17'd4512,17'd4513,17'd4514,17'd4357,17'd4515,17'd4367,17'd4516,17'd4517,17'd4360,17'd4518,17'd4519,17'd4520,17'd4521,17'd4520,17'd4522,17'd4523,17'd4524,17'd4525,17'd4526,17'd4527,17'd4528,17'd4529,17'd4529,17'd4530,17'd4531,17'd4532,17'd4533,17'd4534,17'd4535,17'd4536,17'd4537,17'd4538,17'd4539,17'd4540,17'd4541,17'd4542,17'd4543,17'd4544,17'd4545,17'd4546,17'd4546,17'd4547,17'd4548,17'd4388,17'd4549,17'd4550,17'd4551,17'd4552,17'd4054,17'd4394,17'd3872,17'd4553,17'd4554,17'd4555,17'd4556,17'd4557,17'd4558,17'd3099,17'd4085,17'd4559,17'd4560,17'd4561,17'd2914,17'd3396,17'd3573,17'd4404,17'd4232,17'd4406,17'd4562,17'd4407,17'd4062,17'd4062,17'd4062,17'd4232,17'd3402,17'd3403,17'd4064,17'd4563,17'd4564,17'd4564,17'd4410,17'd4565,17'd4410,17'd3726,17'd4566,17'd4234,17'd4567,17'd4568,17'd2757,17'd3579,17'd3409,17'd4075,17'd4075,17'd3727,17'd3727,17'd4569,17'd4415,17'd4237,17'd4238,17'd4570,17'd3243,17'd4571,17'd4572,17'd4572,17'd3892,17'd4080,17'd3737,17'd2926,17'd4573,17'd4574,17'd3734,17'd3586,17'd2775,17'd1680,17'd445,17'd1261,17'd3098,17'd230,17'd1261,17'd2392,17'd1810,17'd4423,17'd4423,17'd4423,17'd4423,17'd4575,17'd3897,17'd3897,17'd2096,17'd3247,17'd624,17'd446,17'd1544,17'd795,17'd795,17'd1402,17'd3072,17'd3745,17'd3072,17'd623,17'd623,17'd427,17'd954,17'd953,17'd954,17'd260,17'd260,17'd643,17'd644,17'd971,17'd1685,17'd1550,17'd973,17'd803,17'd644,17'd643,17'd643,17'd803,17'd645,17'd1685,17'd1685,17'd1244,17'd1381,17'd202,17'd1382
},
'{
17'd3,17'd3,17'd283,17'd465,17'd651,17'd807,17'd977,17'd2591,17'd977,17'd465,17'd283,17'd0,17'd4576,17'd4577,17'd4245,17'd4244,17'd4578,17'd4426,17'd4087,17'd3903,17'd4428,17'd4428,17'd4088,17'd4088,17'd3901,17'd3751,17'd2934,17'd2784,17'd1689,17'd14,17'd2,17'd2,17'd0,17'd0,17'd0,17'd466,17'd4247,17'd4247,17'd1127,17'd15,17'd1127,17'd14,17'd2,17'd0,17'd19,17'd10,17'd21,17'd21,17'd23,17'd23,17'd23,17'd23,17'd5,17'd5,17'd3753,17'd3753,17'd3753,17'd3753,17'd6,17'd5,17'd4,17'd23,17'd23,17'd22,17'd20,17'd21,17'd9,17'd9,17'd1833,17'd27,17'd980,17'd980,17'd652,17'd652,17'd653,17'd2938,17'd2938,17'd653,17'd653,17'd652,17'd28,17'd652,17'd652,17'd653,17'd652,17'd652,17'd653,17'd653,17'd652,17'd652,17'd4430,17'd4430,17'd4431,17'd4091,17'd3910,17'd3434,17'd4579,17'd4250,17'd4251,17'd2604,17'd4580,17'd4580,17'd4580,17'd4580,17'd4581,17'd4581,17'd4581,17'd4581,17'd4432,17'd4432,17'd3911,17'd4092,17'd4582,17'd4583,17'd4583,17'd4433,17'd3915,17'd4093,17'd4093,17'd4584,17'd4585,17'd4586,17'd4587,17'd4588,17'd4098,17'd4099,17'd4265,17'd4589,17'd4440,17'd4590,17'd4442,17'd4591,17'd4592,17'd4593,17'd4594,17'd4595,17'd4596,17'd4597,17'd4598,17'd4451,17'd4599,17'd4600,17'd4601,17'd4602,17'd4456,17'd4603,17'd4604,17'd4605,17'd4606,17'd4607,17'd4608,17'd4288,17'd4609,17'd4609,17'd4122,17'd4123,17'd3951,17'd4291,17'd4291,17'd4610,17'd4464,17'd4611,17'd4464,17'd4464,17'd4291,17'd4291,17'd4291,17'd4291,17'd3951,17'd3955,17'd4612,17'd4613,17'd4465,17'd4614,17'd4295,17'd2981,17'd4615,17'd2827,17'd4616,17'd2469,17'd4617,17'd2659,17'd2476,17'd4618,17'd3964,17'd3794,17'd2661,17'd2164,17'd4619,17'd4620,17'd4621,17'd4622,17'd4622,17'd4623,17'd4624,17'd4625,17'd3008,17'd4626,17'd4627,17'd4628,17'd4629,17'd4630,17'd4631,17'd4632,17'd4633,17'd4634,17'd4319,17'd4635,17'd4636,17'd4637,17'd4638,17'd4639,17'd3990,17'd4640,17'd4641,17'd4642,17'd4490,17'd4643,17'd4644,17'd4645,17'd4646,17'd4493,17'd4647,17'd2510,17'd2338,17'd4648,17'd4648,17'd4649,17'd4650,17'd4651,17'd4652,17'd4653,17'd3511,17'd3337,17'd541,17'd1480,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd135,17'd3169,17'd2865,17'd4654,17'd4655,17'd4656,17'd4657,17'd4658,17'd4659,17'd4660,17'd4661,17'd4662,17'd4663,17'd4664,17'd4665,17'd4666,17'd4667,17'd4668,17'd4669,17'd4670,17'd4671,17'd4672,17'd4364,17'd4366,17'd4673,17'd4674,17'd4675,17'd4517,17'd4360,17'd4676,17'd4523,17'd4677,17'd4678,17'd4679,17'd4680,17'd4681,17'd4682,17'd4683,17'd4684,17'd4685,17'd4686,17'd4686,17'd4687,17'd4688,17'd4529,17'd4689,17'd4690,17'd4690,17'd4691,17'd4692,17'd4693,17'd4694,17'd4695,17'd4696,17'd4539,17'd4697,17'd4698,17'd4699,17'd4700,17'd4701,17'd4702,17'd4703,17'd4547,17'd4704,17'd4705,17'd3554,17'd4706,17'd4707,17'd4393,17'd4708,17'd4709,17'd4710,17'd4396,17'd4555,17'd4711,17'd4557,17'd4712,17'd3246,17'd4713,17'd4714,17'd3392,17'd3393,17'd4715,17'd4716,17'd3575,17'd4232,17'd4407,17'd4717,17'd4718,17'd4719,17'd4062,17'd4407,17'd4407,17'd4404,17'd3402,17'd3402,17'd3575,17'd4064,17'd4720,17'd3082,17'd2405,17'd2405,17'd4410,17'd3405,17'd3406,17'd3578,17'd4567,17'd4721,17'd3084,17'd3884,17'd3579,17'd3409,17'd3886,17'd3727,17'd4722,17'd4723,17'd4724,17'd4725,17'd4238,17'd2768,17'd3243,17'd4417,17'd4572,17'd4571,17'd3737,17'd4080,17'd3737,17'd3417,17'd4726,17'd4574,17'd3893,17'd3590,17'd2417,17'd445,17'd3743,17'd4727,17'd1401,17'd1262,17'd1261,17'd2392,17'd4423,17'd4728,17'd4713,17'd4729,17'd4730,17'd4575,17'd3897,17'd2096,17'd2096,17'd3247,17'd228,17'd227,17'd1264,17'd1264,17'd795,17'd1402,17'd3072,17'd3745,17'd446,17'd446,17'd227,17'd227,17'd953,17'd953,17'd259,17'd260,17'd260,17'd643,17'd972,17'd971,17'd1963,17'd1963,17'd645,17'd644,17'd643,17'd643,17'd644,17'd645,17'd1685,17'd1098,17'd1381,17'd1381,17'd4731,17'd4731
},
'{
17'd12,17'd3,17'd283,17'd650,17'd4732,17'd651,17'd465,17'd465,17'd465,17'd283,17'd0,17'd1967,17'd4577,17'd4733,17'd4244,17'd4426,17'd4734,17'd4735,17'd3902,17'd4244,17'd4428,17'd4428,17'd3903,17'd4736,17'd4737,17'd4738,17'd2593,17'd3250,17'd1689,17'd14,17'd2,17'd2,17'd1,17'd0,17'd2,17'd466,17'd4247,17'd1127,17'd14,17'd15,17'd1127,17'd14,17'd2,17'd12,17'd11,17'd10,17'd25,17'd25,17'd23,17'd23,17'd23,17'd4,17'd5,17'd6,17'd3753,17'd3753,17'd3753,17'd3753,17'd6,17'd5,17'd23,17'd23,17'd23,17'd23,17'd21,17'd25,17'd9,17'd25,17'd27,17'd980,17'd1278,17'd980,17'd652,17'd652,17'd653,17'd2938,17'd2938,17'd653,17'd652,17'd28,17'd287,17'd28,17'd652,17'd653,17'd653,17'd652,17'd652,17'd652,17'd652,17'd652,17'd4430,17'd4430,17'd4091,17'd3755,17'd3434,17'd3434,17'd4250,17'd4739,17'd4739,17'd2604,17'd4580,17'd4580,17'd4580,17'd4580,17'd4740,17'd4741,17'd4742,17'd4581,17'd4432,17'd4253,17'd3911,17'd2948,17'd3261,17'd4433,17'd3915,17'd4093,17'd4093,17'd4743,17'd4743,17'd4744,17'd4745,17'd4746,17'd4747,17'd4263,17'd4099,17'd4265,17'd4748,17'd4749,17'd4750,17'd4442,17'd4751,17'd4752,17'd4753,17'd4754,17'd4755,17'd4448,17'd4756,17'd4598,17'd4757,17'd4599,17'd4758,17'd4759,17'd4760,17'd4115,17'd4761,17'd4762,17'd4763,17'd4764,17'd4765,17'd4609,17'd4462,17'd3949,17'd3950,17'd3950,17'd3951,17'd4126,17'd4127,17'd4127,17'd4610,17'd4766,17'd4767,17'd4767,17'd4766,17'd4766,17'd4768,17'd4768,17'd4291,17'd4769,17'd4123,17'd4770,17'd3956,17'd3476,17'd4771,17'd3141,17'd4129,17'd4772,17'd4468,17'd2650,17'd4773,17'd4774,17'd4617,17'd4775,17'd2476,17'd2159,17'd4776,17'd2162,17'd4777,17'd4778,17'd4779,17'd4780,17'd4781,17'd4782,17'd4783,17'd4784,17'd4785,17'd4786,17'd3797,17'd4787,17'd4788,17'd4789,17'd4790,17'd4791,17'd4792,17'd4793,17'd4794,17'd4795,17'd4795,17'd4796,17'd4797,17'd4798,17'd4799,17'd4800,17'd4801,17'd4802,17'd4803,17'd4804,17'd4805,17'd4806,17'd4807,17'd4808,17'd4808,17'd4809,17'd4810,17'd4811,17'd4810,17'd4812,17'd4812,17'd4812,17'd4813,17'd4650,17'd4495,17'd3511,17'd540,17'd541,17'd1480,17'd1481,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd135,17'd131,17'd4814,17'd4815,17'd4816,17'd4817,17'd4342,17'd4818,17'd4819,17'd4820,17'd4821,17'd4822,17'd4823,17'd4178,17'd4824,17'd4825,17'd4826,17'd4827,17'd4828,17'd4829,17'd4830,17'd4831,17'd4832,17'd4018,17'd4833,17'd4834,17'd4368,17'd4835,17'd4836,17'd4836,17'd4837,17'd4838,17'd4838,17'd4837,17'd4837,17'd4681,17'd4839,17'd4840,17'd4841,17'd4842,17'd4842,17'd4843,17'd4844,17'd4844,17'd4845,17'd4687,17'd4846,17'd4846,17'd4847,17'd4846,17'd4848,17'd4849,17'd4850,17'd4851,17'd4851,17'd4852,17'd4853,17'd4854,17'd4855,17'd4856,17'd4857,17'd4858,17'd4859,17'd4214,17'd4548,17'd4860,17'd4861,17'd3554,17'd4862,17'd4863,17'd4224,17'd4708,17'd4864,17'd4227,17'd4395,17'd4865,17'd4711,17'd4866,17'd4867,17'd4868,17'd4869,17'd2906,17'd3392,17'd2574,17'd3394,17'd4870,17'd4404,17'd4062,17'd4062,17'd4718,17'd4871,17'd4872,17'd4407,17'd4873,17'd4873,17'd4403,17'd3876,17'd3396,17'd3575,17'd3575,17'd4064,17'd3082,17'd2405,17'd4565,17'd4565,17'd4410,17'd3407,17'd4234,17'd4568,17'd3232,17'd3084,17'd3579,17'd3729,17'd3887,17'd3886,17'd4722,17'd4874,17'd4875,17'd4876,17'd4877,17'd3241,17'd4079,17'd3243,17'd4878,17'd4879,17'd4417,17'd4080,17'd3737,17'd4417,17'd3417,17'd4726,17'd4574,17'd3421,17'd2585,17'd445,17'd4880,17'd4881,17'd1261,17'd1262,17'd1401,17'd445,17'd4085,17'd4882,17'd4713,17'd4729,17'd4730,17'd4883,17'd4883,17'd3897,17'd3897,17'd3247,17'd2586,17'd1119,17'd3426,17'd795,17'd795,17'd795,17'd3072,17'd3745,17'd625,17'd625,17'd446,17'd446,17'd1962,17'd1962,17'd953,17'd260,17'd260,17'd259,17'd425,17'd972,17'd1963,17'd1963,17'd645,17'd643,17'd206,17'd206,17'd644,17'd803,17'd1685,17'd1098,17'd1381,17'd1245,17'd4731,17'd2932
},
'{
17'd2,17'd1,17'd4884,17'd650,17'd650,17'd465,17'd465,17'd465,17'd806,17'd12,17'd4885,17'd4886,17'd4887,17'd4428,17'd4426,17'd4888,17'd4889,17'd4890,17'd4891,17'd4892,17'd4428,17'd3903,17'd4427,17'd4087,17'd4893,17'd4738,17'd2782,17'd2781,17'd1127,17'd2,17'd2,17'd0,17'd0,17'd2,17'd1127,17'd4247,17'd1127,17'd14,17'd14,17'd14,17'd14,17'd14,17'd2,17'd12,17'd11,17'd10,17'd25,17'd25,17'd22,17'd23,17'd4,17'd4,17'd6,17'd6,17'd3753,17'd3753,17'd5,17'd6,17'd5,17'd5,17'd23,17'd23,17'd467,17'd467,17'd9,17'd9,17'd25,17'd21,17'd980,17'd980,17'd980,17'd980,17'd652,17'd652,17'd653,17'd653,17'd1278,17'd980,17'd27,17'd27,17'd28,17'd652,17'd652,17'd652,17'd652,17'd652,17'd652,17'd652,17'd980,17'd980,17'd4430,17'd4248,17'd4091,17'd3595,17'd3434,17'd4249,17'd4250,17'd4739,17'd2604,17'd2946,17'd4580,17'd4894,17'd4740,17'd4740,17'd4895,17'd4895,17'd4740,17'd4740,17'd4581,17'd4896,17'd4253,17'd2948,17'd3913,17'd3913,17'd4255,17'd4254,17'd4743,17'd4897,17'd4898,17'd4899,17'd4900,17'd4746,17'd4901,17'd4902,17'd4265,17'd4903,17'd4904,17'd4905,17'd4906,17'd4907,17'd4752,17'd4908,17'd4909,17'd4910,17'd4911,17'd4912,17'd4913,17'd4914,17'd4915,17'd4916,17'd4917,17'd4918,17'd4602,17'd4281,17'd4919,17'd4920,17'd4763,17'd4764,17'd4921,17'd4922,17'd4463,17'd4923,17'd4924,17'd4924,17'd4610,17'd4610,17'd4925,17'd4925,17'd4925,17'd4926,17'd4927,17'd4927,17'd4925,17'd4928,17'd4768,17'd4291,17'd4125,17'd4124,17'd3631,17'd3632,17'd3956,17'd3476,17'd4771,17'd3141,17'd4129,17'd4929,17'd4930,17'd4931,17'd4932,17'd4774,17'd4617,17'd2659,17'd4302,17'd4131,17'd2161,17'd4933,17'd4934,17'd4935,17'd4936,17'd4937,17'd4938,17'd4939,17'd4783,17'd4940,17'd4941,17'd4942,17'd4943,17'd4140,17'd3976,17'd4944,17'd4945,17'd4946,17'd4794,17'd4947,17'd4948,17'd4949,17'd4950,17'd4951,17'd4952,17'd4953,17'd4954,17'd4955,17'd4956,17'd4957,17'd4958,17'd4959,17'd4960,17'd4961,17'd4962,17'd4963,17'd4964,17'd4965,17'd4965,17'd4966,17'd4967,17'd4968,17'd4969,17'd4969,17'd4970,17'd4971,17'd3336,17'd1196,17'd356,17'd1481,17'd1481,17'd1481,17'd356,17'd356,17'd356,17'd1481,17'd1197,17'd1197,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd132,17'd132,17'd134,17'd1759,17'd4972,17'd4973,17'd4815,17'd4974,17'd4975,17'd4976,17'd4977,17'd4978,17'd4979,17'd4980,17'd4981,17'd4982,17'd4983,17'd3829,17'd4984,17'd4985,17'd4986,17'd4987,17'd4988,17'd4989,17'd4521,17'd4990,17'd4991,17'd4838,17'd4992,17'd4993,17'd4994,17'd4840,17'd4995,17'd4996,17'd4997,17'd4998,17'd4999,17'd4999,17'd5000,17'd5001,17'd4529,17'd4688,17'd4845,17'd5002,17'd5003,17'd5003,17'd5004,17'd5005,17'd4848,17'd5006,17'd5007,17'd5007,17'd4848,17'd5008,17'd5009,17'd5010,17'd5011,17'd5012,17'd5013,17'd5014,17'd5015,17'd5016,17'd5017,17'd5018,17'd5019,17'd5020,17'd4215,17'd5021,17'd4044,17'd4217,17'd4218,17'd5022,17'd5023,17'd5024,17'd4394,17'd5025,17'd3872,17'd4227,17'd4554,17'd5026,17'd5027,17'd5028,17'd4883,17'd4869,17'd5029,17'd5030,17'd5031,17'd2574,17'd2914,17'd4870,17'd5032,17'd4404,17'd5033,17'd4871,17'd5034,17'd4406,17'd4873,17'd5035,17'd5036,17'd3228,17'd3228,17'd3400,17'd3575,17'd4064,17'd5037,17'd5037,17'd5038,17'd5039,17'd4410,17'd4410,17'd4721,17'd3233,17'd3233,17'd3083,17'd3084,17'd3884,17'd3409,17'd4074,17'd5040,17'd5041,17'd5042,17'd5043,17'd5044,17'd4725,17'd5045,17'd4079,17'd3243,17'd5046,17'd4879,17'd4418,17'd4418,17'd5047,17'd5046,17'd5048,17'd4574,17'd5049,17'd4241,17'd2559,17'd5050,17'd5050,17'd1680,17'd1680,17'd1401,17'd1261,17'd3391,17'd4729,17'd4713,17'd4869,17'd4869,17'd4713,17'd4883,17'd4883,17'd4883,17'd3897,17'd3423,17'd2586,17'd625,17'd623,17'd795,17'd795,17'd1402,17'd3072,17'd3898,17'd3898,17'd625,17'd446,17'd625,17'd1262,17'd1962,17'd954,17'd259,17'd259,17'd425,17'd425,17'd645,17'd1963,17'd645,17'd643,17'd206,17'd206,17'd1124,17'd1828,17'd1685,17'd1098,17'd1245,17'd1382,17'd2932,17'd1527
},
'{
17'd2,17'd1,17'd4884,17'd5051,17'd650,17'd283,17'd283,17'd650,17'd12,17'd14,17'd4886,17'd4887,17'd4088,17'd4087,17'd4734,17'd5052,17'd5053,17'd4890,17'd4426,17'd3902,17'd4244,17'd4244,17'd4087,17'd4426,17'd4893,17'd4738,17'd2592,17'd1967,17'd1127,17'd466,17'd2,17'd0,17'd2,17'd1127,17'd4247,17'd4247,17'd14,17'd14,17'd1127,17'd4247,17'd15,17'd2,17'd13,17'd12,17'd1128,17'd11,17'd21,17'd25,17'd22,17'd23,17'd4,17'd8,17'd6,17'd6,17'd3753,17'd3753,17'd5,17'd5,17'd5,17'd5,17'd23,17'd23,17'd1691,17'd2937,17'd1413,17'd25,17'd21,17'd20,17'd980,17'd980,17'd27,17'd27,17'd653,17'd653,17'd652,17'd652,17'd980,17'd27,17'd27,17'd27,17'd652,17'd652,17'd652,17'd28,17'd28,17'd28,17'd652,17'd652,17'd28,17'd652,17'd4430,17'd4091,17'd3595,17'd3255,17'd4249,17'd3104,17'd2604,17'd2604,17'd2604,17'd2604,17'd4894,17'd5054,17'd5055,17'd4741,17'd4895,17'd5056,17'd4740,17'd4740,17'd4896,17'd4896,17'd4253,17'd4253,17'd4254,17'd5057,17'd5057,17'd5058,17'd5059,17'd5059,17'd5060,17'd5061,17'd5062,17'd5063,17'd5064,17'd5065,17'd4748,17'd4904,17'd5066,17'd5067,17'd4751,17'd5068,17'd5069,17'd5070,17'd5071,17'd4911,17'd5072,17'd5073,17'd5074,17'd5075,17'd5076,17'd5077,17'd5078,17'd5079,17'd5080,17'd4456,17'd4603,17'd4763,17'd5081,17'd4921,17'd5082,17'd5083,17'd5084,17'd5085,17'd5086,17'd5087,17'd5088,17'd5088,17'd5089,17'd4925,17'd4925,17'd5090,17'd4767,17'd4767,17'd4926,17'd4766,17'd4291,17'd4292,17'd4123,17'd3955,17'd3632,17'd3956,17'd3634,17'd3789,17'd3635,17'd3141,17'd2988,17'd2981,17'd2825,17'd2656,17'd5091,17'd5092,17'd4617,17'd2659,17'd5093,17'd5094,17'd4302,17'd2306,17'd5095,17'd5096,17'd5097,17'd5098,17'd5099,17'd5100,17'd5101,17'd4479,17'd3319,17'd4480,17'd4481,17'd5102,17'd4483,17'd5103,17'd5103,17'd5104,17'd5104,17'd5105,17'd5106,17'd5107,17'd5108,17'd5109,17'd5110,17'd5111,17'd5112,17'd5113,17'd5114,17'd5115,17'd5116,17'd5117,17'd5118,17'd5119,17'd5120,17'd5121,17'd5122,17'd5123,17'd5124,17'd5125,17'd5126,17'd5127,17'd5128,17'd4969,17'd4652,17'd3511,17'd1195,17'd1480,17'd4163,17'd356,17'd1481,17'd1481,17'd1481,17'd541,17'd541,17'd1196,17'd719,17'd1197,17'd1197,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd135,17'd132,17'd132,17'd132,17'd135,17'd2698,17'd5129,17'd4814,17'd5130,17'd5131,17'd5132,17'd5133,17'd5134,17'd5135,17'd5136,17'd5137,17'd5138,17'd5139,17'd5140,17'd4183,17'd4987,17'd5141,17'd5141,17'd5142,17'd5143,17'd4519,17'd4676,17'd5144,17'd5145,17'd5146,17'd5147,17'd5148,17'd5149,17'd5150,17'd5151,17'd5152,17'd5153,17'd5154,17'd5155,17'd5155,17'd4526,17'd5156,17'd4529,17'd5157,17'd5002,17'd5002,17'd5158,17'd5159,17'd5160,17'd5160,17'd5161,17'd5162,17'd5162,17'd5162,17'd5163,17'd5009,17'd5164,17'd5165,17'd5166,17'd5167,17'd5168,17'd5169,17'd5170,17'd5171,17'd5172,17'd5017,17'd5018,17'd5173,17'd5174,17'd5175,17'd4214,17'd5176,17'd5021,17'd5177,17'd5178,17'd5179,17'd5024,17'd4054,17'd5025,17'd3710,17'd4395,17'd4554,17'd5180,17'd5181,17'd5182,17'd3896,17'd4869,17'd5183,17'd3074,17'd4561,17'd2751,17'd2913,17'd3396,17'd3573,17'd4232,17'd4405,17'd4562,17'd5034,17'd5184,17'd4873,17'd5036,17'd5185,17'd3227,17'd3228,17'd3396,17'd3575,17'd4064,17'd5037,17'd3082,17'd5038,17'd4565,17'd2755,17'd2757,17'd4721,17'd4568,17'd3233,17'd3083,17'd2757,17'd3579,17'd3579,17'd3727,17'd5041,17'd5186,17'd5042,17'd4723,17'd5187,17'd4877,17'd5188,17'd3243,17'd4079,17'd4879,17'd4418,17'd4418,17'd5189,17'd5046,17'd5190,17'd4726,17'd4574,17'd5191,17'd5192,17'd2392,17'd5050,17'd1261,17'd1680,17'd1261,17'd1261,17'd229,17'd5193,17'd4729,17'd4869,17'd5194,17'd4713,17'd4730,17'd4730,17'd4883,17'd3896,17'd3423,17'd3423,17'd2777,17'd2249,17'd795,17'd795,17'd1402,17'd3072,17'd3898,17'd5195,17'd624,17'd228,17'd228,17'd624,17'd1262,17'd953,17'd954,17'd259,17'd1112,17'd606,17'd803,17'd645,17'd803,17'd643,17'd206,17'd206,17'd1829,17'd1687,17'd1685,17'd1098,17'd603,17'd422,17'd2932,17'd1527
},
'{
17'd2,17'd1,17'd283,17'd283,17'd3,17'd283,17'd283,17'd1,17'd4885,17'd5196,17'd4577,17'd4088,17'd4087,17'd5197,17'd5198,17'd5198,17'd5199,17'd5200,17'd5201,17'd5202,17'd5202,17'd5201,17'd5203,17'd5204,17'd3751,17'd2784,17'd2781,17'd14,17'd2,17'd2,17'd14,17'd15,17'd4247,17'd1127,17'd1127,17'd1127,17'd1127,17'd1127,17'd2,17'd2,17'd2,17'd13,17'd18,17'd1128,17'd20,17'd21,17'd21,17'd25,17'd4,17'd4,17'd6,17'd6,17'd5205,17'd3753,17'd3753,17'd3594,17'd5,17'd6,17'd4,17'd23,17'd4,17'd8,17'd5206,17'd4,17'd467,17'd27,17'd980,17'd27,17'd286,17'd286,17'd27,17'd1278,17'd980,17'd980,17'd1278,17'd980,17'd285,17'd285,17'd20,17'd2598,17'd1128,17'd1128,17'd1128,17'd1128,17'd27,17'd27,17'd27,17'd28,17'd4430,17'd4431,17'd5207,17'd5208,17'd5209,17'd4249,17'd4579,17'd4250,17'd3105,17'd3105,17'd4739,17'd5210,17'd5210,17'd5211,17'd5211,17'd5212,17'd5213,17'd5056,17'd5214,17'd5215,17'd5216,17'd5217,17'd5058,17'd5218,17'd5219,17'd5219,17'd5220,17'd5221,17'd5222,17'd5223,17'd5224,17'd5225,17'd5226,17'd5227,17'd5228,17'd5229,17'd5230,17'd4905,17'd4590,17'd5231,17'd5232,17'd5233,17'd5234,17'd5235,17'd5236,17'd5237,17'd5238,17'd5239,17'd5240,17'd5241,17'd5242,17'd5243,17'd5244,17'd5245,17'd5246,17'd5247,17'd5248,17'd5249,17'd4125,17'd4125,17'd4126,17'd5250,17'd5250,17'd5251,17'd5088,17'd5252,17'd5253,17'd5254,17'd4927,17'd5255,17'd5255,17'd5090,17'd5090,17'd5256,17'd4928,17'd4766,17'd4291,17'd4292,17'd4123,17'd4123,17'd4128,17'd3475,17'd5257,17'd4771,17'd3140,17'd3136,17'd3467,17'd5258,17'd5259,17'd5260,17'd5092,17'd5261,17'd4617,17'd4775,17'd5262,17'd5263,17'd5264,17'd5265,17'd5266,17'd5267,17'd5268,17'd5269,17'd5270,17'd5271,17'd4784,17'd5272,17'd5273,17'd5274,17'd5275,17'd5276,17'd5277,17'd5278,17'd5279,17'd5280,17'd5281,17'd5282,17'd5283,17'd5284,17'd5285,17'd5286,17'd5287,17'd5288,17'd5289,17'd5290,17'd5291,17'd5292,17'd5293,17'd5294,17'd5295,17'd5296,17'd5297,17'd5298,17'd5299,17'd5300,17'd5301,17'd5302,17'd5303,17'd5304,17'd5126,17'd5305,17'd5306,17'd5307,17'd5308,17'd3335,17'd1044,17'd718,17'd542,17'd718,17'd1044,17'd5309,17'd5310,17'd5310,17'd1196,17'd541,17'd541,17'd1481,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd134,17'd132,17'd357,17'd3169,17'd5311,17'd5312,17'd4338,17'd5313,17'd5314,17'd5315,17'd5316,17'd5317,17'd5318,17'd5319,17'd5320,17'd5321,17'd4828,17'd4830,17'd4831,17'd4989,17'd4521,17'd4522,17'd4676,17'd5322,17'd5323,17'd5324,17'd5325,17'd4994,17'd5326,17'd5326,17'd4994,17'd5151,17'd5327,17'd5152,17'd5327,17'd5328,17'd4847,17'd4846,17'd4687,17'd4687,17'd5002,17'd5329,17'd5330,17'd5331,17'd5332,17'd5332,17'd5332,17'd5333,17'd5334,17'd5330,17'd5329,17'd5329,17'd5329,17'd5160,17'd5160,17'd5335,17'd5335,17'd5336,17'd5168,17'd5337,17'd5338,17'd5339,17'd5340,17'd5341,17'd5342,17'd5343,17'd5344,17'd5345,17'd5346,17'd5347,17'd4548,17'd5348,17'd5349,17'd5350,17'd5351,17'd5352,17'd5353,17'd3710,17'd4710,17'd5354,17'd5355,17'd5356,17'd5357,17'd3247,17'd2905,17'd5358,17'd5359,17'd5360,17'd5361,17'd5362,17'd5363,17'd5364,17'd3397,17'd4873,17'd5184,17'd5365,17'd5365,17'd5366,17'd3877,17'd5185,17'd3227,17'd3078,17'd3400,17'd3399,17'd5367,17'd4408,17'd4067,17'd2405,17'd2405,17'd5038,17'd4069,17'd3405,17'd3406,17'd3406,17'd3406,17'd3083,17'd3579,17'd3886,17'd5368,17'd5368,17'd5369,17'd5370,17'd5043,17'd5187,17'd4725,17'd2926,17'd2768,17'd4417,17'd5190,17'd5189,17'd5047,17'd4571,17'd4417,17'd3417,17'd4877,17'd4237,17'd3585,17'd2585,17'd2559,17'd2559,17'd445,17'd1261,17'd1261,17'd4881,17'd4880,17'd5371,17'd5372,17'd4728,17'd4882,17'd4882,17'd4882,17'd4730,17'd4883,17'd4867,17'd5373,17'd3247,17'd4424,17'd625,17'd1544,17'd1114,17'd623,17'd625,17'd624,17'd3247,17'd2586,17'd1119,17'd1119,17'd1119,17'd624,17'd2249,17'd953,17'd259,17'd260,17'd206,17'd803,17'd973,17'd1687,17'd269,17'd272,17'd270,17'd272,17'd803,17'd1686,17'd1821,17'd1246,17'd1527,17'd420
},
'{
17'd0,17'd1,17'd283,17'd283,17'd3,17'd1,17'd0,17'd14,17'd4886,17'd4577,17'd3904,17'd3903,17'd4735,17'd5374,17'd5375,17'd5375,17'd5199,17'd5200,17'd5376,17'd5377,17'd5376,17'd4735,17'd5203,17'd3592,17'd2593,17'd2422,17'd1689,17'd14,17'd0,17'd0,17'd14,17'd14,17'd1688,17'd1689,17'd1127,17'd1127,17'd1127,17'd1127,17'd2,17'd2,17'd2,17'd12,17'd1128,17'd11,17'd20,17'd21,17'd25,17'd25,17'd4,17'd4,17'd6,17'd6,17'd3753,17'd3753,17'd3594,17'd3594,17'd5,17'd4,17'd4,17'd4,17'd5206,17'd5378,17'd8,17'd23,17'd286,17'd1833,17'd1833,17'd286,17'd27,17'd980,17'd980,17'd27,17'd1278,17'd980,17'd27,17'd286,17'd285,17'd26,17'd20,17'd2598,17'd1128,17'd1128,17'd1128,17'd11,17'd27,17'd27,17'd27,17'd28,17'd4431,17'd4431,17'd3910,17'd5208,17'd4249,17'd4249,17'd4251,17'd4250,17'd3104,17'd3104,17'd4250,17'd5210,17'd5379,17'd5379,17'd5211,17'd5211,17'd5056,17'd5056,17'd5215,17'd5215,17'd5380,17'd5220,17'd5220,17'd5381,17'd4742,17'd5382,17'd5383,17'd5384,17'd5385,17'd5386,17'd5387,17'd5388,17'd5389,17'd5390,17'd5391,17'd4749,17'd5392,17'd5393,17'd5394,17'd5395,17'd5396,17'd5397,17'd5235,17'd5398,17'd5399,17'd5238,17'd5239,17'd5400,17'd5401,17'd5402,17'd5403,17'd5404,17'd5245,17'd5405,17'd5406,17'd5407,17'd5408,17'd4125,17'd4126,17'd4126,17'd5250,17'd5250,17'd5251,17'd5088,17'd5252,17'd5252,17'd5253,17'd5253,17'd5255,17'd5255,17'd5409,17'd5410,17'd5256,17'd4928,17'd4766,17'd4127,17'd4292,17'd3785,17'd4123,17'd4122,17'd3948,17'd5411,17'd3299,17'd3139,17'd3136,17'd2984,17'd3135,17'd5412,17'd5413,17'd5414,17'd5415,17'd5261,17'd5261,17'd5261,17'd5265,17'd5416,17'd5417,17'd5418,17'd5419,17'd5420,17'd5421,17'd5422,17'd5423,17'd5424,17'd5425,17'd5426,17'd5427,17'd5428,17'd5429,17'd5430,17'd5282,17'd5431,17'd5432,17'd5433,17'd5434,17'd5435,17'd5436,17'd5437,17'd5438,17'd5439,17'd5440,17'd5441,17'd5442,17'd5443,17'd5444,17'd5445,17'd5446,17'd5447,17'd5448,17'd5449,17'd5450,17'd5451,17'd5452,17'd5453,17'd5454,17'd5455,17'd5456,17'd5457,17'd5458,17'd5304,17'd5305,17'd5306,17'd5459,17'd886,17'd5460,17'd5461,17'd5462,17'd5463,17'd5464,17'd5465,17'd3511,17'd540,17'd541,17'd541,17'd541,17'd1480,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd1197,17'd132,17'd131,17'd3168,17'd5466,17'd5467,17'd5468,17'd5469,17'd5470,17'd4503,17'd5471,17'd5472,17'd4982,17'd5473,17'd5474,17'd4353,17'd5475,17'd5476,17'd4356,17'd4018,17'd5477,17'd4990,17'd4523,17'd4837,17'd5323,17'd4993,17'd5150,17'd5478,17'd5326,17'd5326,17'd5479,17'd5326,17'd5150,17'd5480,17'd5328,17'd4841,17'd4686,17'd4686,17'd5005,17'd5002,17'd5002,17'd5329,17'd5330,17'd5481,17'd5158,17'd5158,17'd5331,17'd5331,17'd5482,17'd5482,17'd5334,17'd5334,17'd5330,17'd5330,17'd5160,17'd5160,17'd5335,17'd5335,17'd5336,17'd5336,17'd5337,17'd5337,17'd5169,17'd5339,17'd5483,17'd5484,17'd5485,17'd5486,17'd5487,17'd5488,17'd5489,17'd4214,17'd5490,17'd4047,17'd5491,17'd5492,17'd5493,17'd5494,17'd4708,17'd3872,17'd4710,17'd5495,17'd5496,17'd5497,17'd4424,17'd3742,17'd2576,17'd5358,17'd5498,17'd3075,17'd5499,17'd5500,17'd5363,17'd5364,17'd4403,17'd4873,17'd5501,17'd5501,17'd5502,17'd5366,17'd5185,17'd5503,17'd3227,17'd3227,17'd3399,17'd3399,17'd3575,17'd4408,17'd3082,17'd2405,17'd4069,17'd4069,17'd3405,17'd3405,17'd3405,17'd3405,17'd4721,17'd2756,17'd3886,17'd3887,17'd5504,17'd5505,17'd5370,17'd5369,17'd5043,17'd5187,17'd4877,17'd2926,17'd3243,17'd4417,17'd4879,17'd5189,17'd4571,17'd4571,17'd4079,17'd4726,17'd4877,17'd5506,17'd4241,17'd2765,17'd2417,17'd445,17'd1261,17'd1261,17'd5507,17'd4881,17'd4881,17'd4880,17'd4423,17'd4423,17'd4882,17'd4882,17'd4730,17'd4883,17'd4867,17'd4867,17'd3897,17'd2096,17'd2586,17'd446,17'd231,17'd443,17'd446,17'd624,17'd2586,17'd3246,17'd3246,17'd3246,17'd1119,17'd1119,17'd625,17'd2249,17'd954,17'd259,17'd206,17'd644,17'd973,17'd1687,17'd269,17'd270,17'd270,17'd272,17'd803,17'd191,17'd1099,17'd1246,17'd420,17'd419
},
'{
17'd0,17'd1,17'd1,17'd1,17'd1,17'd0,17'd1127,17'd1831,17'd5508,17'd4246,17'd4428,17'd4426,17'd4888,17'd5509,17'd5375,17'd5510,17'd5199,17'd5199,17'd5376,17'd5376,17'd4735,17'd4578,17'd5511,17'd3427,17'd2592,17'd3250,17'd1689,17'd14,17'd0,17'd0,17'd14,17'd4247,17'd1127,17'd1127,17'd1127,17'd1127,17'd1127,17'd1127,17'd14,17'd2,17'd0,17'd12,17'd1128,17'd11,17'd21,17'd21,17'd23,17'd23,17'd6,17'd6,17'd3753,17'd3753,17'd3753,17'd3753,17'd3594,17'd3594,17'd6,17'd4,17'd8,17'd5512,17'd5513,17'd5514,17'd1413,17'd25,17'd4429,17'd5515,17'd4429,17'd1833,17'd27,17'd980,17'd3906,17'd26,17'd5516,17'd26,17'd467,17'd467,17'd22,17'd5517,17'd5517,17'd5518,17'd20,17'd20,17'd11,17'd11,17'd27,17'd286,17'd28,17'd28,17'd4431,17'd4091,17'd5208,17'd5209,17'd4249,17'd5519,17'd5520,17'd4579,17'd5379,17'd5379,17'd5379,17'd5379,17'd5210,17'd5210,17'd5055,17'd5055,17'd4741,17'd4740,17'd4740,17'd4740,17'd5214,17'd5221,17'd5221,17'd5221,17'd5521,17'd5384,17'd5522,17'd5385,17'd5523,17'd5524,17'd5525,17'd5389,17'd5526,17'd4265,17'd5527,17'd5528,17'd5529,17'd5530,17'd5395,17'd5531,17'd5397,17'd5532,17'd5533,17'd5534,17'd4913,17'd5535,17'd5536,17'd5537,17'd5538,17'd5539,17'd5540,17'd5541,17'd5542,17'd5543,17'd5544,17'd5545,17'd5408,17'd4768,17'd4610,17'd4610,17'd5088,17'd4925,17'd4925,17'd4925,17'd5253,17'd5253,17'd5255,17'd5255,17'd5255,17'd5255,17'd5410,17'd5090,17'd4766,17'd4610,17'd4768,17'd4291,17'd3954,17'd3786,17'd3629,17'd3628,17'd3948,17'd5411,17'd3298,17'd3297,17'd3296,17'd2984,17'd2983,17'd2824,17'd2657,17'd5546,17'd5547,17'd5415,17'd5415,17'd5547,17'd5547,17'd5547,17'd5548,17'd5549,17'd5550,17'd5551,17'd5552,17'd5553,17'd5554,17'd5555,17'd5556,17'd4476,17'd5557,17'd5558,17'd5559,17'd5560,17'd5561,17'd5562,17'd5563,17'd5563,17'd5564,17'd5565,17'd5566,17'd5567,17'd5438,17'd5568,17'd5569,17'd5570,17'd5571,17'd5572,17'd5573,17'd5574,17'd5575,17'd5576,17'd5577,17'd5578,17'd5579,17'd5580,17'd5581,17'd5582,17'd5583,17'd5584,17'd5585,17'd5586,17'd5587,17'd5588,17'd5589,17'd5125,17'd5126,17'd5590,17'd4969,17'd5591,17'd5591,17'd5592,17'd4971,17'd2511,17'd2037,17'd539,17'd540,17'd541,17'd1481,17'd1481,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd542,17'd542,17'd132,17'd132,17'd131,17'd3168,17'd5593,17'd5468,17'd5594,17'd5595,17'd5596,17'd5597,17'd5598,17'd5599,17'd5600,17'd5601,17'd5602,17'd5603,17'd4987,17'd4830,17'd5604,17'd5477,17'd5605,17'd5605,17'd4681,17'd5606,17'd5607,17'd5608,17'd4994,17'd5478,17'd5609,17'd5610,17'd5610,17'd5610,17'd5609,17'd5478,17'd5609,17'd5609,17'd4844,17'd5611,17'd5611,17'd5481,17'd5481,17'd5481,17'd5482,17'd5482,17'd5612,17'd5613,17'd5158,17'd5158,17'd5482,17'd5482,17'd5334,17'd5334,17'd5336,17'd5336,17'd5335,17'd5335,17'd5335,17'd5336,17'd5614,17'd5614,17'd5615,17'd5337,17'd5616,17'd5617,17'd5618,17'd5619,17'd5620,17'd5621,17'd5018,17'd5622,17'd5623,17'd4384,17'd4216,17'd5177,17'd5348,17'd5624,17'd5625,17'd5493,17'd5626,17'd4708,17'd3710,17'd5627,17'd5628,17'd2558,17'd5629,17'd2586,17'd3391,17'd5630,17'd5631,17'd2741,17'd3075,17'd5632,17'd5633,17'd5634,17'd3573,17'd4403,17'd5635,17'd5501,17'd5502,17'd5502,17'd5636,17'd5637,17'd5638,17'd3227,17'd3399,17'd5032,17'd5639,17'd4064,17'd3082,17'd3082,17'd4069,17'd3720,17'd3720,17'd3720,17'd4410,17'd4410,17'd4721,17'd3233,17'd2757,17'd3409,17'd3727,17'd5368,17'd5369,17'd5370,17'd5640,17'd5641,17'd5044,17'd5642,17'd4079,17'd3737,17'd4417,17'd5046,17'd4879,17'd4571,17'd3243,17'd3417,17'd4877,17'd4725,17'd5049,17'd3422,17'd2559,17'd2392,17'd445,17'd1261,17'd3743,17'd3743,17'd5507,17'd5507,17'd5372,17'd5372,17'd4713,17'd4882,17'd4730,17'd4730,17'd4883,17'd4883,17'd4575,17'd2096,17'd2096,17'd2777,17'd446,17'd231,17'd227,17'd625,17'd2586,17'd2586,17'd3423,17'd3423,17'd2586,17'd1119,17'd624,17'd1680,17'd1243,17'd259,17'd206,17'd644,17'd1963,17'd803,17'd270,17'd270,17'd270,17'd272,17'd803,17'd191,17'd1099,17'd1246,17'd420,17'd419
},
'{
17'd0,17'd0,17'd0,17'd1,17'd1830,17'd15,17'd1689,17'd2935,17'd4245,17'd4428,17'd4427,17'd4735,17'd5052,17'd5509,17'd5643,17'd5644,17'd5644,17'd5199,17'd5376,17'd5645,17'd4734,17'd5646,17'd5204,17'd2934,17'd2592,17'd1689,17'd14,17'd15,17'd0,17'd14,17'd1127,17'd4247,17'd1127,17'd1127,17'd14,17'd1127,17'd1127,17'd1127,17'd1127,17'd14,17'd0,17'd0,17'd19,17'd11,17'd21,17'd25,17'd23,17'd23,17'd6,17'd6,17'd3753,17'd3753,17'd3753,17'd3753,17'd3594,17'd5,17'd4,17'd4,17'd5647,17'd5648,17'd5649,17'd5650,17'd5651,17'd5652,17'd5653,17'd5654,17'd5515,17'd286,17'd27,17'd27,17'd3906,17'd3906,17'd26,17'd285,17'd2937,17'd467,17'd22,17'd5517,17'd5518,17'd5518,17'd21,17'd20,17'd11,17'd11,17'd286,17'd28,17'd28,17'd29,17'd4091,17'd4091,17'd5208,17'd5209,17'd4249,17'd4249,17'd4579,17'd5655,17'd5656,17'd5656,17'd5656,17'd5657,17'd5658,17'd5658,17'd5055,17'd5055,17'd4741,17'd4741,17'd4741,17'd4741,17'd5521,17'd5659,17'd5659,17'd5660,17'd5661,17'd5662,17'd5663,17'd5386,17'd5664,17'd5525,17'd5665,17'd5666,17'd5667,17'd5668,17'd5669,17'd5670,17'd5671,17'd5672,17'd5673,17'd5674,17'd5675,17'd5676,17'd5677,17'd5678,17'd5679,17'd5239,17'd5537,17'd5680,17'd5681,17'd5682,17'd5683,17'd5684,17'd5543,17'd5685,17'd5686,17'd5408,17'd5687,17'd5688,17'd5688,17'd4928,17'd4925,17'd4925,17'd4925,17'd4925,17'd5253,17'd5255,17'd5255,17'd5689,17'd5255,17'd5255,17'd5410,17'd4767,17'd4127,17'd4291,17'd4291,17'd3951,17'd3786,17'd3629,17'd3948,17'd3473,17'd3473,17'd3298,17'd3297,17'd3469,17'd3294,17'd5690,17'd2824,17'd5691,17'd5692,17'd5693,17'd5694,17'd5695,17'd5694,17'd5694,17'd5696,17'd5696,17'd5696,17'd5697,17'd5698,17'd5699,17'd5700,17'd5420,17'd5552,17'd5553,17'd5701,17'd5702,17'd5703,17'd5704,17'd5705,17'd5706,17'd5707,17'd5708,17'd5709,17'd5710,17'd5711,17'd5712,17'd5713,17'd5714,17'd5715,17'd5716,17'd5717,17'd5718,17'd5719,17'd5720,17'd5721,17'd5722,17'd5723,17'd5724,17'd5725,17'd5726,17'd5727,17'd5728,17'd5729,17'd5730,17'd5731,17'd5732,17'd5733,17'd5734,17'd5735,17'd5736,17'd5737,17'd5587,17'd5738,17'd5739,17'd5740,17'd5741,17'd5742,17'd5743,17'd2858,17'd2037,17'd1477,17'd2340,17'd541,17'd541,17'd1481,17'd1481,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd542,17'd542,17'd132,17'd132,17'd3168,17'd5744,17'd5745,17'd4338,17'd5746,17'd5747,17'd5748,17'd5598,17'd5749,17'd5750,17'd5751,17'd5752,17'd5753,17'd4984,17'd4829,17'd4831,17'd5754,17'd4676,17'd5755,17'd5756,17'd5606,17'd5757,17'd5608,17'd4994,17'd5478,17'd5478,17'd5610,17'd5610,17'd5758,17'd5758,17'd5758,17'd5758,17'd5758,17'd5759,17'd5482,17'd5482,17'd5482,17'd5760,17'd5760,17'd5760,17'd5760,17'd5760,17'd5761,17'd5761,17'd5331,17'd5158,17'd5481,17'd5481,17'd5334,17'd5334,17'd5336,17'd5336,17'd5336,17'd5762,17'd5762,17'd5762,17'd5614,17'd5615,17'd5615,17'd5615,17'd5763,17'd5764,17'd5765,17'd5618,17'd5172,17'd5620,17'd5766,17'd5767,17'd5488,17'd5768,17'd5769,17'd4043,17'd4217,17'd3858,17'd5770,17'd5771,17'd5772,17'd4224,17'd5773,17'd5774,17'd3874,17'd5775,17'd2391,17'd4400,17'd3099,17'd3744,17'd5776,17'd5777,17'd5360,17'd5778,17'd2912,17'd3226,17'd4870,17'd3573,17'd4233,17'd5366,17'd5502,17'd5779,17'd5780,17'd5781,17'd5782,17'd5638,17'd3227,17'd3574,17'd4233,17'd5639,17'd4720,17'd4564,17'd3082,17'd4069,17'd4069,17'd3720,17'd3405,17'd3405,17'd2756,17'd3233,17'd4721,17'd2756,17'd5783,17'd3727,17'd3727,17'd5369,17'd5186,17'd5042,17'd4875,17'd5784,17'd5785,17'd3243,17'd3243,17'd5046,17'd4879,17'd4879,17'd3243,17'd3243,17'd4573,17'd4725,17'd5786,17'd5787,17'd5788,17'd4422,17'd1810,17'd2392,17'd5050,17'd3743,17'd4881,17'd4881,17'd5371,17'd5371,17'd4713,17'd4882,17'd5789,17'd5789,17'd4730,17'd4883,17'd4730,17'd4575,17'd3897,17'd2096,17'd1119,17'd227,17'd231,17'd446,17'd1119,17'd2586,17'd3897,17'd3897,17'd2586,17'd1119,17'd1119,17'd2777,17'd1380,17'd970,17'd260,17'd644,17'd645,17'd645,17'd272,17'd269,17'd270,17'd272,17'd803,17'd1098,17'd2116,17'd1246,17'd420,17'd416
},
'{
17'd12,17'd0,17'd0,17'd15,17'd3249,17'd2781,17'd4887,17'd4245,17'd4428,17'd4427,17'd5201,17'd5197,17'd5052,17'd5509,17'd5790,17'd5791,17'd5792,17'd5792,17'd5645,17'd5197,17'd4734,17'd4891,17'd3901,17'd2935,17'd3250,17'd1967,17'd15,17'd0,17'd14,17'd1127,17'd1127,17'd1689,17'd1127,17'd1127,17'd14,17'd1127,17'd1689,17'd1689,17'd1127,17'd14,17'd0,17'd12,17'd11,17'd10,17'd25,17'd23,17'd24,17'd5,17'd6,17'd6,17'd3753,17'd3753,17'd5793,17'd5793,17'd3594,17'd3594,17'd5,17'd5647,17'd5794,17'd5795,17'd5796,17'd5797,17'd5798,17'd5799,17'd5800,17'd5799,17'd5801,17'd3748,17'd979,17'd11,17'd26,17'd26,17'd1691,17'd1691,17'd23,17'd22,17'd284,17'd5802,17'd284,17'd22,17'd21,17'd21,17'd11,17'd10,17'd287,17'd28,17'd652,17'd29,17'd3908,17'd3595,17'd5209,17'd5209,17'd5209,17'd5208,17'd5208,17'd3910,17'd5803,17'd5803,17'd5804,17'd5656,17'd5657,17'd5658,17'd5055,17'd5805,17'd5805,17'd5806,17'd5807,17'd5808,17'd5809,17'd5810,17'd5811,17'd5812,17'd5813,17'd5814,17'd5386,17'd5524,17'd5525,17'd5665,17'd5815,17'd3924,17'd5816,17'd5817,17'd5818,17'd5819,17'd5820,17'd5821,17'd5822,17'd5823,17'd5824,17'd5825,17'd5237,17'd5238,17'd5826,17'd5827,17'd5828,17'd5829,17'd5830,17'd5831,17'd5832,17'd5833,17'd5834,17'd5835,17'd5687,17'd5250,17'd4928,17'd5090,17'd5836,17'd5836,17'd5689,17'd5837,17'd5409,17'd5409,17'd5409,17'd5409,17'd5409,17'd5837,17'd5090,17'd5090,17'd4767,17'd4767,17'd4127,17'd3951,17'd3951,17'd3784,17'd3629,17'd3948,17'd3782,17'd5838,17'd5839,17'd5840,17'd5841,17'd5842,17'd5690,17'd5843,17'd5844,17'd5845,17'd5846,17'd5692,17'd5847,17'd5847,17'd5848,17'd5845,17'd5849,17'd5844,17'd5850,17'd5851,17'd5852,17'd5693,17'd5853,17'd5550,17'd5854,17'd5855,17'd5856,17'd5857,17'd5858,17'd5859,17'd5860,17'd5861,17'd5861,17'd5862,17'd5863,17'd5864,17'd5865,17'd5866,17'd5867,17'd5868,17'd5869,17'd5870,17'd5871,17'd5872,17'd5873,17'd5874,17'd5875,17'd5876,17'd5877,17'd5878,17'd5879,17'd5880,17'd5881,17'd5882,17'd5883,17'd5884,17'd5885,17'd5886,17'd5887,17'd5888,17'd5889,17'd5890,17'd5891,17'd5892,17'd5893,17'd5457,17'd5894,17'd5895,17'd5896,17'd5897,17'd2858,17'd2859,17'd1476,17'd1479,17'd3995,17'd541,17'd1197,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd719,17'd3025,17'd5898,17'd4336,17'd5899,17'd5900,17'd2864,17'd5901,17'd5902,17'd5903,17'd5904,17'd5905,17'd5906,17'd5139,17'd5907,17'd5908,17'd5909,17'd5910,17'd5911,17'd5605,17'd4837,17'd4837,17'd4837,17'd5912,17'd4992,17'd5608,17'd5326,17'd5610,17'd5610,17'd5913,17'd5914,17'd5915,17'd5915,17'd5915,17'd5916,17'd5916,17'd5916,17'd5917,17'd5917,17'd5917,17'd5917,17'd5917,17'd5917,17'd5917,17'd5917,17'd5918,17'd5918,17'd5916,17'd5915,17'd5482,17'd5482,17'd5331,17'd5331,17'd5335,17'd5336,17'd5614,17'd5615,17'd5615,17'd5919,17'd5615,17'd5615,17'd5615,17'd5615,17'd5763,17'd5764,17'd5920,17'd5765,17'd5921,17'd5922,17'd5923,17'd5342,17'd5924,17'd5925,17'd5926,17'd5927,17'd5928,17'd5929,17'd5930,17'd5931,17'd5023,17'd5772,17'd5932,17'd5933,17'd5934,17'd5935,17'd5936,17'd5937,17'd5938,17'd5939,17'd3744,17'd5940,17'd5941,17'd5942,17'd5943,17'd5944,17'd3876,17'd3396,17'd3398,17'd3574,17'd5366,17'd5779,17'd5780,17'd5781,17'd5780,17'd5945,17'd3227,17'd3574,17'd3574,17'd4233,17'd5946,17'd5947,17'd4564,17'd3082,17'd4069,17'd4069,17'd3720,17'd5948,17'd2756,17'd2756,17'd5949,17'd3233,17'd2757,17'd4075,17'd4414,17'd4414,17'd5504,17'd5369,17'd5950,17'd4723,17'd5951,17'd3093,17'd3243,17'd3243,17'd5046,17'd5190,17'd5046,17'd4417,17'd4079,17'd5952,17'd5953,17'd5954,17'd5955,17'd5956,17'd5192,17'd2559,17'd445,17'd445,17'd5050,17'd5957,17'd5371,17'd5371,17'd4729,17'd4713,17'd4882,17'd5958,17'd4730,17'd4730,17'd5789,17'd4883,17'd3897,17'd2240,17'd2096,17'd1119,17'd227,17'd231,17'd228,17'd2586,17'd3897,17'd3897,17'd3423,17'd2586,17'd2586,17'd2777,17'd2775,17'd1243,17'd259,17'd970,17'd803,17'd645,17'd273,17'd269,17'd270,17'd272,17'd1828,17'd1098,17'd2116,17'd1246,17'd419,17'd197
},
'{
17'd3,17'd0,17'd15,17'd3249,17'd2781,17'd2782,17'd4428,17'd4244,17'd4427,17'd5202,17'd5645,17'd5374,17'd5374,17'd5959,17'd5790,17'd5644,17'd5792,17'd5960,17'd5197,17'd4734,17'd5646,17'd4244,17'd2593,17'd2592,17'd1688,17'd14,17'd0,17'd2,17'd1127,17'd4247,17'd1689,17'd1967,17'd1127,17'd1127,17'd14,17'd1127,17'd1689,17'd1689,17'd1127,17'd14,17'd0,17'd0,17'd19,17'd10,17'd25,17'd4,17'd5,17'd5,17'd6,17'd6,17'd3753,17'd3753,17'd5793,17'd3753,17'd3753,17'd6,17'd5206,17'd5514,17'd5795,17'd5961,17'd5962,17'd5963,17'd5964,17'd5965,17'd5966,17'd5967,17'd5968,17'd5801,17'd5969,17'd19,17'd286,17'd2937,17'd5970,17'd1691,17'd22,17'd5518,17'd284,17'd284,17'd284,17'd284,17'd22,17'd21,17'd10,17'd10,17'd28,17'd28,17'd29,17'd289,17'd3595,17'd3595,17'd5208,17'd5208,17'd5208,17'd3910,17'd3910,17'd5971,17'd5972,17'd5973,17'd5803,17'd5804,17'd5657,17'd5657,17'd5806,17'd5806,17'd5806,17'd5974,17'd5975,17'd5976,17'd5977,17'd5977,17'd5978,17'd5979,17'd5814,17'd5814,17'd5523,17'd5525,17'd5665,17'd5815,17'd5980,17'd5981,17'd5982,17'd5983,17'd5984,17'd5671,17'd5985,17'd5986,17'd5987,17'd5988,17'd5989,17'd5678,17'd5238,17'd5239,17'd5827,17'd5990,17'd5991,17'd5992,17'd5993,17'd5994,17'd5995,17'd5996,17'd5997,17'd5688,17'd5998,17'd5251,17'd5089,17'd5836,17'd5836,17'd5689,17'd5837,17'd5837,17'd5837,17'd5409,17'd5409,17'd5409,17'd5409,17'd5409,17'd5090,17'd4767,17'd4611,17'd4464,17'd3951,17'd3950,17'd3784,17'd3628,17'd3948,17'd3473,17'd5838,17'd5839,17'd5999,17'd6000,17'd5842,17'd6001,17'd5843,17'd5843,17'd5849,17'd5849,17'd5849,17'd5845,17'd5848,17'd6002,17'd6003,17'd6004,17'd6005,17'd6000,17'd6006,17'd6007,17'd2824,17'd5844,17'd5852,17'd6008,17'd6009,17'd6010,17'd6011,17'd6012,17'd6013,17'd6014,17'd6015,17'd6016,17'd6017,17'd6018,17'd6019,17'd6020,17'd6021,17'd6022,17'd6023,17'd6024,17'd6025,17'd6026,17'd6027,17'd6028,17'd6029,17'd6030,17'd6031,17'd6032,17'd6033,17'd6034,17'd6035,17'd6036,17'd6037,17'd6038,17'd6039,17'd6040,17'd6041,17'd6042,17'd6043,17'd6044,17'd6045,17'd6046,17'd6047,17'd6048,17'd6049,17'd6050,17'd6051,17'd6052,17'd6053,17'd6054,17'd5459,17'd3511,17'd2340,17'd1478,17'd541,17'd541,17'd1197,17'd1197,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd1197,17'd134,17'd6055,17'd6056,17'd3813,17'd6057,17'd5596,17'd6058,17'd6059,17'd6060,17'd6061,17'd6062,17'd6063,17'd6064,17'd6065,17'd6066,17'd5911,17'd4522,17'd4838,17'd4837,17'd4681,17'd6067,17'd5323,17'd5607,17'd4994,17'd5326,17'd5610,17'd5913,17'd5914,17'd5914,17'd5915,17'd5916,17'd5916,17'd5917,17'd5917,17'd5917,17'd6068,17'd6068,17'd6068,17'd6068,17'd6068,17'd6068,17'd6068,17'd5917,17'd5918,17'd5918,17'd5916,17'd5916,17'd5760,17'd5760,17'd5332,17'd5332,17'd5335,17'd5336,17'd5614,17'd5615,17'd5919,17'd5919,17'd5919,17'd5919,17'd5615,17'd5615,17'd5763,17'd5763,17'd5764,17'd5920,17'd6069,17'd5921,17'd6070,17'd6071,17'd6072,17'd6073,17'd6074,17'd6075,17'd6076,17'd6077,17'd6078,17'd4704,17'd6079,17'd6080,17'd6081,17'd6082,17'd6083,17'd6084,17'd4228,17'd5496,17'd6085,17'd5939,17'd3246,17'd5371,17'd2575,17'd5941,17'd4561,17'd6086,17'd2913,17'd3876,17'd3400,17'd3398,17'd5503,17'd5036,17'd5637,17'd5780,17'd5780,17'd5637,17'd6087,17'd6087,17'd3574,17'd3574,17'd4062,17'd5946,17'd4409,17'd3082,17'd4069,17'd4069,17'd3720,17'd5948,17'd4721,17'd2757,17'd2759,17'd6088,17'd2756,17'd3084,17'd3084,17'd4075,17'd5504,17'd5368,17'd6089,17'd5950,17'd6090,17'd5953,17'd5188,17'd3740,17'd5046,17'd5190,17'd5190,17'd5046,17'd3243,17'd5048,17'd6091,17'd5951,17'd6092,17'd6093,17'd5956,17'd3742,17'd2392,17'd445,17'd5957,17'd5957,17'd5371,17'd5371,17'd3744,17'd4729,17'd4882,17'd5958,17'd5789,17'd4730,17'd6094,17'd6095,17'd3896,17'd4575,17'd4575,17'd3247,17'd228,17'd227,17'd1260,17'd1119,17'd3423,17'd3897,17'd3897,17'd3423,17'd3247,17'd3247,17'd2559,17'd1380,17'd1243,17'd970,17'd644,17'd645,17'd274,17'd269,17'd270,17'd270,17'd1828,17'd1098,17'd2116,17'd421,17'd198,17'd197
},
'{
17'd0,17'd0,17'd4885,17'd6096,17'd4887,17'd4428,17'd3902,17'd5202,17'd5377,17'd5960,17'd5198,17'd5198,17'd5198,17'd5643,17'd5645,17'd5960,17'd5792,17'd5960,17'd5197,17'd4888,17'd4426,17'd3904,17'd2592,17'd2781,17'd1689,17'd14,17'd2,17'd466,17'd1127,17'd4247,17'd1689,17'd1967,17'd1127,17'd1127,17'd1689,17'd1689,17'd1689,17'd1689,17'd1127,17'd14,17'd0,17'd12,17'd11,17'd21,17'd23,17'd4,17'd6,17'd3753,17'd6,17'd6,17'd3753,17'd3753,17'd3753,17'd3753,17'd3753,17'd6,17'd6097,17'd6098,17'd6099,17'd6100,17'd6101,17'd6102,17'd6103,17'd6104,17'd6105,17'd6106,17'd6100,17'd6107,17'd5801,17'd6108,17'd5651,17'd5512,17'd8,17'd23,17'd284,17'd5802,17'd284,17'd24,17'd24,17'd284,17'd22,17'd21,17'd27,17'd27,17'd28,17'd652,17'd4091,17'd3595,17'd3595,17'd3595,17'd5208,17'd3910,17'd5207,17'd5971,17'd5971,17'd5971,17'd5973,17'd5973,17'd5803,17'd5803,17'd5656,17'd5656,17'd5657,17'd5657,17'd6109,17'd6110,17'd5976,17'd6111,17'd6111,17'd6112,17'd6113,17'd5979,17'd5814,17'd5224,17'd6114,17'd6115,17'd6116,17'd5815,17'd4264,17'd6117,17'd6118,17'd6119,17'd5529,17'd6120,17'd6121,17'd6122,17'd6123,17'd6124,17'd6125,17'd6126,17'd6127,17'd5536,17'd6128,17'd6129,17'd6130,17'd6131,17'd5994,17'd6132,17'd6133,17'd6134,17'd6135,17'd6136,17'd6137,17'd6138,17'd6139,17'd6140,17'd6141,17'd6141,17'd6142,17'd6142,17'd6142,17'd6142,17'd6143,17'd6143,17'd5409,17'd5409,17'd4767,17'd4926,17'd4464,17'd4127,17'd3951,17'd3784,17'd3784,17'd3628,17'd3782,17'd5838,17'd5838,17'd5839,17'd5999,17'd6000,17'd5842,17'd6144,17'd5843,17'd5843,17'd6145,17'd6145,17'd5844,17'd6146,17'd6147,17'd6148,17'd6149,17'd6150,17'd6150,17'd6151,17'd6152,17'd3469,17'd3468,17'd6007,17'd6005,17'd6153,17'd6154,17'd6155,17'd6155,17'd6155,17'd6156,17'd6157,17'd6158,17'd6159,17'd6160,17'd6160,17'd6161,17'd6162,17'd6163,17'd6164,17'd6165,17'd6166,17'd6167,17'd6168,17'd6169,17'd6170,17'd6171,17'd6172,17'd6173,17'd6174,17'd6175,17'd6176,17'd6177,17'd6178,17'd6179,17'd6180,17'd6181,17'd6182,17'd6183,17'd6184,17'd6185,17'd6186,17'd6187,17'd6188,17'd6189,17'd6190,17'd6191,17'd6192,17'd6193,17'd6194,17'd6195,17'd6196,17'd6197,17'd5460,17'd3335,17'd3337,17'd6198,17'd6198,17'd1197,17'd1197,17'd1197,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd132,17'd133,17'd133,17'd132,17'd357,17'd3512,17'd6199,17'd6200,17'd6201,17'd6202,17'd5472,17'd6203,17'd6204,17'd6205,17'd6206,17'd6065,17'd6207,17'd6208,17'd6209,17'd6210,17'd5322,17'd5607,17'd5607,17'd4993,17'd4994,17'd4994,17'd6211,17'd6212,17'd5913,17'd5913,17'd5915,17'd6213,17'd6214,17'd6214,17'd6215,17'd6215,17'd6215,17'd6215,17'd6216,17'd6216,17'd6216,17'd6216,17'd6217,17'd6217,17'd6216,17'd6216,17'd6216,17'd6215,17'd5917,17'd5916,17'd5916,17'd5916,17'd5332,17'd5332,17'd5332,17'd5332,17'd6218,17'd6218,17'd6219,17'd6219,17'd6220,17'd6220,17'd6221,17'd5919,17'd6222,17'd6222,17'd6223,17'd6224,17'd6224,17'd6069,17'd6225,17'd6226,17'd6227,17'd6228,17'd6229,17'd6230,17'd6231,17'd6232,17'd6233,17'd6234,17'd3856,17'd6079,17'd6235,17'd3869,17'd6236,17'd6237,17'd6238,17'd6239,17'd5497,17'd4712,17'd1119,17'd5050,17'd1668,17'd412,17'd2408,17'd5360,17'd2751,17'd3395,17'd5634,17'd6240,17'd3227,17'd6087,17'd5637,17'd5780,17'd5781,17'd5780,17'd6241,17'd6242,17'd3574,17'd5635,17'd6243,17'd6243,17'd6244,17'd6245,17'd6246,17'd6247,17'd3082,17'd4564,17'd6248,17'd2405,17'd2247,17'd3404,17'd6249,17'd6249,17'd2247,17'd6250,17'd6251,17'd6252,17'd5368,17'd5369,17'd4874,17'd6253,17'd5953,17'd3242,17'd5046,17'd5190,17'd6254,17'd5190,17'd5190,17'd5190,17'd6255,17'd6256,17'd5954,17'd6257,17'd5955,17'd4241,17'd3742,17'd3742,17'd2392,17'd2392,17'd5372,17'd5371,17'd4880,17'd5371,17'd4729,17'd4882,17'd5958,17'd5958,17'd6258,17'd6258,17'd6095,17'd4730,17'd6259,17'd2240,17'd3247,17'd228,17'd1399,17'd228,17'd2586,17'd2096,17'd4575,17'd3897,17'd3423,17'd2586,17'd2559,17'd2417,17'd1823,17'd1666,17'd259,17'd1243,17'd274,17'd269,17'd269,17'd270,17'd1828,17'd1098,17'd2117,17'd1246,17'd419,17'd198
},
'{
17'd14,17'd1127,17'd5196,17'd6260,17'd3904,17'd4244,17'd5201,17'd5377,17'd5792,17'd6261,17'd6262,17'd6262,17'd5643,17'd5790,17'd5645,17'd5197,17'd5792,17'd5960,17'd6263,17'd4888,17'd3902,17'd6264,17'd6265,17'd1689,17'd14,17'd1127,17'd2595,17'd4247,17'd1127,17'd1127,17'd1689,17'd1689,17'd1127,17'd1127,17'd1689,17'd1689,17'd1689,17'd1689,17'd1127,17'd14,17'd2,17'd12,17'd11,17'd21,17'd4,17'd5,17'd3753,17'd3753,17'd6,17'd6,17'd3753,17'd3753,17'd3753,17'd6,17'd6,17'd1413,17'd6098,17'd6266,17'd5965,17'd6101,17'd6267,17'd6268,17'd6269,17'd6270,17'd6271,17'd6272,17'd6273,17'd6274,17'd6275,17'd5799,17'd6276,17'd6277,17'd25,17'd23,17'd22,17'd284,17'd24,17'd24,17'd284,17'd22,17'd22,17'd21,17'd27,17'd27,17'd28,17'd652,17'd4091,17'd3595,17'd3595,17'd3595,17'd3910,17'd6278,17'd5971,17'd5971,17'd5971,17'd5971,17'd5973,17'd5973,17'd5803,17'd5803,17'd5803,17'd5803,17'd5803,17'd5803,17'd6279,17'd6279,17'd6280,17'd6112,17'd6281,17'd6282,17'd6282,17'd5979,17'd5223,17'd6283,17'd6284,17'd5665,17'd5815,17'd4098,17'd6285,17'd6286,17'd6287,17'd5392,17'd5393,17'd6288,17'd6289,17'd6290,17'd6291,17'd6292,17'd6293,17'd6294,17'd6295,17'd6296,17'd6129,17'd6297,17'd6298,17'd6299,17'd6133,17'd6300,17'd6301,17'd6302,17'd5836,17'd6303,17'd6304,17'd6138,17'd6305,17'd6140,17'd6141,17'd6141,17'd6141,17'd6142,17'd6142,17'd6142,17'd6143,17'd5837,17'd5409,17'd5090,17'd4926,17'd6306,17'd4127,17'd3951,17'd3784,17'd3784,17'd3949,17'd6307,17'd5838,17'd5838,17'd5839,17'd3470,17'd6308,17'd6309,17'd6310,17'd6144,17'd6144,17'd6144,17'd6144,17'd5843,17'd6144,17'd6004,17'd6149,17'd6311,17'd6312,17'd6313,17'd6314,17'd6315,17'd5839,17'd6316,17'd6317,17'd6318,17'd6319,17'd6320,17'd6321,17'd6322,17'd6323,17'd6324,17'd6325,17'd6326,17'd6327,17'd6328,17'd6160,17'd6329,17'd6330,17'd6331,17'd6332,17'd6333,17'd6334,17'd6335,17'd6336,17'd6337,17'd6338,17'd6339,17'd6340,17'd6341,17'd6342,17'd6343,17'd6344,17'd6345,17'd6346,17'd6347,17'd6348,17'd6349,17'd6350,17'd6351,17'd6352,17'd6353,17'd6354,17'd6355,17'd6356,17'd6357,17'd6358,17'd6359,17'd6360,17'd6361,17'd6362,17'd6363,17'd6364,17'd6365,17'd6366,17'd6367,17'd6368,17'd1044,17'd6198,17'd6198,17'd3025,17'd1197,17'd1197,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd134,17'd132,17'd3168,17'd6369,17'd6370,17'd6371,17'd6372,17'd6373,17'd6374,17'd6375,17'd6376,17'd6377,17'd6378,17'd6207,17'd6379,17'd6380,17'd4677,17'd6381,17'd5607,17'd5325,17'd4993,17'd4993,17'd4994,17'd5326,17'd6382,17'd6383,17'd6384,17'd6384,17'd6213,17'd6213,17'd6214,17'd6215,17'd6215,17'd6215,17'd6215,17'd6215,17'd6216,17'd6215,17'd6216,17'd6216,17'd6217,17'd6217,17'd6385,17'd6386,17'd6216,17'd6216,17'd5917,17'd5917,17'd5916,17'd5915,17'd5761,17'd5331,17'd6387,17'd6388,17'd6218,17'd6389,17'd6390,17'd6219,17'd6220,17'd6391,17'd6392,17'd6391,17'd6222,17'd6222,17'd6393,17'd6393,17'd6224,17'd6394,17'd6395,17'd6396,17'd6397,17'd6227,17'd6398,17'd6399,17'd6400,17'd6401,17'd6075,17'd6233,17'd6234,17'd3857,17'd6402,17'd6403,17'd4054,17'd6404,17'd6405,17'd6406,17'd4228,17'd3745,17'd2777,17'd2392,17'd6407,17'd2409,17'd2098,17'd5498,17'd2574,17'd2913,17'd5633,17'd5634,17'd3228,17'd3227,17'd5780,17'd5780,17'd5781,17'd5781,17'd6408,17'd6242,17'd3574,17'd5366,17'd4407,17'd6243,17'd6243,17'd6409,17'd6245,17'd6247,17'd3082,17'd2405,17'd3082,17'd4409,17'd3404,17'd2248,17'd4563,17'd4063,17'd3404,17'd2248,17'd6251,17'd3884,17'd6410,17'd5368,17'd6089,17'd4874,17'd4876,17'd5953,17'd3417,17'd5046,17'd5190,17'd6255,17'd6254,17'd5190,17'd6254,17'd6411,17'd6412,17'd6413,17'd6414,17'd5955,17'd5956,17'd5192,17'd1810,17'd1810,17'd6415,17'd5371,17'd4880,17'd4880,17'd4729,17'd4882,17'd5958,17'd6416,17'd6417,17'd6418,17'd6094,17'd6258,17'd4730,17'd6259,17'd4575,17'd3247,17'd1399,17'd1260,17'd2586,17'd2096,17'd4575,17'd4575,17'd3897,17'd3246,17'd2392,17'd2417,17'd2417,17'd1666,17'd260,17'd1243,17'd458,17'd269,17'd269,17'd270,17'd1828,17'd1686,17'd2117,17'd421,17'd198,17'd198
},
'{
17'd6419,17'd4576,17'd6260,17'd6420,17'd4891,17'd4426,17'd6421,17'd6422,17'd5510,17'd6423,17'd6423,17'd6422,17'd5643,17'd5198,17'd6263,17'd5376,17'd5959,17'd5959,17'd5645,17'd4087,17'd3751,17'd6424,17'd2781,17'd1967,17'd1127,17'd4247,17'd4247,17'd1127,17'd14,17'd1967,17'd1689,17'd1688,17'd1689,17'd1689,17'd1689,17'd1689,17'd1689,17'd1689,17'd1127,17'd1127,17'd2,17'd3,17'd808,17'd9,17'd8,17'd6,17'd3753,17'd5793,17'd3753,17'd3594,17'd3594,17'd5205,17'd6,17'd5,17'd6425,17'd6426,17'd6427,17'd6428,17'd6102,17'd6268,17'd6269,17'd6429,17'd6430,17'd6431,17'd6432,17'd6270,17'd6433,17'd6267,17'd6434,17'd6435,17'd6436,17'd5650,17'd5647,17'd8,17'd4,17'd4,17'd23,17'd22,17'd22,17'd22,17'd1832,17'd285,17'd286,17'd27,17'd653,17'd653,17'd4091,17'd4091,17'd3755,17'd3755,17'd5971,17'd5971,17'd6437,17'd6437,17'd6437,17'd6438,17'd5803,17'd5803,17'd5803,17'd5803,17'd5803,17'd5972,17'd5972,17'd6439,17'd6440,17'd6441,17'd6113,17'd6282,17'd6282,17'd6281,17'd6442,17'd6443,17'd5222,17'd6444,17'd6284,17'd5063,17'd6445,17'd6446,17'd6447,17'd6448,17'd5230,17'd6449,17'd6450,17'd6451,17'd6452,17'd6453,17'd6454,17'd6455,17'd6456,17'd6457,17'd6458,17'd6459,17'd6460,17'd6461,17'd6299,17'd6462,17'd6301,17'd6463,17'd6463,17'd6464,17'd6465,17'd6465,17'd6305,17'd6305,17'd6466,17'd6467,17'd6140,17'd6468,17'd6141,17'd6141,17'd6141,17'd6141,17'd5409,17'd5409,17'd5090,17'd4926,17'd4926,17'd4127,17'd3952,17'd6469,17'd6470,17'd3629,17'd3949,17'd3949,17'd6471,17'd3626,17'd5839,17'd3470,17'd2985,17'd2985,17'd5842,17'd5842,17'd5842,17'd5842,17'd5842,17'd5842,17'd5842,17'd6472,17'd6312,17'd6313,17'd6473,17'd6473,17'd6474,17'd6475,17'd6476,17'd6477,17'd6478,17'd6479,17'd6480,17'd6481,17'd6482,17'd6483,17'd6484,17'd6485,17'd6486,17'd6487,17'd6488,17'd6159,17'd6489,17'd6490,17'd6491,17'd6492,17'd6493,17'd6494,17'd6495,17'd6496,17'd6497,17'd6498,17'd6499,17'd6500,17'd6501,17'd6502,17'd6503,17'd6504,17'd6505,17'd6506,17'd6507,17'd6508,17'd6509,17'd6510,17'd6511,17'd6512,17'd6513,17'd6514,17'd6515,17'd6516,17'd6517,17'd6518,17'd6519,17'd6520,17'd6521,17'd6522,17'd6523,17'd6524,17'd6525,17'd6526,17'd6527,17'd6528,17'd6368,17'd6529,17'd6530,17'd6198,17'd719,17'd542,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd133,17'd133,17'd132,17'd131,17'd6531,17'd6532,17'd6533,17'd6534,17'd6535,17'd6536,17'd6537,17'd6538,17'd6539,17'd6540,17'd6541,17'd6542,17'd6209,17'd4677,17'd6543,17'd6544,17'd6545,17'd6546,17'd6547,17'd6548,17'd6549,17'd5913,17'd5914,17'd5914,17'd6384,17'd6384,17'd6215,17'd6550,17'd6550,17'd6550,17'd6550,17'd6550,17'd6550,17'd6550,17'd6550,17'd6386,17'd6386,17'd6386,17'd6386,17'd6385,17'd6385,17'd6551,17'd6215,17'd6215,17'd6214,17'd6213,17'd6213,17'd5915,17'd6552,17'd6552,17'd5332,17'd6388,17'd6553,17'd6553,17'd6390,17'd6554,17'd6219,17'd6220,17'd6222,17'd6555,17'd6556,17'd6557,17'd6558,17'd6558,17'd6559,17'd6560,17'd6561,17'd6562,17'd6563,17'd6564,17'd4541,17'd6565,17'd6566,17'd6567,17'd6568,17'd6569,17'd6233,17'd6570,17'd4218,17'd6571,17'd6572,17'd3869,17'd5025,17'd6405,17'd3071,17'd447,17'd626,17'd625,17'd445,17'd4085,17'd2393,17'd1383,17'd5359,17'd4231,17'd2913,17'd3876,17'd3228,17'd3227,17'd3227,17'd5779,17'd6573,17'd6408,17'd6574,17'd5779,17'd5503,17'd5366,17'd5501,17'd6575,17'd6576,17'd6577,17'd6244,17'd5947,17'd4564,17'd4564,17'd3404,17'd4563,17'd6249,17'd2247,17'd3716,17'd3402,17'd4064,17'd4064,17'd2248,17'd2754,17'd6251,17'd6578,17'd5505,17'd5186,17'd6579,17'd5187,17'd5642,17'd3242,17'd5190,17'd6255,17'd6580,17'd5190,17'd5190,17'd5048,17'd4725,17'd4876,17'd6412,17'd4237,17'd3889,17'd3585,17'd5192,17'd3742,17'd1810,17'd4422,17'd6415,17'd5372,17'd5371,17'd5372,17'd3073,17'd6581,17'd6258,17'd6418,17'd6094,17'd6258,17'd4730,17'd6582,17'd6259,17'd4575,17'd2586,17'd228,17'd228,17'd3247,17'd6259,17'd4575,17'd3425,17'd3246,17'd1119,17'd2392,17'd2559,17'd1262,17'd970,17'd970,17'd273,17'd272,17'd640,17'd269,17'd1687,17'd1098,17'd2116,17'd1246,17'd419,17'd198
},
'{
17'd6583,17'd6260,17'd6584,17'd4892,17'd4426,17'd4735,17'd5790,17'd6585,17'd6586,17'd6423,17'd6423,17'd6586,17'd5510,17'd5643,17'd5959,17'd5645,17'd6263,17'd5197,17'd4735,17'd4427,17'd2783,17'd2592,17'd1967,17'd1967,17'd4247,17'd1127,17'd1127,17'd1127,17'd1689,17'd1689,17'd1689,17'd1689,17'd1689,17'd1689,17'd1689,17'd1689,17'd1689,17'd1127,17'd14,17'd2,17'd12,17'd806,17'd25,17'd4,17'd6,17'd3753,17'd5793,17'd5793,17'd3753,17'd3753,17'd3753,17'd6,17'd6,17'd8,17'd6587,17'd6588,17'd6435,17'd6589,17'd6268,17'd6269,17'd6590,17'd6591,17'd6592,17'd6593,17'd6591,17'd6594,17'd6269,17'd6595,17'd6105,17'd6596,17'd6597,17'd5794,17'd5647,17'd5647,17'd8,17'd4,17'd23,17'd23,17'd23,17'd22,17'd285,17'd285,17'd27,17'd980,17'd653,17'd653,17'd4091,17'd4091,17'd4431,17'd4431,17'd5971,17'd6598,17'd6437,17'd6437,17'd6437,17'd6437,17'd5803,17'd5803,17'd5803,17'd5973,17'd5972,17'd6599,17'd6599,17'd6600,17'd6601,17'd6601,17'd6602,17'd6602,17'd6282,17'd6281,17'd6443,17'd5385,17'd5524,17'd6114,17'd6603,17'd6604,17'd6605,17'd6606,17'd6607,17'd6608,17'd6609,17'd6610,17'd6611,17'd6612,17'd6613,17'd6614,17'd6615,17'd6616,17'd6617,17'd6618,17'd6619,17'd6620,17'd6621,17'd6299,17'd6622,17'd6623,17'd5836,17'd5836,17'd6464,17'd6464,17'd6465,17'd6624,17'd6625,17'd6625,17'd6466,17'd6467,17'd6626,17'd6626,17'd6141,17'd6141,17'd6141,17'd5837,17'd5409,17'd5255,17'd4925,17'd6627,17'd4127,17'd6628,17'd6628,17'd3951,17'd3784,17'd3784,17'd3949,17'd6629,17'd6630,17'd3781,17'd3470,17'd3470,17'd3468,17'd3468,17'd5842,17'd5842,17'd5842,17'd6631,17'd6472,17'd6472,17'd6150,17'd6312,17'd6313,17'd6632,17'd6633,17'd6634,17'd6635,17'd6636,17'd6637,17'd6638,17'd6639,17'd6633,17'd6640,17'd6641,17'd6642,17'd6643,17'd6644,17'd6645,17'd6646,17'd6647,17'd6648,17'd6649,17'd6650,17'd6651,17'd6652,17'd6653,17'd6654,17'd6655,17'd6656,17'd6657,17'd6658,17'd6659,17'd6660,17'd6661,17'd6662,17'd6663,17'd6664,17'd6665,17'd6666,17'd6667,17'd6668,17'd6669,17'd6670,17'd6671,17'd6672,17'd6673,17'd6674,17'd6675,17'd6676,17'd6677,17'd6678,17'd6679,17'd6680,17'd6681,17'd6682,17'd6683,17'd6684,17'd6685,17'd6686,17'd6687,17'd6688,17'd6689,17'd6690,17'd6368,17'd3167,17'd6198,17'd719,17'd542,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd1197,17'd1197,17'd132,17'd357,17'd6691,17'd6692,17'd6693,17'd6694,17'd6695,17'd6696,17'd6697,17'd6698,17'd6699,17'd6700,17'd6701,17'd6380,17'd4677,17'd4679,17'd6702,17'd6545,17'd6547,17'd6211,17'd6548,17'd6549,17'd5913,17'd5914,17'd5914,17'd6384,17'd6384,17'd6703,17'd6550,17'd6550,17'd6550,17'd6550,17'd6550,17'd6550,17'd6550,17'd6550,17'd6550,17'd6550,17'd6550,17'd6386,17'd6550,17'd6386,17'd6386,17'd6385,17'd6386,17'd6216,17'd6215,17'd6215,17'd6215,17'd6215,17'd5918,17'd6704,17'd6705,17'd6706,17'd6707,17'd6707,17'd6390,17'd6390,17'd6390,17'd6390,17'd6708,17'd6222,17'd6557,17'd6557,17'd6557,17'd6557,17'd6709,17'd6710,17'd6711,17'd6712,17'd6713,17'd5923,17'd4540,17'd4541,17'd6073,17'd6714,17'd6715,17'd6716,17'd6717,17'd4041,17'd6078,17'd4218,17'd6718,17'd6719,17'd4393,17'd5933,17'd6720,17'd451,17'd2587,17'd623,17'd625,17'd3247,17'd6415,17'd2393,17'd6721,17'd5942,17'd6722,17'd3395,17'd5634,17'd3227,17'd6087,17'd5779,17'd5636,17'd5636,17'd6723,17'd6574,17'd5185,17'd5779,17'd5502,17'd5365,17'd6724,17'd6576,17'd6577,17'd6244,17'd4564,17'd3082,17'd6249,17'd4563,17'd4563,17'd3404,17'd3403,17'd3403,17'd4064,17'd4720,17'd2247,17'd2248,17'd3084,17'd2757,17'd6725,17'd6725,17'd5950,17'd4875,17'd5784,17'd5642,17'd3417,17'd6255,17'd6580,17'd6580,17'd6255,17'd6254,17'd6091,17'd5784,17'd5187,17'd6412,17'd4237,17'd5955,17'd6726,17'd5788,17'd4422,17'd4422,17'd1946,17'd6415,17'd5371,17'd5371,17'd5940,17'd6727,17'd6094,17'd6418,17'd6094,17'd6258,17'd5789,17'd5789,17'd5789,17'd6259,17'd3897,17'd2586,17'd1119,17'd2586,17'd4575,17'd4575,17'd4883,17'd3896,17'd3246,17'd3247,17'd2392,17'd1680,17'd1396,17'd1243,17'd273,17'd273,17'd640,17'd269,17'd1687,17'd1098,17'd2116,17'd1246,17'd419,17'd198
},
'{
17'd6728,17'd3904,17'd4244,17'd4087,17'd5200,17'd6421,17'd6422,17'd6585,17'd6586,17'd6729,17'd6423,17'd6586,17'd5510,17'd5790,17'd5959,17'd5197,17'd6263,17'd4734,17'd6730,17'd3751,17'd2784,17'd2781,17'd1967,17'd14,17'd4247,17'd1127,17'd14,17'd14,17'd1688,17'd1688,17'd5196,17'd4576,17'd2781,17'd2781,17'd1689,17'd1689,17'd1127,17'd1127,17'd2,17'd13,17'd3,17'd1275,17'd9,17'd8,17'd6,17'd3753,17'd5793,17'd5793,17'd3753,17'd3753,17'd7,17'd6,17'd8,17'd5512,17'd6731,17'd6732,17'd6589,17'd6733,17'd6734,17'd6735,17'd6736,17'd6737,17'd6738,17'd6738,17'd6739,17'd6740,17'd6741,17'd6742,17'd6105,17'd6732,17'd6743,17'd5648,17'd5647,17'd5206,17'd8,17'd4,17'd4,17'd23,17'd25,17'd25,17'd285,17'd26,17'd27,17'd980,17'd653,17'd653,17'd4430,17'd4430,17'd6744,17'd6744,17'd6437,17'd6437,17'd6437,17'd6437,17'd6745,17'd6437,17'd6746,17'd6746,17'd5972,17'd6439,17'd6599,17'd6600,17'd6747,17'd6748,17'd6749,17'd6749,17'd6750,17'd6602,17'd5979,17'd5979,17'd5813,17'd5385,17'd5386,17'd6751,17'd6752,17'd6753,17'd6754,17'd6755,17'd6756,17'd6757,17'd6758,17'd6759,17'd6760,17'd6761,17'd6762,17'd6125,17'd6616,17'd6763,17'd6764,17'd6765,17'd6766,17'd6460,17'd6767,17'd6768,17'd6622,17'd6464,17'd6465,17'd6465,17'd6465,17'd6624,17'd6625,17'd6769,17'd6770,17'd6770,17'd6141,17'd6140,17'd6626,17'd6626,17'd6141,17'd6141,17'd5689,17'd5689,17'd5255,17'd4925,17'd4926,17'd6306,17'd3952,17'd6628,17'd6628,17'd6771,17'd4923,17'd3950,17'd6772,17'd3949,17'd6471,17'd3626,17'd5839,17'd3470,17'd5840,17'd5841,17'd5841,17'd6152,17'd5841,17'd6773,17'd6774,17'd6316,17'd6775,17'd6776,17'd6776,17'd6777,17'd6635,17'd6778,17'd6778,17'd6779,17'd6779,17'd6780,17'd6781,17'd6782,17'd6783,17'd6784,17'd6785,17'd6786,17'd6787,17'd6645,17'd6788,17'd6789,17'd6790,17'd6791,17'd6792,17'd6793,17'd6794,17'd6795,17'd6796,17'd6797,17'd6798,17'd6799,17'd6800,17'd6801,17'd6802,17'd6803,17'd6804,17'd6805,17'd6806,17'd6807,17'd6808,17'd6809,17'd6810,17'd6811,17'd6812,17'd6813,17'd6814,17'd6815,17'd6816,17'd6817,17'd6818,17'd6819,17'd6820,17'd6821,17'd6822,17'd6823,17'd6824,17'd6825,17'd6826,17'd6827,17'd6686,17'd6687,17'd6688,17'd6689,17'd6828,17'd6829,17'd6830,17'd888,17'd542,17'd542,17'd542,17'd542,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd135,17'd132,17'd132,17'd135,17'd5593,17'd6831,17'd4976,17'd3347,17'd6832,17'd6833,17'd6834,17'd6538,17'd6835,17'd6836,17'd6837,17'd6838,17'd6839,17'd6840,17'd6543,17'd6544,17'd6545,17'd6841,17'd6842,17'd6843,17'd6844,17'd6845,17'd6846,17'd6846,17'd6703,17'd6703,17'd6847,17'd6847,17'd6848,17'd6848,17'd6848,17'd6848,17'd6848,17'd6848,17'd6848,17'd6849,17'd6849,17'd6849,17'd6849,17'd6849,17'd6849,17'd6849,17'd6386,17'd6386,17'd6386,17'd6386,17'd6386,17'd6216,17'd6217,17'd6850,17'd6705,17'd6851,17'd6851,17'd6852,17'd6707,17'd6220,17'd6219,17'd6390,17'd6390,17'd6853,17'd6223,17'd6558,17'd6557,17'd6854,17'd6854,17'd6855,17'd6710,17'd6711,17'd6856,17'd6857,17'd6858,17'd6859,17'd6860,17'd6228,17'd6073,17'd6861,17'd6400,17'd6862,17'd6863,17'd6864,17'd6078,17'd4218,17'd6865,17'd3563,17'd6866,17'd6083,17'd6867,17'd235,17'd447,17'd1825,17'd1119,17'd6407,17'd6868,17'd2575,17'd2408,17'd3393,17'd2914,17'd3876,17'd3573,17'd3399,17'd3877,17'd5502,17'd6869,17'd6870,17'd6870,17'd6574,17'd6574,17'd5502,17'd5365,17'd6871,17'd6872,17'd6873,17'd6577,17'd6245,17'd5037,17'd3082,17'd4564,17'd5946,17'd4720,17'd3402,17'd3403,17'd3402,17'd4232,17'd6249,17'd3404,17'd2760,17'd2757,17'd6874,17'd6875,17'd6876,17'd5640,17'd6877,17'd6878,17'd4726,17'd5048,17'd6580,17'd6879,17'd6880,17'd6255,17'd6580,17'd6411,17'd6881,17'd6882,17'd6883,17'd5786,17'd6257,17'd6884,17'd6885,17'd6886,17'd6887,17'd6888,17'd5372,17'd4880,17'd5372,17'd6889,17'd6416,17'd6890,17'd6890,17'd6094,17'd6094,17'd6891,17'd5789,17'd6259,17'd6259,17'd3897,17'd445,17'd1261,17'd3391,17'd4423,17'd4882,17'd4713,17'd3897,17'd3247,17'd2392,17'd2417,17'd1823,17'd1243,17'd641,17'd409,17'd640,17'd269,17'd643,17'd1685,17'd2116,17'd1246,17'd419,17'd416
},
'{
17'd6892,17'd4244,17'd4426,17'd4735,17'd6421,17'd5643,17'd6422,17'd6585,17'd6893,17'd6729,17'd6423,17'd6423,17'd6422,17'd5510,17'd5959,17'd5509,17'd4888,17'd5646,17'd4086,17'd2782,17'd2781,17'd1967,17'd14,17'd1127,17'd1127,17'd1127,17'd14,17'd1689,17'd1688,17'd1688,17'd5196,17'd5196,17'd3250,17'd3250,17'd1689,17'd1689,17'd1127,17'd466,17'd13,17'd2423,17'd1275,17'd2591,17'd4,17'd6,17'd3753,17'd3753,17'd5793,17'd5793,17'd3753,17'd3753,17'd6,17'd8,17'd5647,17'd5648,17'd6099,17'd6434,17'd6268,17'd6429,17'd6593,17'd6894,17'd6738,17'd6895,17'd6896,17'd6896,17'd6894,17'd6897,17'd6898,17'd6899,17'd6105,17'd6900,17'd6901,17'd5794,17'd5647,17'd8,17'd8,17'd4,17'd4,17'd23,17'd25,17'd25,17'd26,17'd26,17'd980,17'd980,17'd652,17'd652,17'd6744,17'd6744,17'd6902,17'd6902,17'd6903,17'd6437,17'd6437,17'd6437,17'd6745,17'd6745,17'd5972,17'd6439,17'd6439,17'd6904,17'd6600,17'd6747,17'd6905,17'd6905,17'd6906,17'd6907,17'd6750,17'd6602,17'd5979,17'd5979,17'd5813,17'd5386,17'd6908,17'd6909,17'd6910,17'd6911,17'd6912,17'd6913,17'd6914,17'd6915,17'd6916,17'd6917,17'd6918,17'd6919,17'd6920,17'd6921,17'd6922,17'd6923,17'd6924,17'd6925,17'd6926,17'd6927,17'd6928,17'd6929,17'd6930,17'd6465,17'd6465,17'd6465,17'd6624,17'd6624,17'd6769,17'd6769,17'd6931,17'd6770,17'd6141,17'd6140,17'd6626,17'd6626,17'd6141,17'd5689,17'd5255,17'd5255,17'd4926,17'd4926,17'd6306,17'd6932,17'd6628,17'd6628,17'd6771,17'd6771,17'd6933,17'd6934,17'd6772,17'd6629,17'd3626,17'd5838,17'd5839,17'd3297,17'd5840,17'd5840,17'd5841,17'd6935,17'd6773,17'd6936,17'd6776,17'd6475,17'd6474,17'd6475,17'd6777,17'd6937,17'd6778,17'd6938,17'd6779,17'd6939,17'd6940,17'd6941,17'd6942,17'd6943,17'd6944,17'd6945,17'd6946,17'd6947,17'd6948,17'd6949,17'd6950,17'd6951,17'd6952,17'd6953,17'd6954,17'd6955,17'd6956,17'd6957,17'd6958,17'd6959,17'd6960,17'd6961,17'd6962,17'd6963,17'd6964,17'd6965,17'd6966,17'd6967,17'd6968,17'd6969,17'd6970,17'd6971,17'd6972,17'd6973,17'd6974,17'd6975,17'd6976,17'd6977,17'd6978,17'd6979,17'd6980,17'd6818,17'd6981,17'd6982,17'd6983,17'd6984,17'd6985,17'd6986,17'd6987,17'd6988,17'd6686,17'd6364,17'd6989,17'd6990,17'd6991,17'd6992,17'd6993,17'd6830,17'd542,17'd542,17'd542,17'd542,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd5898,17'd132,17'd132,17'd357,17'd6531,17'd6994,17'd6995,17'd6996,17'd6997,17'd6998,17'd6999,17'd7000,17'd7001,17'd7002,17'd7003,17'd7004,17'd7005,17'd7006,17'd6702,17'd7007,17'd7008,17'd6841,17'd7009,17'd6845,17'd6845,17'd6846,17'd6703,17'd6703,17'd6703,17'd6847,17'd6847,17'd6848,17'd6848,17'd6848,17'd6848,17'd6848,17'd6848,17'd6848,17'd6848,17'd7010,17'd7010,17'd7010,17'd7010,17'd7010,17'd6849,17'd7010,17'd7010,17'd6386,17'd6386,17'd6386,17'd6385,17'd6217,17'd6217,17'd6850,17'd6850,17'd6705,17'd6705,17'd6707,17'd6852,17'd6391,17'd6391,17'd6220,17'd6219,17'd6708,17'd6223,17'd7011,17'd6558,17'd6854,17'd7012,17'd7013,17'd6855,17'd6711,17'd7014,17'd7015,17'd7016,17'd7017,17'd6859,17'd6860,17'd6228,17'd6566,17'd6567,17'd7018,17'd7019,17'd7020,17'd7021,17'd6234,17'd7022,17'd7023,17'd7024,17'd7025,17'd7026,17'd6084,17'd1121,17'd795,17'd625,17'd2417,17'd5957,17'd2905,17'd7027,17'd4560,17'd3393,17'd4715,17'd3573,17'd3573,17'd4233,17'd5501,17'd5365,17'd5502,17'd6869,17'd6723,17'd6574,17'd6869,17'd6869,17'd7028,17'd6872,17'd7029,17'd7030,17'd6409,17'd6245,17'd3082,17'd3082,17'd4720,17'd7031,17'd4404,17'd3402,17'd3402,17'd3575,17'd4563,17'd6249,17'd2759,17'd2756,17'd6874,17'd3883,17'd7032,17'd7033,17'd7034,17'd6877,17'd7035,17'd5048,17'd5952,17'd7036,17'd7037,17'd6879,17'd6580,17'd6880,17'd7038,17'd7039,17'd7040,17'd4724,17'd6413,17'd6257,17'd6093,17'd7041,17'd6887,17'd6887,17'd1946,17'd5372,17'd5371,17'd4423,17'd5789,17'd6094,17'd6890,17'd6094,17'd6094,17'd6094,17'd6094,17'd5789,17'd5789,17'd6259,17'd3391,17'd1261,17'd3895,17'd4423,17'd4882,17'd4882,17'd4575,17'd3423,17'd3391,17'd2392,17'd5050,17'd1396,17'd970,17'd409,17'd269,17'd640,17'd206,17'd645,17'd1409,17'd1246,17'd419,17'd416
},
'{
17'd7042,17'd5202,17'd4734,17'd5197,17'd6421,17'd5643,17'd7043,17'd7044,17'd7045,17'd7045,17'd6423,17'd7046,17'd5375,17'd5375,17'd7047,17'd7048,17'd7049,17'd5204,17'd2934,17'd2592,17'd1967,17'd14,17'd1127,17'd466,17'd14,17'd1127,17'd1689,17'd1689,17'd1689,17'd2781,17'd4886,17'd4886,17'd3250,17'd3250,17'd1688,17'd1688,17'd4247,17'd466,17'd13,17'd806,17'd2591,17'd2421,17'd6,17'd3753,17'd3753,17'd3753,17'd5793,17'd5793,17'd3753,17'd3753,17'd6,17'd5206,17'd7050,17'd6588,17'd6435,17'd6106,17'd6270,17'd7051,17'd6737,17'd7052,17'd7053,17'd7053,17'd6896,17'd7052,17'd6737,17'd7054,17'd7055,17'd7056,17'd7057,17'd7058,17'd7059,17'd5512,17'd8,17'd6,17'd5,17'd5,17'd1691,17'd1691,17'd467,17'd285,17'd286,17'd27,17'd980,17'd980,17'd980,17'd27,17'd7060,17'd7061,17'd7061,17'd7061,17'd6745,17'd6745,17'd6745,17'd6745,17'd6745,17'd6745,17'd7062,17'd6599,17'd6904,17'd6600,17'd6747,17'd7063,17'd7063,17'd7063,17'd6907,17'd7064,17'd6750,17'd7065,17'd7066,17'd7066,17'd7067,17'd7067,17'd7068,17'd7069,17'd7070,17'd7071,17'd7072,17'd7073,17'd6915,17'd6759,17'd7074,17'd6918,17'd6291,17'd7075,17'd7076,17'd7077,17'd7078,17'd7079,17'd6925,17'd7080,17'd7081,17'd7082,17'd7083,17'd7084,17'd6624,17'd7085,17'd7085,17'd6625,17'd6625,17'd6769,17'd7086,17'd7086,17'd7087,17'd7087,17'd6141,17'd6468,17'd5409,17'd5409,17'd5255,17'd5255,17'd5255,17'd4926,17'd7088,17'd7088,17'd3952,17'd3952,17'd6628,17'd6628,17'd6628,17'd5085,17'd6933,17'd7089,17'd7090,17'd6307,17'd5838,17'd5838,17'd6773,17'd6773,17'd6935,17'd7091,17'd6773,17'd7092,17'd3626,17'd7093,17'd7094,17'd7095,17'd7096,17'd7097,17'd7098,17'd7098,17'd7098,17'd7099,17'd7100,17'd7101,17'd7102,17'd7103,17'd7104,17'd7105,17'd7106,17'd7107,17'd7108,17'd7109,17'd7110,17'd7111,17'd7112,17'd7113,17'd7114,17'd7115,17'd7116,17'd7117,17'd7118,17'd7119,17'd7120,17'd7121,17'd7122,17'd7123,17'd7124,17'd7125,17'd7126,17'd7127,17'd7128,17'd7129,17'd7130,17'd7131,17'd7132,17'd7133,17'd7134,17'd7135,17'd7136,17'd7137,17'd7138,17'd7139,17'd7140,17'd7141,17'd7142,17'd7143,17'd7144,17'd7145,17'd7146,17'd7147,17'd7148,17'd7149,17'd7150,17'd7151,17'd6524,17'd7152,17'd7153,17'd6527,17'd7154,17'd6828,17'd7155,17'd6993,17'd888,17'd717,17'd542,17'd542,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd1759,17'd132,17'd131,17'd131,17'd4815,17'd4344,17'd7156,17'd7157,17'd3670,17'd6375,17'd7158,17'd7001,17'd7159,17'd7160,17'd7161,17'd6839,17'd7162,17'd6544,17'd7163,17'd7164,17'd7165,17'd7009,17'd7166,17'd7167,17'd7167,17'd7168,17'd7168,17'd7169,17'd7169,17'd7170,17'd7170,17'd7171,17'd7172,17'd7172,17'd7172,17'd7172,17'd7173,17'd7174,17'd7174,17'd7175,17'd7175,17'd7175,17'd7175,17'd6849,17'd6849,17'd6849,17'd6849,17'd6550,17'd6550,17'd6386,17'd6386,17'd6386,17'd6386,17'd7176,17'd7176,17'd6705,17'd6705,17'd6707,17'd6852,17'd6392,17'd6392,17'd6391,17'd6220,17'd7177,17'd7178,17'd7011,17'd7011,17'd6709,17'd7179,17'd7180,17'd7180,17'd7014,17'd7014,17'd7181,17'd7182,17'd7183,17'd7184,17'd7185,17'd6860,17'd4380,17'd6399,17'd7186,17'd7187,17'd4210,17'd7188,17'd7189,17'd5929,17'd7022,17'd7023,17'd7190,17'd7191,17'd6405,17'd3071,17'd1121,17'd428,17'd953,17'd1823,17'd6407,17'd2575,17'd2098,17'd2408,17'd7192,17'd3403,17'd4404,17'd5946,17'd6243,17'd7193,17'd4407,17'd4872,17'd7194,17'd7194,17'd6870,17'd6869,17'd5365,17'd6871,17'd7029,17'd6873,17'd7195,17'd7196,17'd4409,17'd3082,17'd4720,17'd7031,17'd4407,17'd4232,17'd7197,17'd3402,17'd4063,17'd4563,17'd3082,17'd2405,17'd4565,17'd4410,17'd7198,17'd7033,17'd7199,17'd7200,17'd6882,17'd6091,17'd4726,17'd7201,17'd7202,17'd7037,17'd7203,17'd7204,17'd7037,17'd6881,17'd7205,17'd7206,17'd4724,17'd6413,17'd7207,17'd7208,17'd4060,17'd4060,17'd7209,17'd7210,17'd6407,17'd5371,17'd4882,17'd5789,17'd6094,17'd6094,17'd6418,17'd6418,17'd6418,17'd6258,17'd5958,17'd7211,17'd4423,17'd3895,17'd3895,17'd4085,17'd4713,17'd4713,17'd4730,17'd3897,17'd3391,17'd1810,17'd5957,17'd1396,17'd970,17'd1243,17'd207,17'd258,17'd269,17'd645,17'd1409,17'd2117,17'd1528,17'd416
},
'{
17'd7212,17'd5645,17'd5197,17'd5959,17'd5643,17'd5643,17'd7043,17'd7043,17'd7045,17'd7213,17'd7046,17'd7046,17'd6262,17'd6262,17'd7047,17'd5509,17'd5203,17'd3901,17'd2784,17'd2781,17'd1967,17'd1127,17'd466,17'd466,17'd14,17'd1689,17'd1688,17'd1689,17'd2781,17'd2781,17'd4886,17'd7214,17'd2422,17'd3250,17'd1688,17'd1688,17'd1127,17'd13,17'd2423,17'd2933,17'd2421,17'd7215,17'd3753,17'd3753,17'd3753,17'd3753,17'd5793,17'd5793,17'd3753,17'd3753,17'd6,17'd7216,17'd6098,17'd6099,17'd6434,17'd6268,17'd7217,17'd7218,17'd6896,17'd6895,17'd7219,17'd7220,17'd6896,17'd7052,17'd7221,17'd6897,17'd6430,17'd6742,17'd7222,17'd7223,17'd7224,17'd1413,17'd8,17'd5,17'd5,17'd5,17'd1691,17'd1691,17'd467,17'd285,17'd286,17'd27,17'd27,17'd27,17'd27,17'd286,17'd7061,17'd7061,17'd7061,17'd7061,17'd6745,17'd6745,17'd6745,17'd6745,17'd6745,17'd7225,17'd7226,17'd7226,17'd6600,17'd6747,17'd7063,17'd7063,17'd7063,17'd7227,17'd7228,17'd6602,17'd7065,17'd7065,17'd7229,17'd7229,17'd7230,17'd7231,17'd6909,17'd6910,17'd6911,17'd7232,17'd7233,17'd7234,17'd7235,17'd7236,17'd7237,17'd7238,17'd7239,17'd6455,17'd7240,17'd7241,17'd7242,17'd7243,17'd7244,17'd7245,17'd7246,17'd7247,17'd7248,17'd6625,17'd7249,17'd7249,17'd6625,17'd6769,17'd6769,17'd7250,17'd7086,17'd7087,17'd7087,17'd7251,17'd6468,17'd6468,17'd5409,17'd5409,17'd5255,17'd5255,17'd4926,17'd7088,17'd7252,17'd7252,17'd3952,17'd3952,17'd6628,17'd6628,17'd4924,17'd4924,17'd6933,17'd7253,17'd7254,17'd7255,17'd7256,17'd5838,17'd6773,17'd6773,17'd7091,17'd7257,17'd6936,17'd6475,17'd6476,17'd6638,17'd7095,17'd7258,17'd7099,17'd7259,17'd7260,17'd7259,17'd7099,17'd7261,17'd7262,17'd7263,17'd7264,17'd7265,17'd7266,17'd7267,17'd7268,17'd7269,17'd7270,17'd7271,17'd7272,17'd7273,17'd7274,17'd7275,17'd7276,17'd7277,17'd7278,17'd7279,17'd7280,17'd7281,17'd7282,17'd7283,17'd7284,17'd7284,17'd7285,17'd7286,17'd7287,17'd7288,17'd7289,17'd7290,17'd7291,17'd7292,17'd7293,17'd7294,17'd7295,17'd7296,17'd7297,17'd7298,17'd7299,17'd7300,17'd7301,17'd7302,17'd7303,17'd7304,17'd7305,17'd7306,17'd7307,17'd7146,17'd7308,17'd7309,17'd7310,17'd7311,17'd7312,17'd7313,17'd7314,17'd6365,17'd7315,17'd7154,17'd6690,17'd7155,17'd6830,17'd888,17'd542,17'd542,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd3168,17'd5593,17'd7316,17'd7317,17'd7318,17'd7319,17'd7320,17'd7321,17'd7322,17'd7002,17'd7323,17'd6701,17'd6380,17'd7006,17'd7324,17'd7325,17'd7326,17'd7165,17'd7327,17'd7166,17'd7328,17'd7167,17'd7169,17'd7168,17'd7168,17'd7169,17'd7169,17'd7170,17'd7171,17'd7172,17'd7172,17'd7173,17'd7173,17'd7173,17'd7173,17'd7174,17'd7174,17'd7175,17'd7175,17'd7175,17'd7175,17'd6849,17'd7329,17'd7329,17'd6849,17'd6550,17'd6550,17'd6550,17'd6550,17'd6550,17'd6550,17'd7176,17'd7176,17'd6705,17'd6705,17'd6707,17'd6707,17'd6221,17'd6221,17'd6220,17'd6220,17'd7177,17'd7177,17'd7011,17'd7011,17'd6559,17'd6710,17'd7180,17'd7180,17'd7014,17'd7014,17'd7330,17'd7331,17'd7182,17'd7183,17'd7332,17'd7333,17'd7334,17'd7335,17'd7336,17'd7337,17'd7187,17'd6568,17'd7338,17'd7339,17'd5929,17'd4219,17'd7340,17'd4863,17'd6404,17'd7341,17'd243,17'd210,17'd428,17'd953,17'd2559,17'd2905,17'd1946,17'd2098,17'd7342,17'd1818,17'd6249,17'd7031,17'd6243,17'd6243,17'd4717,17'd7343,17'd7194,17'd7344,17'd7345,17'd6870,17'd5365,17'd7028,17'd7346,17'd7029,17'd7347,17'd7348,17'd7349,17'd4409,17'd4720,17'd7031,17'd4717,17'd4407,17'd5032,17'd3402,17'd4563,17'd4063,17'd4409,17'd4564,17'd4410,17'd4410,17'd7198,17'd7198,17'd7350,17'd7199,17'd7351,17'd7040,17'd7201,17'd7201,17'd7202,17'd7352,17'd7353,17'd7354,17'd7036,17'd7037,17'd7355,17'd7356,17'd7357,17'd7358,17'd7359,17'd7360,17'd7361,17'd7362,17'd7363,17'd7209,17'd7210,17'd2392,17'd4575,17'd4730,17'd6258,17'd6094,17'd6418,17'd7364,17'd6418,17'd6417,17'd7365,17'd5958,17'd4728,17'd4085,17'd3391,17'd3391,17'd4729,17'd4729,17'd4730,17'd4883,17'd4729,17'd4085,17'd5957,17'd3743,17'd1396,17'd1243,17'd271,17'd261,17'd640,17'd803,17'd1409,17'd1821,17'd1246,17'd416
},
'{
17'd5960,17'd5960,17'd5790,17'd6422,17'd6422,17'd6422,17'd7043,17'd7366,17'd7366,17'd7367,17'd7368,17'd6262,17'd7046,17'd7369,17'd7370,17'd5960,17'd4086,17'd2593,17'd7371,17'd3750,17'd1967,17'd1127,17'd466,17'd466,17'd1127,17'd1689,17'd1689,17'd2781,17'd2781,17'd3250,17'd7214,17'd7372,17'd2422,17'd3250,17'd1689,17'd1127,17'd466,17'd13,17'd1275,17'd2591,17'd2421,17'd7373,17'd3753,17'd3753,17'd5793,17'd5793,17'd3753,17'd3753,17'd3753,17'd3753,17'd7374,17'd7375,17'd6588,17'd6596,17'd6105,17'd7376,17'd6592,17'd6737,17'd6895,17'd7377,17'd7219,17'd7220,17'd7378,17'd7053,17'd6738,17'd6431,17'd6741,17'd7379,17'd7380,17'd7381,17'd5652,17'd8,17'd6,17'd3753,17'd7382,17'd7382,17'd7383,17'd7384,17'd1691,17'd467,17'd286,17'd286,17'd286,17'd286,17'd7385,17'd7385,17'd7385,17'd7385,17'd7385,17'd7385,17'd7386,17'd7387,17'd7225,17'd7225,17'd7225,17'd7388,17'd7389,17'd7389,17'd6748,17'd6905,17'd7390,17'd7390,17'd7227,17'd7391,17'd7392,17'd6282,17'd7393,17'd7393,17'd7229,17'd7230,17'd7230,17'd7231,17'd7069,17'd7394,17'd7395,17'd7396,17'd7397,17'd7398,17'd7399,17'd7400,17'd6613,17'd7401,17'd7402,17'd7403,17'd7404,17'd7405,17'd7406,17'd7407,17'd7081,17'd7408,17'd7409,17'd7410,17'd6770,17'd7411,17'd7411,17'd7412,17'd7412,17'd7413,17'd7413,17'd7413,17'd7414,17'd7415,17'd7416,17'd7417,17'd6468,17'd7418,17'd7418,17'd5409,17'd5090,17'd4767,17'd7088,17'd7252,17'd6932,17'd6932,17'd3952,17'd3952,17'd4127,17'd4127,17'd4127,17'd5250,17'd6933,17'd7253,17'd7254,17'd7255,17'd7256,17'd7256,17'd7092,17'd7419,17'd6314,17'd6314,17'd6475,17'd6777,17'd6637,17'd7420,17'd7421,17'd7099,17'd7422,17'd7422,17'd7422,17'd7422,17'd7423,17'd7424,17'd7425,17'd7426,17'd7427,17'd7428,17'd7429,17'd7430,17'd7431,17'd7432,17'd7433,17'd7434,17'd7435,17'd7436,17'd7437,17'd7438,17'd7439,17'd7440,17'd7441,17'd7442,17'd7443,17'd7444,17'd7445,17'd7446,17'd7447,17'd7448,17'd7449,17'd7450,17'd7451,17'd7452,17'd7453,17'd7454,17'd7455,17'd7456,17'd7457,17'd7458,17'd7459,17'd7460,17'd7461,17'd7462,17'd7463,17'd7464,17'd7465,17'd7466,17'd7467,17'd7468,17'd7469,17'd7470,17'd7471,17'd7472,17'd7473,17'd7474,17'd7475,17'd7476,17'd7477,17'd7478,17'd7479,17'd7480,17'd7481,17'd7482,17'd7483,17'd6368,17'd6830,17'd888,17'd719,17'd542,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd1197,17'd133,17'd3025,17'd3168,17'd7484,17'd7485,17'd7486,17'd7487,17'd7488,17'd5319,17'd7489,17'd7490,17'd7491,17'd6701,17'd7492,17'd7493,17'd6543,17'd6544,17'd7163,17'd7326,17'd7327,17'd7494,17'd7328,17'd7328,17'd7169,17'd7169,17'd6550,17'd6550,17'd6848,17'd6848,17'd7171,17'd7495,17'd7496,17'd7497,17'd7498,17'd7498,17'd7173,17'd7173,17'd7173,17'd7173,17'd7175,17'd7175,17'd7175,17'd7175,17'd6848,17'd6848,17'd6849,17'd6849,17'd6550,17'd6550,17'd6550,17'd6550,17'd6550,17'd6550,17'd6215,17'd6215,17'd7176,17'd6704,17'd6387,17'd6387,17'd5919,17'd5919,17'd5919,17'd6220,17'd7499,17'd7500,17'd6558,17'd6559,17'd7501,17'd7501,17'd6711,17'd7502,17'd7014,17'd7014,17'd7181,17'd7330,17'd7503,17'd7504,17'd7505,17'd7184,17'd7506,17'd7507,17'd7335,17'd6399,17'd4209,17'd7508,17'd7509,17'd7338,17'd7339,17'd7510,17'd5022,17'd7511,17'd5626,17'd7026,17'd784,17'd1093,17'd429,17'd7512,17'd1262,17'd5957,17'd6415,17'd2575,17'd4560,17'd2407,17'd2248,17'd4063,17'd6409,17'd6409,17'd6576,17'd7343,17'd7513,17'd7514,17'd7515,17'd7345,17'd7516,17'd7346,17'd7029,17'd7029,17'd7517,17'd7517,17'd7518,17'd7519,17'd7031,17'd7031,17'd6243,17'd7193,17'd7520,17'd7521,17'd5947,17'd4409,17'd7349,17'd7349,17'd3407,17'd3406,17'd6875,17'd7522,17'd7350,17'd7350,17'd7523,17'd7524,17'd7525,17'd7035,17'd7526,17'd7037,17'd7527,17'd7528,17'd7353,17'd7529,17'd7530,17'd7356,17'd7531,17'd6579,17'd7532,17'd7533,17'd7534,17'd7535,17'd7536,17'd7536,17'd7209,17'd6407,17'd1810,17'd6259,17'd5789,17'd6094,17'd7537,17'd7538,17'd7537,17'd6416,17'd5958,17'd5958,17'd7211,17'd4728,17'd4085,17'd3895,17'd3744,17'd4729,17'd6095,17'd4730,17'd4713,17'd4085,17'd6407,17'd4084,17'd190,17'd1243,17'd642,17'd256,17'd7539,17'd803,17'd1686,17'd1821,17'd1246,17'd601
},
'{
17'd6261,17'd7540,17'd7541,17'd5510,17'd6422,17'd5510,17'd7043,17'd7542,17'd7542,17'd7543,17'd7369,17'd6423,17'd7046,17'd7368,17'd7544,17'd5377,17'd3751,17'd2784,17'd2781,17'd1967,17'd1127,17'd4247,17'd466,17'd2,17'd4247,17'd1689,17'd3750,17'd3750,17'd2781,17'd2422,17'd7214,17'd7545,17'd3250,17'd3250,17'd1689,17'd1127,17'd2,17'd12,17'd2933,17'd2421,17'd7215,17'd7373,17'd3753,17'd3753,17'd5793,17'd5793,17'd3753,17'd3753,17'd6,17'd6,17'd7216,17'd5649,17'd6266,17'd5965,17'd6733,17'd7546,17'd6738,17'd7547,17'd7220,17'd7548,17'd7219,17'd7378,17'd7549,17'd7550,17'd6737,17'd6431,17'd7551,17'd7552,17'd6266,17'd7553,17'd5647,17'd5206,17'd6,17'd6,17'd7554,17'd7383,17'd7383,17'd7383,17'd1691,17'd1691,17'd285,17'd286,17'd286,17'd286,17'd7555,17'd7555,17'd7385,17'd7385,17'd7385,17'd7385,17'd7386,17'd7386,17'd7225,17'd7556,17'd7556,17'd7557,17'd7389,17'd7558,17'd6905,17'd7559,17'd7390,17'd7560,17'd7561,17'd7392,17'd7562,17'd7563,17'd6282,17'd7393,17'd7229,17'd7230,17'd7230,17'd7564,17'd7070,17'd7071,17'd7565,17'd7566,17'd7567,17'd7568,17'd7569,17'd6761,17'd7570,17'd6292,17'd7571,17'd7572,17'd7573,17'd7574,17'd7575,17'd7576,17'd7577,17'd7578,17'd7578,17'd6770,17'd7412,17'd7412,17'd7579,17'd7579,17'd7414,17'd7580,17'd7580,17'd7580,17'd7579,17'd7581,17'd7416,17'd7417,17'd6468,17'd5409,17'd5409,17'd7582,17'd4767,17'd4926,17'd7088,17'd7252,17'd7583,17'd3953,17'd3952,17'd4127,17'd4127,17'd4610,17'd4610,17'd5250,17'd6933,17'd7584,17'd7254,17'd7255,17'd7256,17'd7256,17'd7585,17'd7585,17'd6474,17'd6475,17'd6777,17'd6637,17'd7420,17'd7421,17'd7259,17'd7261,17'd7586,17'd7586,17'd7587,17'd7101,17'd7262,17'd7425,17'd7588,17'd7589,17'd7590,17'd7591,17'd7592,17'd7593,17'd7594,17'd7595,17'd7596,17'd7597,17'd7598,17'd7599,17'd7600,17'd7601,17'd7602,17'd7603,17'd7604,17'd7605,17'd7606,17'd7607,17'd7608,17'd7609,17'd7610,17'd7611,17'd7612,17'd7613,17'd7614,17'd7615,17'd7616,17'd7617,17'd7618,17'd7619,17'd7620,17'd7621,17'd7622,17'd7623,17'd7624,17'd7625,17'd7626,17'd7627,17'd7628,17'd7629,17'd7630,17'd7631,17'd7632,17'd7633,17'd7634,17'd7635,17'd7636,17'd7637,17'd7638,17'd7639,17'd7640,17'd7641,17'd7642,17'd7643,17'd7644,17'd7645,17'd7646,17'd7647,17'd7648,17'd6830,17'd889,17'd1197,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd1197,17'd135,17'd7649,17'd7650,17'd7651,17'd3347,17'd7652,17'd4982,17'd7653,17'd7654,17'd7655,17'd6701,17'd7656,17'd7657,17'd7658,17'd7659,17'd7163,17'd7326,17'd7327,17'd7660,17'd7661,17'd7662,17'd6703,17'd7169,17'd6847,17'd6847,17'd6848,17'd6848,17'd7663,17'd7173,17'd7173,17'd7498,17'd7498,17'd7498,17'd7498,17'd7498,17'd7173,17'd7664,17'd7664,17'd7665,17'd7666,17'd7666,17'd7666,17'd7175,17'd7175,17'd7010,17'd7010,17'd6386,17'd6550,17'd6550,17'd6550,17'd6550,17'd6550,17'd6550,17'd6216,17'd7667,17'd7667,17'd6704,17'd6387,17'd6553,17'd6553,17'd6707,17'd6221,17'd6220,17'd7668,17'd7669,17'd6557,17'd6559,17'd7670,17'd7670,17'd6711,17'd6711,17'd7014,17'd7671,17'd7330,17'd7331,17'd7503,17'd7503,17'd7672,17'd7673,17'd7674,17'd7675,17'd6714,17'd7676,17'd7677,17'd7678,17'd7509,17'd7679,17'd7339,17'd3856,17'd6718,17'd7680,17'd3567,17'd6867,17'd633,17'd1681,17'd7681,17'd443,17'd1680,17'd1810,17'd2097,17'd7682,17'd4402,17'd1954,17'd6249,17'd6245,17'd7031,17'd6724,17'd7343,17'd5184,17'd7344,17'd7514,17'd7683,17'd7344,17'd7684,17'd7685,17'd7686,17'd7687,17'd7687,17'd7688,17'd7689,17'd6577,17'd6244,17'd6244,17'd7193,17'd6576,17'd7193,17'd4563,17'd6248,17'd7519,17'd7518,17'd3578,17'd3408,17'd3881,17'd3724,17'd7350,17'd7690,17'd7691,17'd7692,17'd7356,17'd7693,17'd7526,17'd7036,17'd7694,17'd7527,17'd7695,17'd7696,17'd7352,17'd7697,17'd7698,17'd7699,17'd7700,17'd7700,17'd7701,17'd7360,17'd7702,17'd7703,17'd7704,17'd6885,17'd1810,17'd6259,17'd5789,17'd6094,17'd7537,17'd7705,17'd7705,17'd7537,17'd6416,17'd5958,17'd5958,17'd7211,17'd4423,17'd3895,17'd5193,17'd4713,17'd6095,17'd6258,17'd4882,17'd4729,17'd5372,17'd6407,17'd4084,17'd410,17'd642,17'd261,17'd7539,17'd644,17'd1686,17'd1099,17'd1246,17'd601
},
'{
17'd5197,17'd5792,17'd5644,17'd5790,17'd6422,17'd6422,17'd7213,17'd7706,17'd7707,17'd7708,17'd7709,17'd7709,17'd7710,17'd5374,17'd5201,17'd4244,17'd2934,17'd2422,17'd2781,17'd1967,17'd14,17'd466,17'd466,17'd466,17'd4247,17'd1689,17'd6096,17'd6583,17'd7545,17'd5508,17'd7545,17'd7711,17'd3250,17'd3250,17'd1689,17'd2,17'd18,17'd21,17'd24,17'd5,17'd3753,17'd3753,17'd7382,17'd7712,17'd7712,17'd7712,17'd3753,17'd6,17'd5206,17'd1413,17'd7050,17'd7713,17'd6596,17'd6106,17'd7714,17'd7715,17'd7547,17'd7716,17'd7717,17'd7718,17'd7220,17'd7719,17'd7720,17'd7221,17'd7721,17'd7722,17'd7723,17'd7724,17'd7725,17'd7726,17'd7727,17'd5,17'd4,17'd4,17'd4,17'd5,17'd5,17'd5,17'd1690,17'd1690,17'd21,17'd25,17'd1833,17'd1833,17'd7728,17'd7728,17'd7061,17'd7061,17'd7555,17'd7385,17'd7385,17'd7385,17'd7386,17'd7388,17'd6747,17'd6748,17'd7729,17'd7729,17'd7559,17'd7390,17'd7228,17'd7730,17'd7392,17'd7731,17'd7392,17'd6282,17'd6602,17'd7065,17'd7229,17'd7230,17'd7732,17'd7733,17'd7734,17'd7735,17'd7736,17'd7737,17'd7738,17'd7569,17'd7739,17'd5988,17'd6614,17'd7740,17'd7741,17'd7742,17'd7743,17'd7744,17'd7745,17'd7746,17'd7747,17'd6931,17'd6931,17'd7413,17'd7413,17'd7414,17'd7748,17'd7748,17'd7748,17'd7749,17'd7749,17'd7579,17'd7087,17'd7417,17'd7417,17'd6141,17'd7750,17'd7750,17'd5410,17'd5090,17'd4767,17'd7751,17'd7751,17'd3953,17'd3952,17'd3952,17'd6628,17'd4924,17'd5087,17'd5087,17'd6306,17'd6628,17'd7090,17'd6629,17'd6307,17'd7256,17'd7752,17'd7753,17'd7754,17'd7754,17'd6637,17'd7097,17'd7421,17'd7098,17'd7260,17'd7755,17'd7756,17'd7422,17'd7757,17'd7758,17'd7759,17'd7102,17'd7760,17'd7761,17'd7762,17'd7763,17'd7265,17'd7266,17'd7764,17'd7765,17'd7766,17'd7767,17'd7768,17'd7769,17'd7770,17'd7771,17'd7772,17'd7773,17'd7774,17'd7775,17'd7776,17'd7777,17'd7778,17'd7778,17'd7778,17'd7779,17'd7779,17'd7780,17'd7781,17'd7782,17'd7783,17'd7784,17'd7785,17'd7786,17'd7787,17'd7788,17'd7789,17'd7790,17'd7620,17'd7458,17'd7791,17'd7792,17'd7793,17'd7794,17'd7795,17'd7630,17'd7796,17'd7797,17'd7798,17'd7799,17'd7800,17'd7801,17'd7802,17'd7803,17'd7804,17'd7805,17'd7806,17'd7807,17'd7641,17'd7808,17'd7809,17'd7810,17'd7811,17'd7646,17'd7812,17'd7813,17'd889,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd542,17'd133,17'd132,17'd132,17'd131,17'd132,17'd133,17'd542,17'd3025,17'd5593,17'd7814,17'd7815,17'd7816,17'd7817,17'd7818,17'd7819,17'd7820,17'd7490,17'd7821,17'd7822,17'd4679,17'd7658,17'd7659,17'd7823,17'd7824,17'd7327,17'd7166,17'd6844,17'd7825,17'd7167,17'd7169,17'd7826,17'd7170,17'd7827,17'd7827,17'd7172,17'd7828,17'd7829,17'd7830,17'd7831,17'd7832,17'd7833,17'd7834,17'd7828,17'd7835,17'd7835,17'd7173,17'd7664,17'd7173,17'd7175,17'd7666,17'd6385,17'd6385,17'd6385,17'd6386,17'd6849,17'd6849,17'd7329,17'd7329,17'd7329,17'd6550,17'd6550,17'd6550,17'd6550,17'd6215,17'd7667,17'd6704,17'd6704,17'd6387,17'd6707,17'd6707,17'd6221,17'd6391,17'd6391,17'd6555,17'd6557,17'd6559,17'd7836,17'd7837,17'd7838,17'd7839,17'd7839,17'd7840,17'd7330,17'd7841,17'd7016,17'd7016,17'd7842,17'd7843,17'd5766,17'd5018,17'd4381,17'd7019,17'd7844,17'd7678,17'd7845,17'd7846,17'd7847,17'd4861,17'd7848,17'd7849,17'd4864,17'd6084,17'd450,17'd799,17'd7850,17'd2249,17'd1680,17'd6407,17'd7027,17'd7851,17'd7852,17'd2106,17'd4063,17'd4719,17'd4719,17'd5034,17'd7853,17'd7344,17'd7344,17'd7854,17'd7855,17'd7514,17'd7684,17'd7684,17'd7856,17'd7857,17'd7858,17'd7859,17'd7860,17'd7196,17'd7196,17'd7519,17'd7518,17'd4871,17'd6243,17'd7031,17'd7031,17'd6409,17'd7860,17'd7861,17'd3723,17'd7862,17'd7863,17'd7864,17'd7865,17'd7866,17'd7867,17'd7355,17'd7868,17'd7869,17'd7870,17'd7871,17'd7871,17'd7872,17'd7872,17'd7355,17'd7873,17'd7874,17'd6877,17'd7875,17'd7876,17'd7877,17'd7534,17'd7534,17'd7702,17'd7361,17'd4728,17'd4085,17'd4713,17'd6416,17'd6890,17'd6418,17'd6418,17'd7878,17'd6418,17'd6094,17'd6095,17'd4730,17'd5958,17'd4713,17'd3895,17'd3391,17'd4882,17'd5958,17'd4882,17'd4882,17'd4882,17'd3391,17'd445,17'd3742,17'd1243,17'd3899,17'd7879,17'd643,17'd1098,17'd1099,17'd1246,17'd415
},
'{
17'd5197,17'd5645,17'd5644,17'd5790,17'd6422,17'd6423,17'd7880,17'd7708,17'd7881,17'd7881,17'd7882,17'd7883,17'd7047,17'd5197,17'd4087,17'd4428,17'd2784,17'd3250,17'd1967,17'd14,17'd466,17'd466,17'd466,17'd466,17'd1127,17'd1689,17'd6096,17'd7711,17'd7545,17'd5508,17'd7545,17'd7711,17'd3250,17'd1688,17'd1127,17'd2,17'd11,17'd22,17'd5,17'd3753,17'd3753,17'd3753,17'd7712,17'd7712,17'd7712,17'd7884,17'd3753,17'd6,17'd5647,17'd5794,17'd5796,17'd6428,17'd6589,17'd7885,17'd6592,17'd7547,17'd7886,17'd7887,17'd7887,17'd7888,17'd7377,17'd7719,17'd7889,17'd6592,17'd7890,17'd7891,17'd7892,17'd7893,17'd7894,17'd7895,17'd3753,17'd5,17'd4,17'd9,17'd4,17'd4,17'd5,17'd5,17'd1690,17'd1690,17'd21,17'd25,17'd1833,17'd1833,17'd7728,17'd7728,17'd7061,17'd7061,17'd7555,17'd7555,17'd7385,17'd7385,17'd7388,17'd7557,17'd6747,17'd6905,17'd7896,17'd7896,17'd7559,17'd7063,17'd7228,17'd7730,17'd7730,17'd7392,17'd7392,17'd6602,17'd6602,17'd7393,17'd7897,17'd7231,17'd6909,17'd7898,17'd7899,17'd7900,17'd7901,17'd7902,17'd7903,17'd7904,17'd7905,17'd6762,17'd7906,17'd7907,17'd7908,17'd7573,17'd7909,17'd7910,17'd7911,17'd7749,17'd7413,17'd6770,17'd7413,17'd7413,17'd7414,17'd7414,17'd7748,17'd7748,17'd7748,17'd7748,17'd7579,17'd7087,17'd7417,17'd6141,17'd6141,17'd5837,17'd5255,17'd4927,17'd4767,17'd4611,17'd7912,17'd7751,17'd3953,17'd3952,17'd4291,17'd4291,17'd4924,17'd5250,17'd5087,17'd5087,17'd6306,17'd6628,17'd7090,17'd6629,17'd7093,17'd7913,17'd7754,17'd7754,17'd7914,17'd7915,17'd7097,17'd7421,17'd7755,17'd7916,17'd7755,17'd7756,17'd7756,17'd7756,17'd7917,17'd7918,17'd7919,17'd7920,17'd7921,17'd7763,17'd7922,17'd7923,17'd7924,17'd7925,17'd7926,17'd7927,17'd7928,17'd7929,17'd7930,17'd7931,17'd7932,17'd7933,17'd7934,17'd7935,17'd7936,17'd7937,17'd7938,17'd7939,17'd7940,17'd7941,17'd7941,17'd7942,17'd7943,17'd7944,17'd7945,17'd7946,17'd7947,17'd7948,17'd7949,17'd7950,17'd7951,17'd7952,17'd7953,17'd7954,17'd7955,17'd7620,17'd7621,17'd7956,17'd7957,17'd7958,17'd7959,17'd7960,17'd7961,17'd7962,17'd7963,17'd7964,17'd7965,17'd7966,17'd7967,17'd7968,17'd7969,17'd7970,17'd7971,17'd7972,17'd7973,17'd7974,17'd7975,17'd7976,17'd7977,17'd7978,17'd7812,17'd7979,17'd7980,17'd1045,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd132,17'd131,17'd131,17'd132,17'd542,17'd542,17'd133,17'd132,17'd131,17'd131,17'd132,17'd133,17'd542,17'd132,17'd7981,17'd7982,17'd7983,17'd7984,17'd7985,17'd7986,17'd7987,17'd6539,17'd7988,17'd4989,17'd4678,17'd7658,17'd7325,17'd7326,17'd7824,17'd7989,17'd7494,17'd7990,17'd7825,17'd7991,17'd7168,17'd7169,17'd7169,17'd7992,17'd7827,17'd7993,17'd7828,17'd7994,17'd7995,17'd7996,17'd7997,17'd7998,17'd7832,17'd7832,17'd7834,17'd7828,17'd7498,17'd7828,17'd7173,17'd7173,17'd7174,17'd7175,17'd7010,17'd6386,17'd6386,17'd6386,17'd6849,17'd6849,17'd6849,17'd7329,17'd7329,17'd7329,17'd6550,17'd6550,17'd6550,17'd6550,17'd7667,17'd7667,17'd6704,17'd6704,17'd7999,17'd8000,17'd6707,17'd5919,17'd6220,17'd6220,17'd7500,17'd6557,17'd8001,17'd8002,17'd7501,17'd6711,17'd7838,17'd7839,17'd6712,17'd7331,17'd8003,17'd8003,17'd8003,17'd7842,17'd7184,17'd8004,17'd8005,17'd8006,17'd7019,17'd7677,17'd8007,17'd8008,17'd7846,17'd8009,17'd8010,17'd8011,17'd8012,17'd4708,17'd6720,17'd8013,17'd8014,17'd8015,17'd624,17'd2392,17'd6888,17'd5358,17'd1392,17'd8016,17'd2247,17'd4063,17'd4405,17'd4562,17'd8017,17'd7853,17'd7684,17'd8018,17'd7855,17'd7854,17'd7344,17'd7344,17'd8018,17'd8019,17'd8020,17'd8021,17'd8022,17'd8023,17'd7196,17'd7196,17'd4234,17'd4567,17'd4718,17'd4407,17'd6243,17'd6577,17'd7860,17'd7861,17'd3725,17'd8024,17'd8025,17'd7864,17'd8026,17'd7865,17'd8027,17'd8028,17'd8029,17'd8030,17'd7872,17'd7871,17'd7871,17'd8031,17'd7870,17'd7871,17'd8032,17'd7873,17'd8033,17'd8033,17'd8034,17'd7532,17'd8035,17'd7534,17'd8036,17'd7702,17'd3712,17'd6415,17'd4713,17'd5958,17'd6890,17'd6094,17'd7364,17'd7878,17'd6418,17'd6418,17'd6258,17'd6258,17'd6581,17'd4713,17'd3391,17'd4085,17'd4882,17'd5958,17'd5958,17'd4882,17'd4882,17'd3744,17'd3895,17'd1810,17'd1396,17'd3899,17'd7879,17'd606,17'd952,17'd193,17'd421,17'd415
},
'{
17'd5790,17'd5790,17'd5790,17'd5644,17'd5510,17'd7046,17'd7706,17'd8037,17'd8038,17'd8038,17'd8039,17'd7046,17'd5374,17'd5201,17'd3903,17'd4733,17'd3250,17'd1689,17'd14,17'd14,17'd466,17'd2595,17'd466,17'd466,17'd1127,17'd1689,17'd7711,17'd7545,17'd4887,17'd4246,17'd4887,17'd7545,17'd3250,17'd1688,17'd1127,17'd12,17'd21,17'd23,17'd6,17'd3753,17'd5793,17'd8040,17'd5205,17'd5205,17'd5205,17'd5205,17'd7,17'd7,17'd8041,17'd6588,17'd6099,17'd8042,17'd6733,17'd7722,17'd6738,17'd8043,17'd7718,17'd7716,17'd7888,17'd7219,17'd7548,17'd7550,17'd6896,17'd6737,17'd8044,17'd8045,17'd6435,17'd7050,17'd8046,17'd7894,17'd5,17'd5206,17'd5647,17'd1413,17'd8,17'd5,17'd7383,17'd7383,17'd1690,17'd2937,17'd25,17'd25,17'd467,17'd467,17'd7555,17'd7555,17'd7555,17'd7555,17'd7555,17'd7555,17'd7555,17'd8047,17'd7557,17'd8048,17'd7063,17'd7063,17'd7559,17'd7390,17'd6907,17'd7228,17'd6602,17'd6113,17'd6602,17'd6602,17'd8049,17'd6602,17'd7065,17'd8050,17'd8051,17'd8052,17'd7070,17'd8053,17'd8054,17'd7234,17'd8055,17'd8056,17'd8057,17'd6761,17'd6919,17'd8058,17'd8059,17'd8060,17'd8061,17'd8062,17'd7080,17'd8063,17'd7911,17'd8064,17'd7580,17'd7413,17'd7413,17'd7413,17'd7414,17'd7414,17'd7748,17'd8065,17'd7748,17'd7748,17'd7579,17'd7087,17'd7417,17'd6468,17'd6468,17'd5409,17'd5255,17'd4611,17'd8066,17'd8067,17'd7751,17'd8068,17'd7751,17'd4464,17'd4127,17'd4127,17'd5250,17'd5250,17'd5251,17'd5087,17'd5087,17'd4924,17'd7253,17'd7090,17'd7584,17'd7584,17'd8069,17'd7915,17'd7097,17'd7099,17'd8070,17'd7755,17'd8071,17'd8072,17'd8073,17'd8074,17'd7917,17'd8075,17'd8076,17'd8076,17'd7760,17'd8077,17'd7763,17'd8078,17'd7105,17'd8079,17'd7105,17'd8080,17'd8081,17'd8082,17'd8083,17'd8084,17'd8085,17'd8086,17'd8087,17'd8088,17'd8089,17'd8090,17'd8091,17'd8092,17'd8093,17'd8094,17'd8095,17'd8094,17'd8096,17'd8097,17'd8097,17'd8098,17'd8099,17'd8100,17'd8101,17'd8102,17'd8103,17'd7948,17'd8104,17'd7950,17'd8105,17'd7953,17'd8106,17'd7955,17'd8107,17'd8108,17'd8109,17'd8110,17'd8111,17'd8112,17'd8113,17'd8114,17'd8115,17'd8116,17'd7964,17'd8117,17'd8118,17'd8119,17'd8120,17'd8121,17'd8122,17'd8123,17'd8124,17'd8125,17'd8126,17'd8127,17'd8128,17'd8129,17'd8130,17'd8131,17'd8132,17'd889,17'd1197,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd131,17'd132,17'd133,17'd542,17'd133,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd131,17'd6532,17'd8133,17'd8134,17'd8135,17'd8136,17'd8137,17'd8138,17'd8139,17'd8140,17'd8141,17'd8142,17'd8143,17'd7163,17'd7164,17'd8144,17'd7494,17'd7661,17'd8145,17'd8145,17'd7992,17'd7827,17'd8146,17'd8147,17'd7992,17'd7827,17'd7173,17'd8148,17'd8149,17'd8150,17'd8151,17'd8152,17'd8153,17'd7995,17'd7995,17'd7994,17'd7832,17'd7830,17'd7830,17'd7829,17'd7174,17'd7174,17'd7174,17'd7174,17'd7175,17'd7010,17'd7010,17'd7010,17'd6849,17'd6849,17'd6849,17'd7329,17'd7329,17'd7329,17'd6849,17'd6550,17'd6550,17'd7667,17'd7667,17'd7667,17'd7176,17'd6704,17'd6704,17'd6553,17'd6553,17'd8154,17'd6220,17'd7668,17'd7500,17'd6557,17'd8155,17'd6559,17'd7501,17'd7501,17'd7838,17'd8156,17'd8157,17'd6562,17'd8003,17'd8003,17'd7016,17'd8158,17'd8159,17'd8160,17'd8005,17'd8161,17'd7019,17'd6400,17'd7678,17'd7679,17'd4545,17'd4045,17'd5022,17'd8162,17'd8163,17'd5025,17'd8164,17'd1943,17'd1120,17'd2249,17'd1667,17'd2577,17'd8165,17'd2762,17'd1392,17'd8166,17'd2759,17'd5033,17'd4718,17'd8167,17'd8168,17'd7685,17'd8169,17'd8170,17'd8170,17'd7854,17'd7514,17'd8018,17'd8171,17'd8172,17'd8173,17'd8174,17'd8022,17'd8023,17'd8175,17'd3578,17'd7518,17'd6576,17'd7193,17'd6577,17'd6577,17'd7860,17'd7195,17'd8176,17'd8177,17'd7350,17'd8178,17'd7691,17'd8026,17'd8179,17'd8027,17'd8028,17'd7697,17'd7872,17'd8031,17'd8180,17'd8180,17'd7871,17'd7871,17'd7697,17'd7873,17'd8181,17'd7874,17'd7875,17'd7876,17'd8182,17'd8035,17'd8183,17'd8183,17'd8184,17'd2097,17'd8185,17'd5630,17'd8186,17'd8187,17'd7364,17'd7364,17'd7364,17'd7364,17'd6418,17'd6094,17'd6581,17'd4882,17'd4085,17'd4085,17'd4882,17'd5958,17'd5958,17'd5958,17'd5958,17'd4085,17'd445,17'd2559,17'd410,17'd426,17'd8188,17'd643,17'd1098,17'd1099,17'd1246,17'd415
},
'{
17'd5790,17'd5643,17'd5790,17'd7541,17'd6586,17'd7883,17'd8037,17'd8037,17'd8189,17'd7882,17'd7883,17'd5375,17'd5645,17'd4427,17'd4088,17'd4887,17'd2781,17'd1967,17'd14,17'd14,17'd466,17'd466,17'd466,17'd1127,17'd1689,17'd3250,17'd7545,17'd7545,17'd4246,17'd4887,17'd4887,17'd7545,17'd1688,17'd1127,17'd2,17'd3,17'd25,17'd5,17'd5205,17'd5205,17'd8040,17'd8040,17'd8190,17'd5205,17'd5205,17'd6,17'd7,17'd5206,17'd6098,17'd6266,17'd8042,17'd6272,17'd7722,17'd7218,17'd8191,17'd7888,17'd7887,17'd7378,17'd7220,17'd7719,17'd8192,17'd6895,17'd6895,17'd7889,17'd8193,17'd8194,17'd5963,17'd6588,17'd8195,17'd8196,17'd5206,17'd5514,17'd5512,17'd5647,17'd8,17'd5,17'd7383,17'd1690,17'd2937,17'd2937,17'd25,17'd25,17'd467,17'd285,17'd7385,17'd7555,17'd7555,17'd7555,17'd7555,17'd7555,17'd8047,17'd8197,17'd8048,17'd8198,17'd7390,17'd7390,17'd7390,17'd7560,17'd7228,17'd7228,17'd6602,17'd6602,17'd6602,17'd6750,17'd8199,17'd8200,17'd8201,17'd8051,17'd8052,17'd8202,17'd8203,17'd8204,17'd8205,17'd8206,17'd8207,17'd6917,17'd7400,17'd6613,17'd8208,17'd8209,17'd8060,17'd8210,17'd8211,17'd8212,17'd8213,17'd8214,17'd8215,17'd8216,17'd8217,17'd7580,17'd7413,17'd7413,17'd7414,17'd7414,17'd8065,17'd8065,17'd7748,17'd8218,17'd7087,17'd6142,17'd6468,17'd5409,17'd5409,17'd5410,17'd4767,17'd8066,17'd8067,17'd8067,17'd7751,17'd7751,17'd7912,17'd4766,17'd4610,17'd4610,17'd5250,17'd5250,17'd5251,17'd5087,17'd5087,17'd5085,17'd4923,17'd7090,17'd7095,17'd7258,17'd7097,17'd7099,17'd7260,17'd7423,17'd8219,17'd8219,17'd8071,17'd8220,17'd8074,17'd8220,17'd8075,17'd8221,17'd8221,17'd8222,17'd8223,17'd7762,17'd7923,17'd8224,17'd8080,17'd8225,17'd8225,17'd8226,17'd8227,17'd8228,17'd8229,17'd8230,17'd8231,17'd8232,17'd8233,17'd8234,17'd8235,17'd8236,17'd8237,17'd8238,17'd8239,17'd8240,17'd8241,17'd8242,17'd8243,17'd8244,17'd8245,17'd8246,17'd8247,17'd8247,17'd8248,17'd8249,17'd8249,17'd8250,17'd8251,17'd8252,17'd7948,17'd8253,17'd8254,17'd8255,17'd8256,17'd7954,17'd8257,17'd8258,17'd8259,17'd8260,17'd8261,17'd8262,17'd8263,17'd8264,17'd8265,17'd8266,17'd8267,17'd8268,17'd8269,17'd8270,17'd8271,17'd8272,17'd8273,17'd8274,17'd8275,17'd8276,17'd8277,17'd8278,17'd8279,17'd7812,17'd8131,17'd889,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd3811,17'd7650,17'd8280,17'd8281,17'd8282,17'd8283,17'd8284,17'd8285,17'd8286,17'd8287,17'd8288,17'd8289,17'd6544,17'd7164,17'd7165,17'd6383,17'd7328,17'd8145,17'd8290,17'd8291,17'd8291,17'd8291,17'd8292,17'd8292,17'd7663,17'd7173,17'd7828,17'd8293,17'd8294,17'd8295,17'd8296,17'd8297,17'd8298,17'd8298,17'd8299,17'd8152,17'd7997,17'd8300,17'd8300,17'd7830,17'd7829,17'd7174,17'd7174,17'd7174,17'd7174,17'd8301,17'd7010,17'd7010,17'd7010,17'd6849,17'd6849,17'd6849,17'd7329,17'd7329,17'd7329,17'd6550,17'd6550,17'd8302,17'd7667,17'd7667,17'd7667,17'd6704,17'd6704,17'd7999,17'd6553,17'd8303,17'd8154,17'd8304,17'd7668,17'd7500,17'd6557,17'd6557,17'd6709,17'd6559,17'd7501,17'd6394,17'd8305,17'd8305,17'd8306,17'd8306,17'd7330,17'd7672,17'd8307,17'd8308,17'd8309,17'd4542,17'd8310,17'd7186,17'd8311,17'd6401,17'd7189,17'd6570,17'd5930,17'd5931,17'd8312,17'd4393,17'd8313,17'd6405,17'd8314,17'd794,17'd1380,17'd8315,17'd8316,17'd1393,17'd8317,17'd4230,17'd2402,17'd5949,17'd4718,17'd4871,17'd8318,17'd7346,17'd8169,17'd8018,17'd8170,17'd7855,17'd7854,17'd8018,17'd8171,17'd8172,17'd8319,17'd8320,17'd8174,17'd8022,17'd8321,17'd7861,17'd7861,17'd7689,17'd6576,17'd6577,17'd6577,17'd7196,17'd7860,17'd8322,17'd8323,17'd4072,17'd7690,17'd8324,17'd7691,17'd8325,17'd8179,17'd8326,17'd8327,17'd8031,17'd8031,17'd8180,17'd8328,17'd8329,17'd8180,17'd7355,17'd7697,17'd7698,17'd7698,17'd8330,17'd8330,17'd5950,17'd8182,17'd8331,17'd8332,17'd8333,17'd8334,17'd5630,17'd8185,17'd7365,17'd8187,17'd7364,17'd7364,17'd7364,17'd7364,17'd7364,17'd6418,17'd6416,17'd5958,17'd4713,17'd4085,17'd4713,17'd5958,17'd6581,17'd6581,17'd5958,17'd4713,17'd3895,17'd2392,17'd1823,17'd260,17'd3746,17'd606,17'd1272,17'd193,17'd421,17'd415
},
'{
17'd5510,17'd6422,17'd5510,17'd6585,17'd6423,17'd7709,17'd8335,17'd8336,17'd7882,17'd7883,17'd8337,17'd5959,17'd5201,17'd3903,17'd2593,17'd2422,17'd1689,17'd14,17'd2,17'd466,17'd466,17'd466,17'd1127,17'd14,17'd1689,17'd3250,17'd7545,17'd4246,17'd4887,17'd4887,17'd4887,17'd7545,17'd1127,17'd2,17'd12,17'd1275,17'd4,17'd6,17'd5205,17'd8040,17'd8338,17'd8339,17'd8340,17'd5205,17'd3753,17'd6,17'd7,17'd5514,17'd6588,17'd6435,17'd8341,17'd8342,17'd8343,17'd8191,17'd8344,17'd7887,17'd7718,17'd7886,17'd7550,17'd8345,17'd8343,17'd7221,17'd8192,17'd8346,17'd6271,17'd6102,17'd5962,17'd8347,17'd6098,17'd6097,17'd7375,17'd7375,17'd5513,17'd5378,17'd6,17'd5,17'd1690,17'd1690,17'd2937,17'd4429,17'd25,17'd25,17'd285,17'd285,17'd7385,17'd7555,17'd7555,17'd8047,17'd8047,17'd8047,17'd8197,17'd8197,17'd8198,17'd8198,17'd7390,17'd7390,17'd7227,17'd7391,17'd7392,17'd7228,17'd6602,17'd6750,17'd8348,17'd8348,17'd8349,17'd8350,17'd8351,17'd8352,17'd8353,17'd8354,17'd8355,17'd8356,17'd7901,17'd8357,17'd8358,17'd8057,17'd6290,17'd8359,17'd8360,17'd8361,17'd8362,17'd8363,17'd8364,17'd8063,17'd8365,17'd8217,17'd8217,17'd8217,17'd7749,17'd7749,17'd8366,17'd8366,17'd8367,17'd8367,17'd7748,17'd7748,17'd8218,17'd8218,17'd8368,17'd8369,17'd8370,17'd7750,17'd4927,17'd4611,17'd8066,17'd8371,17'd8372,17'd8371,17'd8066,17'd8066,17'd7088,17'd4926,17'd6627,17'd6627,17'd5087,17'd5251,17'd8373,17'd8373,17'd8373,17'd8374,17'd5085,17'd5085,17'd8375,17'd8376,17'd8070,17'd7756,17'd8377,17'd8378,17'd8379,17'd8379,17'd8380,17'd8381,17'd8382,17'd8383,17'd8384,17'd8222,17'd8385,17'd8077,17'd8386,17'd8387,17'd7924,17'd8388,17'd8389,17'd7432,17'd8390,17'd8391,17'd8392,17'd8393,17'd8394,17'd8395,17'd8396,17'd8397,17'd8398,17'd8399,17'd8400,17'd8401,17'd8402,17'd8403,17'd8404,17'd8405,17'd8406,17'd8407,17'd8407,17'd8408,17'd8409,17'd8410,17'd8411,17'd8412,17'd8413,17'd8414,17'd8414,17'd8415,17'd8416,17'd8417,17'd8418,17'd8249,17'd8419,17'd8252,17'd8420,17'd7949,17'd8421,17'd8422,17'd8423,17'd8424,17'd8425,17'd8426,17'd8427,17'd8428,17'd8429,17'd8430,17'd8431,17'd8432,17'd8433,17'd8434,17'd8435,17'd8436,17'd8437,17'd8438,17'd8439,17'd8440,17'd8441,17'd8442,17'd8443,17'd7646,17'd8444,17'd6830,17'd719,17'd542,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd542,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd542,17'd133,17'd357,17'd8445,17'd8446,17'd8447,17'd8448,17'd8136,17'd8449,17'd8450,17'd8451,17'd6836,17'd6700,17'd6542,17'd6543,17'd7163,17'd7165,17'd7166,17'd5914,17'd6384,17'd7662,17'd8452,17'd8453,17'd8454,17'd8454,17'd8455,17'd7172,17'd7498,17'd7828,17'd7834,17'd8456,17'd8457,17'd8458,17'd8295,17'd8459,17'd8460,17'd8461,17'd8461,17'd8462,17'd8463,17'd8464,17'd8465,17'd8466,17'd8467,17'd8468,17'd8469,17'd8470,17'd8470,17'd8470,17'd7174,17'd7175,17'd7175,17'd7175,17'd6848,17'd6848,17'd6848,17'd8146,17'd8146,17'd7329,17'd7168,17'd7168,17'd7168,17'd7667,17'd7667,17'd7667,17'd7667,17'd7176,17'd6704,17'd7999,17'd6707,17'd8154,17'd6220,17'd7668,17'd7500,17'd7669,17'd8471,17'd6557,17'd6559,17'd8472,17'd8473,17'd8473,17'd8474,17'd8306,17'd7331,17'd7331,17'd8475,17'd7017,17'd8159,17'd8476,17'd6228,17'd8477,17'd6714,17'd8478,17'd7188,17'd6233,17'd8479,17'd4044,17'd3860,17'd8480,17'd8481,17'd8482,17'd2557,17'd1122,17'd8483,17'd8484,17'd8485,17'd8486,17'd2921,17'd4061,17'd8487,17'd8488,17'd8489,17'd4871,17'd7688,17'd7688,17'd8490,17'd7856,17'd8171,17'd8491,17'd8170,17'd8170,17'd7856,17'd8172,17'd8492,17'd8493,17'd8494,17'd8495,17'd8496,17'd8176,17'd7861,17'd7688,17'd7030,17'd8497,17'd6577,17'd7519,17'd7860,17'd8322,17'd8496,17'd8323,17'd8177,17'd7690,17'd7864,17'd8026,17'd8498,17'd8499,17'd8500,17'd8501,17'd8180,17'd8180,17'd8328,17'd8501,17'd8328,17'd8329,17'd8329,17'd8032,17'd8028,17'd8502,17'd8330,17'd8503,17'd8503,17'd8504,17'd8035,17'd8505,17'd7703,17'd2097,17'd8185,17'd7365,17'd8187,17'd7705,17'd7537,17'd8506,17'd8506,17'd7537,17'd8507,17'd6416,17'd5958,17'd4882,17'd4729,17'd4713,17'd5958,17'd6581,17'd6581,17'd5958,17'd4423,17'd2392,17'd2559,17'd190,17'd259,17'd3746,17'd643,17'd1685,17'd603,17'd1246,17'd415
},
'{
17'd5510,17'd6585,17'd6586,17'd6729,17'd7883,17'd8508,17'd8336,17'd7882,17'd8039,17'd8509,17'd6261,17'd5201,17'd4244,17'd4245,17'd2422,17'd1688,17'd1127,17'd1127,17'd466,17'd466,17'd466,17'd466,17'd1127,17'd1967,17'd3250,17'd2422,17'd4887,17'd4246,17'd4887,17'd4887,17'd4577,17'd7711,17'd14,17'd12,17'd806,17'd2591,17'd8,17'd7,17'd5205,17'd8040,17'd8339,17'd8339,17'd8340,17'd5205,17'd6,17'd5206,17'd8510,17'd6098,17'd6099,17'd8511,17'd6899,17'd6897,17'd7378,17'd8512,17'd8513,17'd8514,17'd8515,17'd7219,17'd8516,17'd8517,17'd6738,17'd8517,17'd8345,17'd7054,17'd6103,17'd8518,17'd6732,17'd6266,17'd6731,17'd6588,17'd8519,17'd8520,17'd5648,17'd5514,17'd8,17'd23,17'd1691,17'd467,17'd1833,17'd1833,17'd808,17'd25,17'd285,17'd285,17'd7555,17'd7555,17'd7555,17'd8047,17'd8047,17'd8047,17'd8197,17'd8521,17'd8198,17'd8198,17'd7390,17'd7390,17'd7227,17'd7391,17'd7392,17'd7228,17'd8199,17'd8199,17'd8522,17'd8523,17'd8524,17'd8525,17'd6909,17'd7070,17'd8526,17'd8527,17'd8356,17'd8528,17'd8529,17'd8530,17'd8531,17'd6918,17'd7238,17'd8360,17'd8532,17'd8533,17'd8534,17'd8364,17'd8063,17'd7911,17'd8217,17'd7580,17'd7580,17'd7580,17'd7749,17'd7414,17'd8366,17'd8366,17'd8367,17'd8367,17'd7748,17'd8218,17'd8535,17'd8536,17'd8369,17'd8537,17'd7750,17'd8538,17'd4611,17'd8066,17'd8371,17'd8372,17'd8372,17'd8539,17'd4611,17'd4767,17'd4926,17'd4925,17'd6627,17'd6627,17'd5251,17'd5251,17'd8373,17'd8373,17'd8540,17'd8540,17'd8373,17'd8541,17'd8376,17'd7422,17'd7756,17'd7917,17'd8378,17'd8542,17'd8542,17'd8381,17'd8543,17'd8544,17'd8545,17'd8546,17'd8545,17'd8547,17'd8077,17'd7264,17'd8387,17'd8548,17'd7924,17'd8549,17'd7432,17'd8550,17'd8551,17'd8552,17'd8553,17'd8554,17'd8555,17'd8556,17'd8557,17'd8558,17'd8559,17'd8560,17'd8561,17'd8562,17'd8563,17'd8564,17'd8565,17'd8566,17'd8567,17'd8567,17'd8568,17'd8568,17'd8569,17'd8569,17'd8570,17'd8570,17'd8571,17'd8572,17'd8413,17'd8413,17'd8413,17'd8573,17'd8574,17'd8574,17'd8575,17'd8576,17'd8577,17'd8578,17'd8579,17'd8580,17'd8581,17'd7949,17'd8582,17'd8583,17'd8584,17'd8585,17'd8586,17'd8587,17'd8588,17'd8589,17'd8590,17'd8268,17'd8591,17'd8592,17'd7639,17'd8593,17'd8274,17'd8594,17'd8595,17'd8596,17'd7481,17'd7811,17'd8597,17'd8444,17'd6529,17'd719,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd132,17'd133,17'd542,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd542,17'd132,17'd5593,17'd8598,17'd8599,17'd8600,17'd8601,17'd8602,17'd8603,17'd6540,17'd8604,17'd8605,17'd8606,17'd8607,17'd7658,17'd8608,17'd7327,17'd7328,17'd6846,17'd6846,17'd8290,17'd8452,17'd8453,17'd8609,17'd8610,17'd8611,17'd8612,17'd8613,17'd7833,17'd8614,17'd8615,17'd8616,17'd8617,17'd8618,17'd8619,17'd8460,17'd8620,17'd8621,17'd8622,17'd8623,17'd8624,17'd8625,17'd8626,17'd8627,17'd8467,17'd8468,17'd8470,17'd8470,17'd8470,17'd8470,17'd7174,17'd7175,17'd7175,17'd7175,17'd6848,17'd6848,17'd6848,17'd6848,17'd7329,17'd7329,17'd7168,17'd7168,17'd8628,17'd7667,17'd7667,17'd7667,17'd7176,17'd7176,17'd7999,17'd7999,17'd8629,17'd8154,17'd8304,17'd7499,17'd7668,17'd7500,17'd7669,17'd6557,17'd6558,17'd8472,17'd8630,17'd8631,17'd8632,17'd8633,17'd8633,17'd8634,17'd8475,17'd7017,17'd8635,17'd5766,17'd8636,17'd8310,17'd8637,17'd4211,17'd4701,17'd5927,17'd5927,17'd4044,17'd8638,17'd4863,17'd8481,17'd3389,17'd451,17'd8639,17'd8640,17'd8641,17'd8642,17'd8643,17'd7536,17'd8644,17'd8645,17'd6088,17'd7518,17'd7688,17'd7688,17'd8490,17'd8169,17'd7856,17'd8491,17'd8491,17'd8491,17'd8170,17'd8019,17'd7857,17'd8493,17'd8493,17'd8646,17'd8495,17'd8323,17'd8176,17'd7348,17'd6873,17'd7030,17'd8497,17'd7519,17'd7519,17'd4567,17'd8322,17'd8647,17'd8648,17'd8649,17'd8650,17'd8026,17'd8651,17'd7865,17'd8652,17'd8653,17'd8501,17'd8180,17'd8329,17'd8654,17'd8654,17'd8328,17'd8329,17'd7697,17'd8327,17'd8502,17'd7351,17'd8330,17'd8655,17'd8656,17'd8657,17'd8658,17'd8659,17'd8660,17'd5940,17'd7365,17'd8187,17'd7705,17'd7537,17'd8506,17'd8506,17'd7537,17'd7537,17'd6416,17'd6416,17'd5958,17'd4713,17'd4729,17'd5958,17'd6581,17'd5958,17'd5958,17'd4882,17'd4085,17'd1810,17'd4084,17'd970,17'd2779,17'd206,17'd971,17'd603,17'd1246,17'd1529
},
'{
17'd6585,17'd6585,17'd6586,17'd7883,17'd8508,17'd8336,17'd7882,17'd7882,17'd7883,17'd5375,17'd5645,17'd4427,17'd3751,17'd2935,17'd1688,17'd1127,17'd14,17'd2,17'd2,17'd2,17'd466,17'd466,17'd1127,17'd1689,17'd7545,17'd7545,17'd2784,17'd2784,17'd2784,17'd2784,17'd3250,17'd1689,17'd2,17'd806,17'd10,17'd9,17'd5206,17'd5205,17'd8040,17'd8040,17'd8339,17'd8339,17'd8340,17'd5205,17'd8,17'd5512,17'd7893,17'd8661,17'd6105,17'd6899,17'd6898,17'd7221,17'd8515,17'd8514,17'd8662,17'd8663,17'd8664,17'd8665,17'd7720,17'd8343,17'd8666,17'd8667,17'd8668,17'd6431,17'd8669,17'd8670,17'd7223,17'd6428,17'd6435,17'd6732,17'd8671,17'd5961,17'd5649,17'd5514,17'd5970,17'd1691,17'd1832,17'd467,17'd1833,17'd286,17'd10,17'd10,17'd467,17'd467,17'd7555,17'd7555,17'd7388,17'd7388,17'd8197,17'd8197,17'd8048,17'd8048,17'd7063,17'd7063,17'd7063,17'd7063,17'd7228,17'd7228,17'd6602,17'd6602,17'd8348,17'd8348,17'd8523,17'd8672,17'd8673,17'd6908,17'd6910,17'd8674,17'd7899,17'd8675,17'd8676,17'd8677,17'd8530,17'd8678,17'd7237,17'd8679,17'd8680,17'd8681,17'd8533,17'd8363,17'd8364,17'd8682,17'd8683,17'd8216,17'd8216,17'd8684,17'd8685,17'd8685,17'd7748,17'd8367,17'd8686,17'd8686,17'd8367,17'd8367,17'd8218,17'd8218,17'd8535,17'd8687,17'd8369,17'd8537,17'd7750,17'd8538,17'd8066,17'd8371,17'd7751,17'd7751,17'd8371,17'd8688,17'd4767,17'd4767,17'd5254,17'd5253,17'd5254,17'd5252,17'd8689,17'd8689,17'd8690,17'd8373,17'd8691,17'd8691,17'd8692,17'd8693,17'd8074,17'd8220,17'd8379,17'd8382,17'd8382,17'd8694,17'd8694,17'd8695,17'd8696,17'd8697,17'd8698,17'd8699,17'd8700,17'd8701,17'd8702,17'd8702,17'd8703,17'd7427,17'd8078,17'd8079,17'd8704,17'd8705,17'd8706,17'd8707,17'd8708,17'd8709,17'd8710,17'd8711,17'd8712,17'd8713,17'd8714,17'd8715,17'd8716,17'd8717,17'd8718,17'd8719,17'd8720,17'd8720,17'd8721,17'd8721,17'd8722,17'd8722,17'd8723,17'd8723,17'd8569,17'd8724,17'd8725,17'd8725,17'd8726,17'd8410,17'd8409,17'd8727,17'd8568,17'd8728,17'd8569,17'd8724,17'd8569,17'd8729,17'd8729,17'd8730,17'd8731,17'd8575,17'd8732,17'd8733,17'd8734,17'd8735,17'd8736,17'd8737,17'd8738,17'd8739,17'd8740,17'd8741,17'd8742,17'd8743,17'd8744,17'd8745,17'd8746,17'd8747,17'd8748,17'd8749,17'd8128,17'd8750,17'd8751,17'd7647,17'd6529,17'd6830,17'd542,17'd542,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd542,17'd542,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd542,17'd131,17'd8752,17'd8753,17'd3346,17'd8754,17'd8755,17'd6538,17'd8756,17'd8757,17'd8606,17'd8758,17'd6380,17'd8289,17'd6544,17'd7164,17'd7327,17'd7990,17'd7167,17'd7167,17'd8290,17'd8452,17'd8453,17'd8759,17'd8760,17'd8761,17'd8762,17'd8763,17'd8764,17'd8765,17'd8766,17'd8767,17'd8768,17'd8769,17'd8770,17'd8460,17'd8771,17'd8622,17'd8772,17'd8773,17'd8774,17'd8775,17'd8776,17'd8777,17'd8778,17'd8466,17'd7830,17'd7829,17'd8470,17'd8470,17'd7174,17'd7174,17'd7174,17'd7174,17'd7663,17'd7663,17'd7663,17'd7663,17'd8146,17'd8146,17'd7329,17'd7168,17'd7168,17'd6550,17'd8302,17'd8302,17'd7667,17'd7667,17'd8779,17'd7999,17'd7999,17'd6707,17'd8154,17'd6220,17'd7499,17'd7668,17'd8780,17'd7669,17'd7669,17'd6557,17'd7011,17'd8472,17'd8781,17'd8632,17'd8632,17'd8157,17'd8782,17'd8783,17'd7843,17'd8784,17'd8476,17'd8785,17'd8161,17'd6074,17'd4700,17'd4212,17'd4212,17'd5769,17'd3857,17'd8638,17'd8786,17'd8787,17'd8788,17'd442,17'd8789,17'd8790,17'd3733,17'd6093,17'd7361,17'd8791,17'd8792,17'd2756,17'd8793,17'd7195,17'd7347,17'd7348,17'd8490,17'd8794,17'd8170,17'd8795,17'd8491,17'd8491,17'd8796,17'd8797,17'd8493,17'd8798,17'd8799,17'd8800,17'd8801,17'd8802,17'd8022,17'd7347,17'd7347,17'd7348,17'd7518,17'd7519,17'd7518,17'd7518,17'd8803,17'd8804,17'd8648,17'd8805,17'd8806,17'd8807,17'd8808,17'd7866,17'd8027,17'd8809,17'd8328,17'd8329,17'd8501,17'd8654,17'd8501,17'd8328,17'd8032,17'd7873,17'd7698,17'd7698,17'd8330,17'd7034,17'd8810,17'd8811,17'd8792,17'd8505,17'd8791,17'd3712,17'd5940,17'd4714,17'd7537,17'd7537,17'd7538,17'd7538,17'd7537,17'd7537,17'd6416,17'd6416,17'd6416,17'd4869,17'd4729,17'd5958,17'd6581,17'd5958,17'd5958,17'd4728,17'd1810,17'd3742,17'd8812,17'd970,17'd206,17'd206,17'd971,17'd603,17'd1246,17'd2763
},
'{
17'd6585,17'd8813,17'd6893,17'd7709,17'd8335,17'd8336,17'd7882,17'd7883,17'd7046,17'd5198,17'd5201,17'd3903,17'd2593,17'd3250,17'd1127,17'd2,17'd2,17'd2,17'd2,17'd2,17'd2,17'd1127,17'd1688,17'd1688,17'd5508,17'd7545,17'd2784,17'd2784,17'd2784,17'd2422,17'd3250,17'd1127,17'd12,17'd8814,17'd25,17'd8,17'd7,17'd5205,17'd8040,17'd8040,17'd8339,17'd8340,17'd8190,17'd6,17'd5647,17'd5794,17'd8347,17'd8815,17'd7056,17'd6592,17'd8343,17'd7220,17'd8515,17'd8816,17'd8817,17'd8663,17'd8818,17'd8819,17'd6895,17'd7221,17'd8820,17'd8821,17'd8822,17'd8823,17'd8824,17'd8825,17'd6435,17'd6434,17'd8518,17'd6434,17'd8826,17'd8671,17'd6436,17'd5794,17'd8827,17'd467,17'd285,17'd286,17'd287,17'd287,17'd10,17'd10,17'd467,17'd467,17'd7555,17'd7555,17'd7388,17'd7388,17'd8197,17'd8197,17'd8048,17'd8048,17'd7063,17'd7063,17'd7063,17'd7063,17'd6907,17'd7228,17'd6602,17'd8049,17'd8200,17'd8350,17'd8828,17'd8829,17'd6908,17'd8830,17'd8831,17'd6912,17'd8832,17'd8833,17'd8834,17'd8835,17'd8836,17'd7237,17'd8837,17'd8838,17'd8839,17'd8840,17'd8841,17'd8842,17'd8682,17'd8843,17'd8217,17'd8684,17'd8684,17'd8684,17'd8685,17'd8844,17'd7748,17'd8367,17'd8686,17'd8686,17'd8367,17'd8366,17'd8218,17'd8536,17'd8687,17'd8369,17'd8537,17'd7582,17'd7582,17'd8538,17'd8539,17'd8372,17'd7912,17'd7751,17'd8539,17'd8688,17'd4767,17'd4767,17'd5254,17'd5253,17'd5253,17'd5252,17'd8693,17'd8693,17'd8690,17'd8690,17'd8691,17'd8845,17'd8846,17'd8847,17'd8847,17'd8542,17'd8382,17'd8383,17'd8848,17'd8849,17'd8696,17'd8697,17'd8850,17'd8851,17'd8851,17'd8852,17'd8853,17'd8854,17'd7590,17'd8855,17'd8856,17'd8856,17'd8857,17'd8858,17'd8859,17'd8860,17'd8861,17'd8862,17'd8863,17'd8864,17'd8865,17'd8866,17'd8867,17'd8868,17'd8869,17'd8870,17'd8562,17'd8871,17'd8564,17'd8872,17'd8873,17'd8874,17'd8873,17'd8873,17'd8875,17'd8876,17'd8877,17'd8723,17'd8569,17'd8878,17'd8879,17'd8880,17'd8880,17'd8881,17'd8881,17'd8881,17'd8882,17'd8882,17'd8881,17'd8883,17'd8883,17'd8884,17'd8885,17'd8886,17'd8886,17'd8724,17'd8569,17'd8730,17'd8887,17'd8888,17'd8889,17'd8890,17'd8891,17'd8892,17'd8893,17'd8894,17'd8895,17'd7801,17'd8896,17'd8897,17'd8898,17'd8899,17'd8900,17'd8901,17'd8902,17'd7810,17'd7811,17'd7646,17'd7648,17'd888,17'd542,17'd542,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd132,17'd133,17'd542,17'd542,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd131,17'd8903,17'd8904,17'd8905,17'd8906,17'd8907,17'd8908,17'd8909,17'd6701,17'd8910,17'd8911,17'd6543,17'd8912,17'd7164,17'd8913,17'd8914,17'd8452,17'd7827,17'd7827,17'd8290,17'd8452,17'd8915,17'd8759,17'd8760,17'd8916,17'd8917,17'd8918,17'd8919,17'd8919,17'd8920,17'd8921,17'd8922,17'd8769,17'd8923,17'd8924,17'd8622,17'd8622,17'd8772,17'd8925,17'd8926,17'd8927,17'd8928,17'd8929,17'd8777,17'd8778,17'd8930,17'd7830,17'd7830,17'd7829,17'd7174,17'd7174,17'd7174,17'd7174,17'd7174,17'd7663,17'd7663,17'd7663,17'd8146,17'd8146,17'd7329,17'd7329,17'd7168,17'd6550,17'd8302,17'd8302,17'd8931,17'd7667,17'd8779,17'd8932,17'd7999,17'd8000,17'd8629,17'd8154,17'd8933,17'd7499,17'd7668,17'd8780,17'd8934,17'd7669,17'd7177,17'd6558,17'd8935,17'd8936,17'd8781,17'd7838,17'd8305,17'd8937,17'd8938,17'd8939,17'd8940,17'd8941,17'd8942,17'd8943,17'd8944,17'd8945,17'd8945,17'd4212,17'd8479,17'd4218,17'd8946,17'd8947,17'd8948,17'd8949,17'd225,17'd8950,17'd8951,17'd6726,17'd7362,17'd8952,17'd8953,17'd5783,17'd3407,17'd7860,17'd7347,17'd7348,17'd7688,17'd7687,17'd8171,17'd8795,17'd8795,17'd8491,17'd8954,17'd8796,17'd8955,17'd8798,17'd8956,17'd8957,17'd8958,17'd8959,17'd8802,17'd8960,17'd7517,17'd7347,17'd7689,17'd7519,17'd4718,17'd4871,17'd4567,17'd8803,17'd8961,17'd8323,17'd8962,17'd8963,17'd8808,17'd7866,17'd8964,17'd8326,17'd8654,17'd8329,17'd8329,17'd8501,17'd8654,17'd8654,17'd8327,17'd7873,17'd7874,17'd7698,17'd7034,17'd7034,17'd8810,17'd8810,17'd8965,17'd8966,17'd8967,17'd8334,17'd3073,17'd4714,17'd7537,17'd7537,17'd7538,17'd7538,17'd7705,17'd7705,17'd6416,17'd8187,17'd8187,17'd7365,17'd4729,17'd5958,17'd6581,17'd5958,17'd5958,17'd4882,17'd4423,17'd1810,17'd4084,17'd1243,17'd206,17'd206,17'd971,17'd603,17'd1246,17'd2763
},
'{
17'd8968,17'd8969,17'd7880,17'd8970,17'd8335,17'd8336,17'd7709,17'd7046,17'd5960,17'd5376,17'd4893,17'd2783,17'd2784,17'd1689,17'd17,17'd18,17'd8971,17'd13,17'd0,17'd0,17'd14,17'd4247,17'd7214,17'd7214,17'd7545,17'd4887,17'd2592,17'd2784,17'd2422,17'd1831,17'd1689,17'd0,17'd10,17'd23,17'd4,17'd8,17'd7,17'd5205,17'd8040,17'd8040,17'd8040,17'd8040,17'd8972,17'd7725,17'd7050,17'd7713,17'd8973,17'd6272,17'd6592,17'd8192,17'd8974,17'd8975,17'd8976,17'd8977,17'd8662,17'd8978,17'd8977,17'd8979,17'd6895,17'd8980,17'd8981,17'd8982,17'd8983,17'd8984,17'd8985,17'd6266,17'd6435,17'd7380,17'd8669,17'd8669,17'd8986,17'd8987,17'd5795,17'd5652,17'd285,17'd285,17'd26,17'd27,17'd287,17'd28,17'd27,17'd286,17'd8988,17'd7728,17'd7388,17'd7388,17'd7557,17'd8048,17'd8048,17'd8048,17'd8048,17'd8048,17'd7063,17'd7063,17'd7064,17'd7064,17'd8989,17'd6907,17'd8199,17'd8049,17'd8200,17'd7229,17'd7897,17'd7068,17'd7733,17'd8990,17'd6754,17'd7072,17'd8991,17'd8992,17'd8993,17'd8994,17'd8995,17'd8996,17'd8997,17'd8998,17'd8999,17'd9000,17'd9001,17'd9002,17'd8365,17'd9003,17'd9003,17'd9003,17'd8684,17'd7414,17'd7748,17'd7748,17'd8686,17'd8686,17'd8686,17'd8367,17'd8366,17'd9004,17'd8535,17'd8687,17'd9005,17'd9006,17'd8537,17'd8538,17'd9007,17'd8371,17'd8371,17'd8371,17'd8688,17'd8688,17'd4611,17'd4611,17'd5255,17'd5689,17'd6139,17'd6139,17'd9008,17'd9009,17'd9010,17'd9010,17'd8845,17'd9011,17'd8220,17'd8220,17'd8543,17'd9012,17'd9012,17'd8694,17'd8848,17'd8849,17'd8696,17'd9013,17'd9013,17'd9014,17'd9015,17'd9016,17'd9017,17'd9018,17'd9019,17'd7427,17'd8855,17'd9020,17'd9020,17'd7266,17'd9021,17'd9022,17'd9023,17'd9024,17'd9025,17'd9026,17'd9027,17'd9028,17'd9029,17'd9030,17'd9031,17'd9032,17'd9033,17'd9034,17'd9035,17'd9036,17'd9037,17'd8875,17'd9038,17'd9039,17'd9038,17'd9038,17'd9038,17'd8875,17'd8721,17'd8721,17'd9040,17'd9041,17'd9042,17'd9043,17'd9043,17'd8720,17'd8720,17'd8721,17'd8721,17'd8720,17'd8720,17'd9044,17'd9044,17'd9044,17'd8720,17'd8720,17'd9044,17'd9045,17'd9041,17'd9040,17'd9046,17'd9047,17'd9048,17'd9049,17'd9050,17'd9051,17'd9052,17'd9053,17'd9054,17'd9055,17'd9056,17'd8435,17'd8745,17'd8274,17'd9057,17'd7808,17'd9058,17'd7644,17'd8129,17'd8130,17'd7648,17'd9059,17'd8132,17'd889,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd542,17'd542,17'd542,17'd133,17'd132,17'd135,17'd132,17'd132,17'd132,17'd133,17'd1197,17'd132,17'd9060,17'd9061,17'd9062,17'd3348,17'd9063,17'd9064,17'd8603,17'd9065,17'd9066,17'd9067,17'd6702,17'd6545,17'd6841,17'd7009,17'd8145,17'd8452,17'd9068,17'd8455,17'd8455,17'd9068,17'd8291,17'd8915,17'd9069,17'd9070,17'd8916,17'd9071,17'd9072,17'd9073,17'd9074,17'd9075,17'd9076,17'd9077,17'd9078,17'd8459,17'd9079,17'd8771,17'd9080,17'd8774,17'd8927,17'd9081,17'd9082,17'd9082,17'd9083,17'd9084,17'd9085,17'd9086,17'd9087,17'd9088,17'd9089,17'd9089,17'd9089,17'd7665,17'd7174,17'd7174,17'd7174,17'd7663,17'd7663,17'd7174,17'd7663,17'd7329,17'd7329,17'd7329,17'd7329,17'd6550,17'd6550,17'd6216,17'd6216,17'd7667,17'd7667,17'd7667,17'd6704,17'd8000,17'd6707,17'd9090,17'd8154,17'd9091,17'd7499,17'd8780,17'd7669,17'd7669,17'd6557,17'd6710,17'd7501,17'd7670,17'd9092,17'd8473,17'd9093,17'd8783,17'd7843,17'd9094,17'd9095,17'd9096,17'd9097,17'd8944,17'd8944,17'd6074,17'd4212,17'd7021,17'd4216,17'd9098,17'd9099,17'd9100,17'd9101,17'd9102,17'd1257,17'd9103,17'd9104,17'd9105,17'd7361,17'd9106,17'd3730,17'd9107,17'd8175,17'd7861,17'd9108,17'd8490,17'd8490,17'd8794,17'd8954,17'd8795,17'd8795,17'd8795,17'd7856,17'd9109,17'd8798,17'd9110,17'd9111,17'd9112,17'd9113,17'd9114,17'd9115,17'd8174,17'd7347,17'd7688,17'd7518,17'd4718,17'd4718,17'd9116,17'd7689,17'd9108,17'd8495,17'd8801,17'd8959,17'd9117,17'd9118,17'd8499,17'd8499,17'd8326,17'd8327,17'd8501,17'd8654,17'd9119,17'd8654,17'd8654,17'd8654,17'd8327,17'd8327,17'd7698,17'd8181,17'd9120,17'd8655,17'd9121,17'd3886,17'd9122,17'd8333,17'd4559,17'd9123,17'd7537,17'd7705,17'd9124,17'd9124,17'd7705,17'd7537,17'd7537,17'd7537,17'd6094,17'd6258,17'd4713,17'd5958,17'd6416,17'd6416,17'd5958,17'd4882,17'd4423,17'd1810,17'd2764,17'd1823,17'd2779,17'd643,17'd205,17'd1409,17'd2117,17'd2763
},
'{
17'd8969,17'd9125,17'd7706,17'd8970,17'd8335,17'd7709,17'd7369,17'd5375,17'd5645,17'd4087,17'd3901,17'd2935,17'd1688,17'd1127,17'd17,17'd3905,17'd3430,17'd13,17'd0,17'd0,17'd14,17'd1688,17'd4886,17'd7545,17'd4887,17'd4887,17'd2784,17'd2422,17'd1831,17'd4247,17'd14,17'd12,17'd25,17'd4,17'd8,17'd7,17'd5205,17'd5205,17'd8040,17'd8040,17'd8040,17'd5205,17'd7726,17'd8041,17'd5796,17'd6435,17'd6105,17'd6741,17'd7549,17'd7716,17'd9126,17'd9127,17'd9128,17'd9129,17'd9130,17'd9131,17'd9129,17'd8979,17'd7719,17'd8980,17'd7055,17'd9132,17'd9133,17'd9134,17'd8661,17'd9135,17'd9136,17'd9137,17'd6104,17'd6272,17'd9138,17'd9139,17'd5653,17'd10,17'd980,17'd286,17'd27,17'd28,17'd287,17'd2424,17'd286,17'd286,17'd7728,17'd7728,17'd7388,17'd7557,17'd7557,17'd8048,17'd8048,17'd8048,17'd8048,17'd8048,17'd7063,17'd7063,17'd7064,17'd6907,17'd6906,17'd9140,17'd8199,17'd8200,17'd8201,17'd9141,17'd9142,17'd6910,17'd9143,17'd7071,17'd9144,17'd9145,17'd9146,17'd9147,17'd9148,17'd9149,17'd9150,17'd8997,17'd9151,17'd9152,17'd9153,17'd9154,17'd9155,17'd9156,17'd8217,17'd9003,17'd9003,17'd9003,17'd7749,17'd8366,17'd8367,17'd9157,17'd8686,17'd8367,17'd8367,17'd8366,17'd9004,17'd8536,17'd8687,17'd9158,17'd9006,17'd9159,17'd8538,17'd9007,17'd8371,17'd8371,17'd8371,17'd8539,17'd8688,17'd4611,17'd4611,17'd4767,17'd5255,17'd6139,17'd6139,17'd6139,17'd9008,17'd9009,17'd9160,17'd9010,17'd9160,17'd8074,17'd8220,17'd8381,17'd9012,17'd9012,17'd9012,17'd9161,17'd8849,17'd9162,17'd9013,17'd9163,17'd9014,17'd9164,17'd9016,17'd9165,17'd9018,17'd9019,17'd9166,17'd9167,17'd9168,17'd9169,17'd9170,17'd7764,17'd9171,17'd9172,17'd9173,17'd9174,17'd9175,17'd9176,17'd9177,17'd9178,17'd9179,17'd9180,17'd9181,17'd9182,17'd9183,17'd9184,17'd9185,17'd9186,17'd9187,17'd9188,17'd9038,17'd9039,17'd9038,17'd9038,17'd9038,17'd8873,17'd8873,17'd8873,17'd9189,17'd8874,17'd9190,17'd9191,17'd9192,17'd9192,17'd9193,17'd9038,17'd9038,17'd8874,17'd8874,17'd9189,17'd9189,17'd9043,17'd9189,17'd9189,17'd8720,17'd8720,17'd9189,17'd9189,17'd9194,17'd9195,17'd8731,17'd9196,17'd8250,17'd9197,17'd9198,17'd9199,17'd9200,17'd9201,17'd9202,17'd7969,17'd8436,17'd9203,17'd9204,17'd9205,17'd9206,17'd8902,17'd7481,17'd7978,17'd7812,17'd8444,17'd8132,17'd889,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd542,17'd542,17'd133,17'd132,17'd131,17'd131,17'd132,17'd134,17'd133,17'd134,17'd357,17'd9207,17'd9208,17'd9209,17'd9210,17'd9211,17'd9212,17'd9213,17'd9214,17'd9215,17'd8143,17'd9216,17'd9217,17'd9218,17'd9219,17'd7992,17'd8291,17'd9220,17'd9221,17'd9221,17'd8455,17'd7993,17'd7496,17'd9069,17'd9222,17'd9223,17'd9224,17'd9225,17'd9226,17'd9227,17'd9228,17'd8921,17'd9229,17'd9230,17'd8298,17'd9231,17'd8462,17'd8623,17'd9232,17'd9233,17'd9082,17'd9234,17'd9234,17'd9235,17'd9082,17'd9084,17'd9085,17'd9236,17'd9237,17'd9238,17'd9088,17'd9089,17'd7665,17'd7174,17'd7174,17'd7174,17'd7663,17'd7663,17'd7663,17'd7663,17'd6849,17'd6849,17'd7329,17'd7329,17'd7168,17'd7168,17'd6550,17'd6215,17'd7667,17'd7667,17'd7667,17'd7176,17'd7999,17'd7999,17'd8154,17'd8154,17'd7668,17'd7668,17'd7668,17'd7668,17'd7669,17'd7669,17'd6709,17'd6559,17'd8472,17'd8472,17'd8630,17'd8474,17'd9239,17'd8938,17'd9240,17'd8940,17'd9241,17'd9242,17'd4857,17'd8943,17'd8943,17'd8945,17'd4701,17'd9243,17'd4387,17'd9244,17'd3703,17'd9245,17'd9246,17'd9247,17'd7850,17'd3422,17'd9248,17'd6884,17'd7207,17'd3237,17'd9249,17'd3576,17'd7861,17'd9250,17'd9251,17'd7687,17'd8794,17'd9252,17'd8795,17'd9253,17'd8795,17'd8170,17'd8954,17'd8955,17'd9254,17'd9255,17'd9256,17'd9257,17'd9115,17'd9115,17'd8495,17'd8960,17'd7348,17'd7689,17'd4871,17'd4718,17'd9116,17'd7689,17'd9108,17'd9250,17'd8648,17'd8805,17'd8963,17'd9258,17'd7866,17'd8499,17'd9259,17'd8809,17'd8327,17'd8654,17'd8654,17'd9119,17'd8654,17'd8654,17'd8327,17'd8327,17'd7698,17'd7698,17'd9120,17'd7034,17'd9260,17'd3727,17'd3731,17'd9122,17'd8184,17'd6889,17'd6416,17'd9261,17'd9124,17'd9124,17'd7705,17'd7537,17'd7537,17'd7537,17'd6094,17'd6258,17'd4713,17'd5958,17'd6416,17'd6416,17'd5958,17'd4882,17'd4423,17'd4085,17'd6407,17'd1823,17'd2779,17'd643,17'd205,17'd1099,17'd1246,17'd2763
},
'{
17'd8509,17'd7883,17'd8508,17'd9262,17'd8508,17'd7883,17'd7544,17'd5960,17'd5201,17'd4244,17'd2934,17'd2422,17'd1127,17'd466,17'd13,17'd13,17'd2,17'd0,17'd0,17'd2,17'd6419,17'd4886,17'd4886,17'd7711,17'd4887,17'd4887,17'd2422,17'd2422,17'd4247,17'd466,17'd12,17'd806,17'd4,17'd6,17'd7,17'd7,17'd5205,17'd5205,17'd8340,17'd8340,17'd8190,17'd8190,17'd9263,17'd6098,17'd6435,17'd8669,17'd9132,17'd8666,17'd9264,17'd9265,17'd8663,17'd9266,17'd9267,17'd8818,17'd8976,17'd9268,17'd7377,17'd7377,17'd9269,17'd8346,17'd9270,17'd6272,17'd9271,17'd8973,17'd6596,17'd8973,17'd7057,17'd6595,17'd6272,17'd9272,17'd9273,17'd9274,17'd5969,17'd18,17'd652,17'd28,17'd28,17'd28,17'd6902,17'd9275,17'd2424,17'd287,17'd7061,17'd7061,17'd9276,17'd9276,17'd6747,17'd6747,17'd7063,17'd7063,17'd7063,17'd7063,17'd7228,17'd9277,17'd8049,17'd8199,17'd9140,17'd9140,17'd9278,17'd7229,17'd8051,17'd9279,17'd9280,17'd9281,17'd9282,17'd9283,17'd9145,17'd9284,17'd9285,17'd9286,17'd9287,17'd9288,17'd9289,17'd9290,17'd9291,17'd9292,17'd9293,17'd9294,17'd9295,17'd8686,17'd9296,17'd9296,17'd9297,17'd7580,17'd8684,17'd8367,17'd9298,17'd9299,17'd8367,17'd8366,17'd9004,17'd9004,17'd8535,17'd8687,17'd9158,17'd9159,17'd8537,17'd9300,17'd9007,17'd9301,17'd8372,17'd8371,17'd8539,17'd8688,17'd4611,17'd9302,17'd4927,17'd5255,17'd6139,17'd9303,17'd9303,17'd6138,17'd9009,17'd9009,17'd9009,17'd9009,17'd9008,17'd9304,17'd9305,17'd9305,17'd9012,17'd9306,17'd9307,17'd9308,17'd9013,17'd9013,17'd9014,17'd9014,17'd9309,17'd9309,17'd9310,17'd9311,17'd9312,17'd9166,17'd9313,17'd9314,17'd9315,17'd9316,17'd9317,17'd9318,17'd9319,17'd9320,17'd9321,17'd9322,17'd9323,17'd9324,17'd9325,17'd9326,17'd9327,17'd9328,17'd9329,17'd9330,17'd9331,17'd9332,17'd9333,17'd9334,17'd9335,17'd9335,17'd9335,17'd9335,17'd9335,17'd9336,17'd9336,17'd9337,17'd9338,17'd9339,17'd9340,17'd9341,17'd9342,17'd9342,17'd9343,17'd9343,17'd9343,17'd9343,17'd9343,17'd9344,17'd9345,17'd9344,17'd9346,17'd9339,17'd9347,17'd9192,17'd8873,17'd8873,17'd9189,17'd9189,17'd9189,17'd9041,17'd9348,17'd8726,17'd9349,17'd8249,17'd9350,17'd9351,17'd9352,17'd9353,17'd7633,17'd7966,17'd9354,17'd9355,17'd9356,17'd9205,17'd9357,17'd9358,17'd8128,17'd8279,17'd9359,17'd9360,17'd6830,17'd888,17'd542,17'd542,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd542,17'd542,17'd133,17'd132,17'd131,17'd131,17'd132,17'd1197,17'd132,17'd132,17'd3996,17'd9361,17'd9362,17'd9363,17'd9364,17'd9365,17'd9366,17'd9367,17'd6700,17'd9215,17'd7163,17'd6841,17'd9368,17'd9369,17'd7990,17'd7827,17'd8291,17'd8455,17'd9370,17'd9370,17'd9371,17'd7993,17'd9372,17'd9373,17'd8916,17'd9374,17'd9375,17'd9376,17'd9377,17'd9378,17'd9228,17'd8921,17'd8296,17'd9379,17'd9380,17'd8462,17'd9381,17'd9382,17'd8776,17'd9232,17'd9383,17'd9082,17'd9384,17'd9385,17'd9385,17'd9386,17'd9387,17'd9388,17'd9389,17'd9390,17'd9391,17'd9087,17'd9392,17'd9393,17'd7665,17'd7174,17'd7174,17'd7663,17'd7663,17'd7663,17'd6848,17'd6848,17'd6849,17'd7329,17'd7329,17'd7991,17'd7168,17'd7168,17'd7168,17'd6550,17'd7667,17'd7667,17'd5918,17'd5918,17'd6218,17'd6707,17'd9394,17'd9394,17'd7499,17'd7499,17'd7668,17'd7669,17'd6557,17'd6557,17'd6558,17'd7011,17'd6223,17'd8630,17'd9395,17'd9396,17'd7017,17'd9094,17'd9095,17'd9397,17'd9398,17'd8943,17'd8006,17'd9097,17'd5345,17'd9399,17'd5928,17'd9400,17'd9401,17'd4053,17'd6082,17'd9402,17'd9403,17'd9404,17'd3422,17'd3894,17'd3414,17'd3584,17'd3413,17'd5041,17'd4411,17'd8322,17'd8804,17'd8804,17'd8490,17'd7687,17'd8019,17'd9405,17'd8795,17'd8491,17'd8796,17'd8797,17'd9406,17'd8956,17'd9111,17'd8957,17'd9407,17'd9408,17'd8495,17'd9409,17'd7347,17'd7348,17'd7518,17'd7519,17'd7519,17'd7689,17'd9108,17'd8496,17'd8805,17'd9410,17'd8963,17'd8806,17'd8026,17'd7691,17'd9411,17'd9412,17'd8028,17'd7873,17'd8654,17'd9119,17'd8654,17'd8654,17'd8327,17'd8327,17'd8327,17'd8327,17'd7698,17'd8330,17'd7033,17'd5186,17'd8182,17'd8658,17'd9413,17'd6727,17'd6416,17'd9414,17'd7705,17'd9261,17'd7705,17'd7537,17'd7537,17'd7537,17'd6094,17'd6258,17'd4713,17'd5958,17'd6416,17'd6416,17'd8186,17'd5958,17'd4728,17'd1810,17'd2764,17'd1667,17'd206,17'd643,17'd205,17'd1409,17'd2117,17'd2763
},
'{
17'd7709,17'd8508,17'd8508,17'd9262,17'd7709,17'd7046,17'd5959,17'd5201,17'd4244,17'd6420,17'd2422,17'd1689,17'd1127,17'd2,17'd13,17'd13,17'd0,17'd0,17'd2,17'd14,17'd5196,17'd4886,17'd7711,17'd7711,17'd4887,17'd4887,17'd3252,17'd1831,17'd2595,17'd12,17'd806,17'd2933,17'd6,17'd6,17'd7,17'd7,17'd5205,17'd5205,17'd8040,17'd8190,17'd5205,17'd7,17'd6097,17'd6588,17'd6434,17'd9415,17'd9416,17'd8517,17'd8664,17'd9417,17'd9266,17'd9131,17'd8663,17'd8818,17'd9128,17'd9267,17'd7377,17'd9418,17'd8345,17'd8822,17'd9419,17'd9420,17'd8824,17'd5962,17'd8670,17'd7380,17'd6595,17'd6595,17'd7885,17'd6272,17'd9421,17'd9422,17'd1277,17'd18,17'd652,17'd288,17'd288,17'd29,17'd4430,17'd6744,17'd2424,17'd287,17'd7061,17'd7728,17'd7556,17'd9276,17'd6747,17'd6747,17'd7063,17'd7063,17'd7063,17'd7063,17'd9277,17'd9277,17'd8049,17'd8199,17'd9140,17'd9278,17'd8828,17'd6908,17'd9279,17'd9143,17'd6911,17'd8354,17'd9283,17'd9423,17'd9284,17'd9424,17'd9425,17'd9287,17'd9426,17'd9427,17'd9428,17'd9429,17'd9430,17'd9431,17'd9432,17'd9433,17'd9434,17'd9435,17'd9436,17'd9296,17'd7749,17'd8684,17'd8366,17'd9437,17'd9437,17'd9438,17'd8366,17'd9004,17'd9004,17'd9439,17'd8687,17'd9158,17'd9159,17'd9159,17'd9440,17'd9300,17'd9007,17'd9301,17'd8372,17'd8371,17'd8539,17'd4611,17'd9302,17'd4927,17'd5255,17'd5689,17'd6139,17'd9303,17'd6138,17'd6138,17'd9009,17'd9009,17'd9008,17'd9008,17'd9304,17'd9441,17'd9442,17'd9306,17'd9307,17'd9307,17'd9308,17'd9443,17'd9013,17'd9163,17'd9164,17'd9164,17'd9444,17'd9445,17'd9311,17'd9446,17'd9166,17'd9447,17'd9314,17'd9020,17'd9448,17'd9449,17'd9450,17'd9451,17'd9452,17'd9453,17'd9454,17'd9455,17'd9456,17'd9457,17'd9458,17'd9459,17'd9460,17'd9461,17'd9462,17'd9463,17'd9464,17'd9465,17'd9466,17'd9466,17'd9467,17'd9335,17'd9335,17'd9468,17'd9468,17'd9469,17'd9470,17'd9470,17'd9471,17'd9472,17'd9473,17'd9473,17'd9474,17'd9475,17'd9475,17'd9476,17'd9476,17'd9476,17'd9477,17'd9478,17'd9478,17'd9479,17'd9480,17'd9346,17'd9339,17'd9347,17'd8874,17'd8874,17'd9481,17'd9481,17'd9043,17'd9043,17'd9045,17'd8881,17'd9482,17'd9483,17'd9484,17'd9485,17'd9486,17'd9487,17'd9488,17'd9489,17'd9490,17'd9491,17'd9492,17'd9493,17'd9494,17'd7809,17'd8128,17'd9495,17'd9359,17'd9360,17'd6529,17'd6830,17'd542,17'd542,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd542,17'd133,17'd132,17'd132,17'd131,17'd131,17'd132,17'd1197,17'd132,17'd131,17'd3811,17'd7650,17'd9496,17'd9497,17'd7985,17'd9498,17'd9499,17'd9500,17'd9501,17'd9502,17'd9503,17'd6842,17'd9369,17'd7825,17'd7992,17'd7172,17'd7993,17'd9371,17'd9504,17'd9370,17'd9505,17'd8761,17'd9506,17'd8916,17'd9374,17'd9507,17'd9508,17'd9509,17'd9510,17'd9511,17'd9512,17'd9513,17'd8296,17'd9379,17'd9514,17'd8462,17'd8623,17'd9515,17'd9232,17'd9232,17'd9516,17'd9383,17'd9517,17'd9517,17'd9518,17'd9518,17'd9518,17'd9387,17'd9388,17'd9519,17'd9520,17'd9086,17'd9237,17'd9392,17'd9521,17'd7665,17'd7665,17'd7174,17'd7663,17'd7663,17'd6848,17'd6848,17'd6849,17'd7329,17'd7329,17'd9522,17'd7168,17'd7168,17'd7168,17'd6550,17'd8302,17'd7667,17'd7667,17'd5918,17'd9523,17'd6553,17'd9090,17'd9090,17'd8304,17'd7499,17'd7668,17'd8780,17'd7669,17'd7500,17'd7500,17'd7177,17'd6393,17'd6223,17'd8473,17'd8305,17'd9524,17'd7017,17'd8308,17'd9525,17'd8941,17'd9526,17'd9527,17'd9097,17'd9097,17'd4701,17'd5769,17'd9528,17'd6079,17'd9529,17'd9530,17'd5494,17'd6238,17'd5775,17'd9531,17'd4241,17'd3239,17'd9532,17'd9533,17'd3732,17'd6874,17'd4411,17'd9108,17'd9250,17'd8490,17'd8490,17'd7856,17'd8171,17'd8491,17'd8795,17'd9534,17'd8796,17'd9535,17'd9536,17'd9255,17'd9537,17'd9538,17'd9539,17'd9540,17'd9409,17'd9250,17'd7347,17'd7689,17'd7519,17'd7349,17'd7518,17'd9108,17'd8322,17'd8323,17'd9410,17'd9541,17'd8806,17'd8498,17'd7691,17'd9411,17'd9542,17'd7867,17'd8327,17'd8501,17'd9119,17'd8654,17'd8654,17'd8327,17'd8327,17'd8327,17'd8327,17'd7698,17'd7698,17'd7034,17'd6876,17'd5950,17'd8182,17'd8332,17'd9543,17'd6727,17'd9544,17'd7705,17'd9261,17'd7705,17'd7537,17'd7537,17'd7537,17'd6094,17'd6258,17'd4882,17'd5958,17'd6416,17'd6416,17'd8186,17'd8186,17'd4882,17'd4085,17'd6407,17'd1667,17'd206,17'd644,17'd205,17'd1686,17'd2116,17'd2763
},
'{
17'd7709,17'd8508,17'd8508,17'd8508,17'd7369,17'd5375,17'd5376,17'd4087,17'd4088,17'd4246,17'd1688,17'd1127,17'd2,17'd2,17'd2,17'd2,17'd1,17'd0,17'd14,17'd1127,17'd5196,17'd4886,17'd7711,17'd4577,17'd4887,17'd4887,17'd2422,17'd4247,17'd13,17'd806,17'd23,17'd5,17'd6,17'd5205,17'd5205,17'd5205,17'd5205,17'd5205,17'd5205,17'd5205,17'd8972,17'd7725,17'd6098,17'd9135,17'd9545,17'd7714,17'd8517,17'd7220,17'd9546,17'd8662,17'd9547,17'd8662,17'd8978,17'd9131,17'd9268,17'd9548,17'd9418,17'd9549,17'd7055,17'd9550,17'd9272,17'd7057,17'd6434,17'd6596,17'd7892,17'd9137,17'd6595,17'd9551,17'd7885,17'd9552,17'd9553,17'd1415,17'd16,17'd18,17'd29,17'd2118,17'd9554,17'd4431,17'd4430,17'd6744,17'd6902,17'd6902,17'd9555,17'd9555,17'd6904,17'd6904,17'd6747,17'd7063,17'd7063,17'd7063,17'd7228,17'd7228,17'd8049,17'd8049,17'd8200,17'd8200,17'd9278,17'd8828,17'd7732,17'd9556,17'd7070,17'd9557,17'd9558,17'd9559,17'd9145,17'd9284,17'd9424,17'd9147,17'd9560,17'd9561,17'd8997,17'd9562,17'd9563,17'd9564,17'd9000,17'd9565,17'd9566,17'd9567,17'd9568,17'd9434,17'd9569,17'd9570,17'd8686,17'd8686,17'd9571,17'd9572,17'd9437,17'd8367,17'd8366,17'd7086,17'd8536,17'd9573,17'd9158,17'd9574,17'd9159,17'd9300,17'd8538,17'd9007,17'd9575,17'd9575,17'd8067,17'd8066,17'd4611,17'd4611,17'd7750,17'd6468,17'd6140,17'd6140,17'd6139,17'd6138,17'd6138,17'd6138,17'd9009,17'd9009,17'd9576,17'd9304,17'd9577,17'd9578,17'd9578,17'd9579,17'd9579,17'd9580,17'd9580,17'd9580,17'd9581,17'd9582,17'd9309,17'd9583,17'd9584,17'd9584,17'd9585,17'd9586,17'd9447,17'd9587,17'd9588,17'd9589,17'd9590,17'd9591,17'd9451,17'd9592,17'd9593,17'd9594,17'd9595,17'd9596,17'd9597,17'd9598,17'd9599,17'd9600,17'd9601,17'd9602,17'd9603,17'd9604,17'd9605,17'd9606,17'd9607,17'd9607,17'd9607,17'd9608,17'd9608,17'd9608,17'd9608,17'd9606,17'd9609,17'd9475,17'd9610,17'd9611,17'd9612,17'd9613,17'd9614,17'd9615,17'd9615,17'd9615,17'd9614,17'd9616,17'd9617,17'd9618,17'd9618,17'd9619,17'd9479,17'd9620,17'd9346,17'd9347,17'd8874,17'd8874,17'd9191,17'd9191,17'd9043,17'd9043,17'd9621,17'd8882,17'd9482,17'd8247,17'd8418,17'd9622,17'd9623,17'd9624,17'd7795,17'd9625,17'd9626,17'd9627,17'd9628,17'd9629,17'd9494,17'd9630,17'd9631,17'd8750,17'd8130,17'd9360,17'd6529,17'd6830,17'd889,17'd542,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd542,17'd133,17'd132,17'd132,17'd131,17'd135,17'd133,17'd1197,17'd132,17'd131,17'd3026,17'd9632,17'd9633,17'd9634,17'd9635,17'd9636,17'd8286,17'd6837,17'd9637,17'd9638,17'd8608,17'd7165,17'd8913,17'd7990,17'd7827,17'd7173,17'd7172,17'd9371,17'd9639,17'd9640,17'd9641,17'd9642,17'd8917,17'd9374,17'd9507,17'd9643,17'd9644,17'd9645,17'd9646,17'd9647,17'd9076,17'd9648,17'd9649,17'd8297,17'd9650,17'd8463,17'd8625,17'd8623,17'd8776,17'd9232,17'd9516,17'd9383,17'd9651,17'd9651,17'd9517,17'd9651,17'd9518,17'd9651,17'd9652,17'd9653,17'd9654,17'd9655,17'd9656,17'd9087,17'd9392,17'd9521,17'd9393,17'd8301,17'd7665,17'd7174,17'd6848,17'd8146,17'd8146,17'd8146,17'd8146,17'd8146,17'd7329,17'd7329,17'd6849,17'd6550,17'd6550,17'd6215,17'd6215,17'd5917,17'd5918,17'd6704,17'd8000,17'd6707,17'd9090,17'd9090,17'd9657,17'd7668,17'd7668,17'd7669,17'd7669,17'd7500,17'd7500,17'd6558,17'd8472,17'd6394,17'd9395,17'd9524,17'd6858,17'd9658,17'd8476,17'd5018,17'd5487,17'd9659,17'd8943,17'd4382,17'd5768,17'd9660,17'd4045,17'd5022,17'd9661,17'd4225,17'd3568,17'd1120,17'd2578,17'd3240,17'd3733,17'd9662,17'd9663,17'd4077,17'd3727,17'd9664,17'd8322,17'd9250,17'd7347,17'd7347,17'd7686,17'd7856,17'd8491,17'd8795,17'd8795,17'd8019,17'd8797,17'd8798,17'd9254,17'd8956,17'd9256,17'd9538,17'd9665,17'd8495,17'd8804,17'd9250,17'd7688,17'd7518,17'd7519,17'd7518,17'd8322,17'd8322,17'd8323,17'd9410,17'd9541,17'd8962,17'd9666,17'd8650,17'd9411,17'd9542,17'd9412,17'd9667,17'd8654,17'd8654,17'd8654,17'd8654,17'd8654,17'd8654,17'd8327,17'd8028,17'd8181,17'd8181,17'd7698,17'd9668,17'd8655,17'd8504,17'd8658,17'd9669,17'd9670,17'd8187,17'd7705,17'd9261,17'd7705,17'd7537,17'd7537,17'd7537,17'd6890,17'd6094,17'd4882,17'd5958,17'd6416,17'd6416,17'd6416,17'd5958,17'd4728,17'd1810,17'd2764,17'd1667,17'd643,17'd644,17'd1966,17'd1686,17'd2116,17'd9671
},
'{
17'd7709,17'd7709,17'd7709,17'd7369,17'd5375,17'd5790,17'd5202,17'd3903,17'd4733,17'd7545,17'd1127,17'd14,17'd2,17'd2,17'd2,17'd0,17'd0,17'd0,17'd14,17'd1127,17'd5196,17'd7711,17'd4577,17'd4577,17'd4887,17'd7545,17'd1688,17'd1127,17'd12,17'd2933,17'd4,17'd6,17'd3753,17'd5205,17'd5205,17'd5205,17'd5205,17'd3753,17'd5205,17'd5205,17'd9672,17'd8196,17'd9673,17'd7223,17'd8823,17'd6897,17'd8192,17'd8515,17'd9265,17'd9131,17'd9674,17'd9675,17'd9676,17'd9677,17'd9129,17'd9678,17'd9679,17'd8346,17'd9680,17'd9681,17'd9682,17'd6434,17'd6100,17'd7892,17'd9137,17'd6272,17'd7885,17'd9551,17'd9683,17'd9684,17'd2596,17'd17,17'd17,17'd16,17'd981,17'd981,17'd9554,17'd3907,17'd4430,17'd6902,17'd6744,17'd6902,17'd9685,17'd9555,17'd6599,17'd6599,17'd6747,17'd7390,17'd7063,17'd7063,17'd7228,17'd7228,17'd8049,17'd8049,17'd8200,17'd8200,17'd7229,17'd7067,17'd9556,17'd9686,17'd9687,17'd9558,17'd9559,17'd9688,17'd9689,17'd9690,17'd9691,17'd9148,17'd9149,17'd9692,17'd9693,17'd9694,17'd9695,17'd9696,17'd9697,17'd9698,17'd9433,17'd9567,17'd9699,17'd9700,17'd9569,17'd9435,17'd9435,17'd9438,17'd9571,17'd9572,17'd8367,17'd9004,17'd7086,17'd9701,17'd9573,17'd9702,17'd9702,17'd9300,17'd9300,17'd9703,17'd9007,17'd9301,17'd9575,17'd9704,17'd8066,17'd4611,17'd4611,17'd9302,17'd6468,17'd6141,17'd6140,17'd6305,17'd6138,17'd6138,17'd6138,17'd6138,17'd9008,17'd9008,17'd9304,17'd9441,17'd9578,17'd9578,17'd9705,17'd9705,17'd9580,17'd9580,17'd9580,17'd9706,17'd9582,17'd9707,17'd9583,17'd9444,17'd9584,17'd9585,17'd9446,17'd9708,17'd9587,17'd9709,17'd9589,17'd9590,17'd9710,17'd9711,17'd9712,17'd9713,17'd9714,17'd9715,17'd9716,17'd9717,17'd9718,17'd9719,17'd9720,17'd9721,17'd9722,17'd9723,17'd9724,17'd9725,17'd9726,17'd9727,17'd9727,17'd9728,17'd9607,17'd9607,17'd9607,17'd9606,17'd9729,17'd9730,17'd9731,17'd9614,17'd9614,17'd9732,17'd9732,17'd9733,17'd9734,17'd9735,17'd9735,17'd9734,17'd9733,17'd9736,17'd9737,17'd9738,17'd9739,17'd9740,17'd9741,17'd9742,17'd9620,17'd9339,17'd9743,17'd8874,17'd9339,17'd9339,17'd9189,17'd9043,17'd9045,17'd8879,17'd9482,17'd9744,17'd9745,17'd7949,17'd9746,17'd9747,17'd9748,17'd9749,17'd9750,17'd9751,17'd9752,17'd9753,17'd9754,17'd9630,17'd9631,17'd9755,17'd9756,17'd7812,17'd8444,17'd6529,17'd889,17'd542,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd131,17'd135,17'd133,17'd133,17'd132,17'd3996,17'd9757,17'd9758,17'd9759,17'd9760,17'd9761,17'd9762,17'd9763,17'd9764,17'd8911,17'd7659,17'd7823,17'd7824,17'd9765,17'd9068,17'd7993,17'd7173,17'd7835,17'd9766,17'd9371,17'd9505,17'd9767,17'd9374,17'd9768,17'd9769,17'd9375,17'd9375,17'd9644,17'd9770,17'd9771,17'd9772,17'd9773,17'd9774,17'd9775,17'd9776,17'd9777,17'd9514,17'd8625,17'd8625,17'd9778,17'd8776,17'd9779,17'd9516,17'd9651,17'd9651,17'd9517,17'd9780,17'd9518,17'd9651,17'd9781,17'd9781,17'd9782,17'd9654,17'd9520,17'd9783,17'd9087,17'd9521,17'd9393,17'd8301,17'd7665,17'd7665,17'd7175,17'd6848,17'd8146,17'd8146,17'd8146,17'd8146,17'd7329,17'd7329,17'd7329,17'd6849,17'd6550,17'd6550,17'd6550,17'd6216,17'd7176,17'd6704,17'd7999,17'd8000,17'd9090,17'd9394,17'd9657,17'd8304,17'd7668,17'd8780,17'd7669,17'd7669,17'd7500,17'd7177,17'd6558,17'd6559,17'd9092,17'd8305,17'd8782,17'd9784,17'd9658,17'd9525,17'd9785,17'd9786,17'd8161,17'd9097,17'd5345,17'd9787,17'd4215,17'd5177,17'd9788,17'd9789,17'd4864,17'd3711,17'd627,17'd2924,17'd9790,17'd3733,17'd9791,17'd7207,17'd8332,17'd9792,17'd4411,17'd9108,17'd7347,17'd7517,17'd7858,17'd7686,17'd8171,17'd8491,17'd8795,17'd8795,17'd8796,17'd8955,17'd9793,17'd9254,17'd9794,17'd9795,17'd9796,17'd9665,17'd9797,17'd8804,17'd8490,17'd7688,17'd7518,17'd7518,17'd8322,17'd8322,17'd8323,17'd8648,17'd9541,17'd9541,17'd9666,17'd8962,17'd9411,17'd9542,17'd8652,17'd9798,17'd9119,17'd8654,17'd8654,17'd8654,17'd9119,17'd9119,17'd8028,17'd8028,17'd8181,17'd8181,17'd7698,17'd9799,17'd9800,17'd9801,17'd9802,17'd9803,17'd9804,17'd9414,17'd7705,17'd7705,17'd7705,17'd7537,17'd7537,17'd7537,17'd6890,17'd6094,17'd5958,17'd6581,17'd6416,17'd6416,17'd6416,17'd6416,17'd4882,17'd4085,17'd6407,17'd4084,17'd643,17'd644,17'd1966,17'd1098,17'd2116,17'd9671
},
'{
17'd7709,17'd7883,17'd7883,17'd7046,17'd6261,17'd5377,17'd4736,17'd4088,17'd4887,17'd4886,17'd1127,17'd2,17'd2,17'd2,17'd15,17'd15,17'd15,17'd14,17'd1127,17'd1127,17'd5196,17'd7711,17'd4577,17'd4887,17'd4887,17'd7711,17'd1967,17'd0,17'd806,17'd4242,17'd6,17'd5205,17'd8040,17'd8040,17'd5205,17'd5205,17'd7,17'd7,17'd5205,17'd5205,17'd9805,17'd9806,17'd8347,17'd9136,17'd8342,17'd8343,17'd7718,17'd8512,17'd8818,17'd9266,17'd9807,17'd9674,17'd9808,17'd9809,17'd8514,17'd9810,17'd9811,17'd8342,17'd6595,17'd7057,17'd8815,17'd8042,17'd9812,17'd9813,17'd8511,17'd6595,17'd7885,17'd6268,17'd9814,17'd9815,17'd1414,17'd16,17'd289,17'd29,17'd809,17'd31,17'd9816,17'd9554,17'd4430,17'd7061,17'd6744,17'd6902,17'd9555,17'd9555,17'd6904,17'd6904,17'd9817,17'd7228,17'd7228,17'd7228,17'd7228,17'd7228,17'd6602,17'd6602,17'd7393,17'd7229,17'd7067,17'd9818,17'd8830,17'd9819,17'd9820,17'd9821,17'd9822,17'd9823,17'd9824,17'd9825,17'd9826,17'd9827,17'd9828,17'd9829,17'd9830,17'd9831,17'd9832,17'd9833,17'd9834,17'd9835,17'd9836,17'd9837,17'd9700,17'd9838,17'd9838,17'd9839,17'd9840,17'd9841,17'd9571,17'd9437,17'd9004,17'd8535,17'd8536,17'd9573,17'd9158,17'd9574,17'd9159,17'd9703,17'd9703,17'd9704,17'd9704,17'd9575,17'd8371,17'd8371,17'd4611,17'd4767,17'd4767,17'd4927,17'd6141,17'd7417,17'd6140,17'd6140,17'd6139,17'd6138,17'd8693,17'd8846,17'd8846,17'd9842,17'd9304,17'd9441,17'd9578,17'd9843,17'd9844,17'd9844,17'd9845,17'd9845,17'd9846,17'd9847,17'd9848,17'd9849,17'd9444,17'd9850,17'd9584,17'd9585,17'd9312,17'd9447,17'd9709,17'd9588,17'd9851,17'd9852,17'd9853,17'd9712,17'd9854,17'd9855,17'd9856,17'd9857,17'd9858,17'd9859,17'd9860,17'd9861,17'd9862,17'd9863,17'd9864,17'd9865,17'd9866,17'd9725,17'd9867,17'd9867,17'd9868,17'd9869,17'd9727,17'd9729,17'd9870,17'd9871,17'd9731,17'd9872,17'd9734,17'd9873,17'd9874,17'd9874,17'd9875,17'd9876,17'd9877,17'd9878,17'd9878,17'd9879,17'd9880,17'd9881,17'd9736,17'd9882,17'd9739,17'd9883,17'd9884,17'd9885,17'd9620,17'd9346,17'd9743,17'd9743,17'd9346,17'd9339,17'd9189,17'd8720,17'd9348,17'd8879,17'd9886,17'd9887,17'd9888,17'd9889,17'd9890,17'd9891,17'd9892,17'd9893,17'd9894,17'd9895,17'd8436,17'd9896,17'd9897,17'd9898,17'd9631,17'd9899,17'd7978,17'd7647,17'd9059,17'd6529,17'd8132,17'd889,17'd133,17'd133,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd131,17'd135,17'd542,17'd133,17'd132,17'd5311,17'd9900,17'd9901,17'd9363,17'd9902,17'd9903,17'd9904,17'd9905,17'd6380,17'd9906,17'd9907,17'd7823,17'd9908,17'd9909,17'd9910,17'd8915,17'd7496,17'd7835,17'd9911,17'd8455,17'd8611,17'd9912,17'd9913,17'd9914,17'd9915,17'd9916,17'd9917,17'd9918,17'd9919,17'd8618,17'd9920,17'd9921,17'd9922,17'd9923,17'd9924,17'd9925,17'd9926,17'd9926,17'd8623,17'd9927,17'd8776,17'd9782,17'd9085,17'd9516,17'd9383,17'd9517,17'd9780,17'd9928,17'd9928,17'd9928,17'd9082,17'd9929,17'd9388,17'd9654,17'd9520,17'd9391,17'd9087,17'd9392,17'd9393,17'd7665,17'd7665,17'd7175,17'd6848,17'd6848,17'd8146,17'd8146,17'd8146,17'd9930,17'd9930,17'd7329,17'd7329,17'd7329,17'd6550,17'd6550,17'd6216,17'd6850,17'd7176,17'd9523,17'd7999,17'd9931,17'd9932,17'd9090,17'd9090,17'd7668,17'd7668,17'd9933,17'd9933,17'd9934,17'd9934,17'd9934,17'd6557,17'd6558,17'd6224,17'd8473,17'd9239,17'd8938,17'd9658,17'd9935,17'd9936,17'd9527,17'd9097,17'd5488,17'd9937,17'd9938,17'd9939,17'd9940,17'd9941,17'd4709,17'd3711,17'd609,17'd935,17'd9942,17'd9943,17'd5955,17'd3889,17'd7360,17'd8792,17'd6874,17'd3578,17'd8022,17'd8174,17'd8021,17'd7686,17'd9944,17'd9945,17'd8795,17'd9253,17'd8796,17'd8797,17'd9946,17'd9254,17'd9947,17'd9948,17'd9949,17'd9538,17'd9950,17'd8495,17'd7517,17'd7347,17'd7348,17'd7195,17'd7860,17'd8322,17'd8323,17'd8648,17'd9951,17'd9952,17'd9541,17'd9541,17'd9953,17'd7864,17'd8652,17'd9412,17'd8500,17'd9954,17'd9119,17'd9119,17'd9119,17'd9119,17'd8809,17'd8809,17'd8809,17'd8809,17'd9955,17'd8181,17'd9956,17'd8655,17'd8656,17'd9957,17'd9669,17'd9958,17'd9544,17'd7705,17'd7705,17'd7537,17'd7537,17'd7537,17'd6890,17'd6094,17'd5958,17'd6581,17'd6416,17'd6416,17'd6416,17'd6581,17'd4728,17'd1810,17'd2922,17'd4084,17'd644,17'd644,17'd1966,17'd1098,17'd2116,17'd9671
},
'{
17'd7883,17'd7369,17'd7046,17'd5375,17'd5960,17'd9959,17'd9960,17'd4733,17'd7711,17'd6419,17'd14,17'd2,17'd2,17'd2,17'd15,17'd15,17'd14,17'd14,17'd1127,17'd1688,17'd6583,17'd7711,17'd4577,17'd4887,17'd7545,17'd4886,17'd15,17'd3,17'd2933,17'd4242,17'd6,17'd8190,17'd8040,17'd8340,17'd8190,17'd5205,17'd7,17'd7,17'd7,17'd7374,17'd9961,17'd9673,17'd9135,17'd8511,17'd9962,17'd7549,17'd9963,17'd8513,17'd8976,17'd9127,17'd8662,17'd9809,17'd8817,17'd8978,17'd9964,17'd9269,17'd7715,17'd9550,17'd9420,17'd9965,17'd8042,17'd6105,17'd9271,17'd6105,17'd9420,17'd9966,17'd9415,17'd9967,17'd9968,17'd3750,17'd9969,17'd1415,17'd981,17'd2118,17'd31,17'd1129,17'd3754,17'd3907,17'd4091,17'd4430,17'd6902,17'd6902,17'd6903,17'd6903,17'd9970,17'd9970,17'd7228,17'd7228,17'd7228,17'd7228,17'd7228,17'd6602,17'd7065,17'd7393,17'd7229,17'd7897,17'd9142,17'd9971,17'd8990,17'd9557,17'd9972,17'd9973,17'd9974,17'd9975,17'd9976,17'd9826,17'd9977,17'd9150,17'd9829,17'd9978,17'd9979,17'd9980,17'd9981,17'd9982,17'd9983,17'd9983,17'd9836,17'd9837,17'd9984,17'd9838,17'd9839,17'd9840,17'd9840,17'd9841,17'd9438,17'd9437,17'd9004,17'd8536,17'd9573,17'd9702,17'd9574,17'd9574,17'd9703,17'd9703,17'd9704,17'd9704,17'd9704,17'd9575,17'd8371,17'd8371,17'd8066,17'd4767,17'd5090,17'd5255,17'd6626,17'd6140,17'd6140,17'd6305,17'd6138,17'd6138,17'd6304,17'd6304,17'd9985,17'd9842,17'd9986,17'd9987,17'd9843,17'd9843,17'd9844,17'd9844,17'd9845,17'd9988,17'd9989,17'd9990,17'd9991,17'd9992,17'd9850,17'd9584,17'd9585,17'd9312,17'd9166,17'd9314,17'd9588,17'd9993,17'd9852,17'd9450,17'd9994,17'd9995,17'd9996,17'd9997,17'd9998,17'd9999,17'd10000,17'd10001,17'd10002,17'd10003,17'd10004,17'd10005,17'd10006,17'd10007,17'd10008,17'd9868,17'd10009,17'd10009,17'd10010,17'd9868,17'd10011,17'd10012,17'd9731,17'd9615,17'd9872,17'd9735,17'd9874,17'd10013,17'd10013,17'd10014,17'd10014,17'd10015,17'd10016,17'd10017,17'd10018,17'd9879,17'd10019,17'd10020,17'd10021,17'd10022,17'd10023,17'd9883,17'd9884,17'd10024,17'd9742,17'd10025,17'd10026,17'd10026,17'd9339,17'd9339,17'd9189,17'd9041,17'd8884,17'd10027,17'd9886,17'd9887,17'd10028,17'd8255,17'd10029,17'd7622,17'd10030,17'd10031,17'd10032,17'd10033,17'd10034,17'd8593,17'd10035,17'd9898,17'd10036,17'd10037,17'd8279,17'd9359,17'd8444,17'd6529,17'd8132,17'd719,17'd1197,17'd133,17'd1481,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd133,17'd133,17'd131,17'd5467,17'd3031,17'd10038,17'd10039,17'd10040,17'd10041,17'd6540,17'd8288,17'd7658,17'd9216,17'd10042,17'd10043,17'd10044,17'd10045,17'd10046,17'd7496,17'd7497,17'd7835,17'd9221,17'd10047,17'd9641,17'd10048,17'd10049,17'd10050,17'd9915,17'd9377,17'd9510,17'd10051,17'd10052,17'd9920,17'd10053,17'd10054,17'd10055,17'd10056,17'd10057,17'd9925,17'd9926,17'd10058,17'd10059,17'd8925,17'd9233,17'd9232,17'd10060,17'd10061,17'd10062,17'd10063,17'd9780,17'd10064,17'd10064,17'd10064,17'd10064,17'd9651,17'd9781,17'd9779,17'd9085,17'd9655,17'd9086,17'd9237,17'd9392,17'd9393,17'd7665,17'd7666,17'd7175,17'd7175,17'd6848,17'd8146,17'd8147,17'd9930,17'd9930,17'd7329,17'd9522,17'd7329,17'd7329,17'd6550,17'd6550,17'd7176,17'd7176,17'd8932,17'd7999,17'd8629,17'd9931,17'd9931,17'd9090,17'd8304,17'd7668,17'd8780,17'd9933,17'd9933,17'd9934,17'd9934,17'd9934,17'd7500,17'd7011,17'd8631,17'd8305,17'd9396,17'd10065,17'd7185,17'd8940,17'd8785,17'd9526,17'd4857,17'd10066,17'd10067,17'd10068,17'd10069,17'd10070,17'd10071,17'd10072,17'd447,17'd1679,17'd10073,17'd3586,17'd9104,17'd10074,17'd10075,17'd3412,17'd5368,17'd3726,17'd3577,17'd7348,17'd7347,17'd7029,17'd8169,17'd8170,17'd8795,17'd10076,17'd9534,17'd8954,17'd8955,17'd10077,17'd9947,17'd10078,17'd9256,17'd9538,17'd9408,17'd8495,17'd8495,17'd7517,17'd7347,17'd7195,17'd7860,17'd7195,17'd9108,17'd8323,17'd8648,17'd10079,17'd8962,17'd8807,17'd8963,17'd7864,17'd9542,17'd9412,17'd9412,17'd8500,17'd9119,17'd9119,17'd9119,17'd9119,17'd8809,17'd8809,17'd8809,17'd7867,17'd9799,17'd7698,17'd8181,17'd10080,17'd8810,17'd10081,17'd10082,17'd10083,17'd8187,17'd7705,17'd7705,17'd7537,17'd7537,17'd7705,17'd6890,17'd6094,17'd6581,17'd6581,17'd6416,17'd6416,17'd6416,17'd6581,17'd4728,17'd4085,17'd2905,17'd4084,17'd970,17'd425,17'd1966,17'd952,17'd2116,17'd9671
},
'{
17'd6262,17'd6262,17'd5198,17'd5053,17'd4087,17'd4428,17'd6584,17'd7711,17'd1689,17'd14,17'd14,17'd15,17'd0,17'd0,17'd0,17'd2,17'd2,17'd466,17'd4247,17'd1689,17'd2781,17'd2592,17'd2422,17'd3250,17'd1831,17'd466,17'd12,17'd2933,17'd23,17'd6,17'd5205,17'd5205,17'd8340,17'd8340,17'd8340,17'd8340,17'd5205,17'd6,17'd9263,17'd6097,17'd7713,17'd6596,17'd8511,17'd10084,17'd7054,17'd7052,17'd8515,17'd9964,17'd10085,17'd8664,17'd8977,17'd10086,17'd7717,17'd10087,17'd9269,17'd8666,17'd6269,17'd9551,17'd8984,17'd8341,17'd10088,17'd7056,17'd6742,17'd7885,17'd9966,17'd10089,17'd10090,17'd10091,17'd10092,17'd10092,17'd2936,17'd9969,17'd654,17'd31,17'd3255,17'd3255,17'd3595,17'd3907,17'd6598,17'd10093,17'd6437,17'd7225,17'd7556,17'd7556,17'd6904,17'd9970,17'd7064,17'd6907,17'd7064,17'd7064,17'd6602,17'd7065,17'd7229,17'd7067,17'd7068,17'd7069,17'd9280,17'd9143,17'd8831,17'd9820,17'd10094,17'd10095,17'd10096,17'd10097,17'd10098,17'd10099,17'd10100,17'd8838,17'd10101,17'd10102,17'd10103,17'd10104,17'd10105,17'd10106,17'd10107,17'd10108,17'd10108,17'd10109,17'd10110,17'd10110,17'd9841,17'd9568,17'd9841,17'd9572,17'd9437,17'd8064,17'd10111,17'd10112,17'd9574,17'd9300,17'd9300,17'd9300,17'd9300,17'd9703,17'd9703,17'd9703,17'd10113,17'd10113,17'd9007,17'd8538,17'd7750,17'd7750,17'd5255,17'd5255,17'd9303,17'd6139,17'd6139,17'd5252,17'd9009,17'd9009,17'd9008,17'd10114,17'd10115,17'd10116,17'd10117,17'd10118,17'd10119,17'd10120,17'd10121,17'd9988,17'd9988,17'd9989,17'd10122,17'd10123,17'd10124,17'd10125,17'd10126,17'd9446,17'd10127,17'd9166,17'd10128,17'd10129,17'd9170,17'd9317,17'd10130,17'd9712,17'd10131,17'd10132,17'd10133,17'd10134,17'd10135,17'd10136,17'd10137,17'd10138,17'd10139,17'd10140,17'd10141,17'd10142,17'd10143,17'd10144,17'd10145,17'd10146,17'd10147,17'd10148,17'd10149,17'd10150,17'd10151,17'd9872,17'd9734,17'd9873,17'd9878,17'd10152,17'd10015,17'd10153,17'd10154,17'd10155,17'd10155,17'd10156,17'd10157,17'd10158,17'd10159,17'd10160,17'd10161,17'd10162,17'd10163,17'd10164,17'd10165,17'd10166,17'd10167,17'd10168,17'd10169,17'd10170,17'd10171,17'd10172,17'd10026,17'd10173,17'd10174,17'd10175,17'd10176,17'd8884,17'd10177,17'd10178,17'd8252,17'd10179,17'd10180,17'd10181,17'd8892,17'd10182,17'd7469,17'd10183,17'd10184,17'd10185,17'd10186,17'd10187,17'd10188,17'd10189,17'd8279,17'd8130,17'd7647,17'd6529,17'd6198,17'd541,17'd356,17'd356,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd1197,17'd133,17'd134,17'd132,17'd3168,17'd10190,17'd10191,17'd10192,17'd9497,17'd10193,17'd10194,17'd10195,17'd6380,17'd8143,17'd10196,17'd10197,17'd10198,17'd10199,17'd10046,17'd10200,17'd7496,17'd9766,17'd9221,17'd10201,17'd10202,17'd10203,17'd10204,17'd9507,17'd9375,17'd10205,17'd10206,17'd10207,17'd10208,17'd10209,17'd10210,17'd9923,17'd10055,17'd10056,17'd10211,17'd10212,17'd10213,17'd10214,17'd10215,17'd10215,17'd10216,17'd10217,17'd8928,17'd10218,17'd10219,17'd10220,17'd10221,17'd10222,17'd10223,17'd10224,17'd10225,17'd10226,17'd10227,17'd9385,17'd9652,17'd10228,17'd10229,17'd9389,17'd10230,17'd10231,17'd10232,17'd10233,17'd10234,17'd10235,17'd10234,17'd10235,17'd7010,17'd7329,17'd7329,17'd7329,17'd7329,17'd7329,17'd8146,17'd8146,17'd7169,17'd7169,17'd6386,17'd6217,17'd6850,17'd7176,17'd8779,17'd7999,17'd10236,17'd10237,17'd8154,17'd8154,17'd9090,17'd8780,17'd8780,17'd7499,17'd10238,17'd9934,17'd8001,17'd6557,17'd6559,17'd8156,17'd8157,17'd9396,17'd10239,17'd9240,17'd8160,17'd10240,17'd10241,17'd10066,17'd10242,17'd10243,17'd10244,17'd10245,17'd10246,17'd10247,17'd4228,17'd627,17'd1240,17'd10073,17'd3586,17'd3585,17'd3239,17'd9532,17'd3888,17'd5369,17'd4411,17'd9108,17'd9250,17'd8490,17'd10248,17'd7858,17'd8020,17'd9405,17'd10076,17'd9405,17'd9405,17'd9946,17'd9254,17'd9794,17'd10249,17'd9256,17'd9538,17'd9408,17'd9115,17'd8495,17'd7347,17'd7348,17'd6873,17'd7348,17'd7348,17'd9250,17'd9540,17'd8801,17'd10250,17'd10250,17'd10251,17'd8959,17'd7864,17'd8178,17'd7523,17'd9412,17'd9119,17'd10252,17'd10253,17'd10254,17'd9119,17'd7867,17'd9798,17'd10255,17'd8028,17'd7867,17'd8809,17'd8181,17'd10256,17'd8655,17'd9802,17'd10082,17'd10257,17'd7878,17'd7537,17'd9124,17'd9261,17'd7537,17'd8187,17'd10258,17'd6416,17'd6416,17'd6416,17'd8187,17'd6889,17'd3073,17'd4728,17'd4422,17'd5192,17'd4084,17'd1823,17'd425,17'd205,17'd424,17'd2116,17'd10259
},
'{
17'd6262,17'd5198,17'd5053,17'd5200,17'd4244,17'd4733,17'd7545,17'd4886,17'd1127,17'd14,17'd15,17'd15,17'd0,17'd0,17'd0,17'd2,17'd13,17'd466,17'd1127,17'd1689,17'd2781,17'd2784,17'd2422,17'd1688,17'd4247,17'd13,17'd806,17'd10260,17'd5,17'd6,17'd5205,17'd5205,17'd8190,17'd8340,17'd8340,17'd8340,17'd8040,17'd5205,17'd8196,17'd6098,17'd6435,17'd6106,17'd9551,17'd10261,17'd7221,17'd6895,17'd7219,17'd7716,17'd10085,17'd8976,17'd9128,17'd10262,17'd7548,17'd9269,17'd8667,17'd6431,17'd9551,17'd10263,17'd8983,17'd10264,17'd8342,17'd8982,17'd6431,17'd7714,17'd9420,17'd10265,17'd10266,17'd10267,17'd10267,17'd10092,17'd10268,17'd10268,17'd31,17'd31,17'd3255,17'd3255,17'd3755,17'd3907,17'd10269,17'd10093,17'd6903,17'd7225,17'd7556,17'd9970,17'd9970,17'd9817,17'd7228,17'd9277,17'd7228,17'd6602,17'd7065,17'd7066,17'd7067,17'd7068,17'd10270,17'd6910,17'd10271,17'd8203,17'd8526,17'd9821,17'd10272,17'd10273,17'd10274,17'd10098,17'd9561,17'd10275,17'd8359,17'd9830,17'd9979,17'd10276,17'd10277,17'd10278,17'd10279,17'd10280,17'd10110,17'd10110,17'd10109,17'd10109,17'd10281,17'd10281,17'd9841,17'd9568,17'd10282,17'd10283,17'd10284,17'd10111,17'd10285,17'd10286,17'd9574,17'd9300,17'd9300,17'd9300,17'd9703,17'd9703,17'd9703,17'd9703,17'd10113,17'd9703,17'd9007,17'd8538,17'd7750,17'd5409,17'd5255,17'd5689,17'd6139,17'd6138,17'd6138,17'd6138,17'd9009,17'd9008,17'd10114,17'd10114,17'd10116,17'd10117,17'd8685,17'd10287,17'd10119,17'd10120,17'd9988,17'd9988,17'd9989,17'd10288,17'd10289,17'd10123,17'd10290,17'd10291,17'd10292,17'd9708,17'd9313,17'd10293,17'd10294,17'd10295,17'd9317,17'd9450,17'd10296,17'd9854,17'd10297,17'd10298,17'd9997,17'd10299,17'd10300,17'd10301,17'd10302,17'd10303,17'd10304,17'd10305,17'd10306,17'd10307,17'd10007,17'd10308,17'd10309,17'd10310,17'd10146,17'd10148,17'd10311,17'd10312,17'd10313,17'd10314,17'd10315,17'd9878,17'd10016,17'd10153,17'd10316,17'd10317,17'd10317,17'd10318,17'd10318,17'd10319,17'd10320,17'd10321,17'd10322,17'd10323,17'd10324,17'd10325,17'd10326,17'd10165,17'd10327,17'd10328,17'd10328,17'd10329,17'd10330,17'd10331,17'd10332,17'd10333,17'd10334,17'd10173,17'd10335,17'd10336,17'd10175,17'd10337,17'd10338,17'd10339,17'd10340,17'd7953,17'd10341,17'd10342,17'd10343,17'd10344,17'd10345,17'd10346,17'd10347,17'd10034,17'd10348,17'd10349,17'd10350,17'd9631,17'd8750,17'd10351,17'd9359,17'd9360,17'd1044,17'd541,17'd356,17'd1481,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd131,17'd132,17'd132,17'd133,17'd133,17'd542,17'd542,17'd134,17'd131,17'd2861,17'd10352,17'd10353,17'd10354,17'd10355,17'd10356,17'd10357,17'd10358,17'd7006,17'd10196,17'd10359,17'd10359,17'd10360,17'd10361,17'd8609,17'd9372,17'd10362,17'd7835,17'd10363,17'd8762,17'd10203,17'd10364,17'd10049,17'd9643,17'd10365,17'd10366,17'd9918,17'd9770,17'd10367,17'd10368,17'd10210,17'd10369,17'd10370,17'd10371,17'd10372,17'd10373,17'd10374,17'd10214,17'd10215,17'd10215,17'd8928,17'd10217,17'd10375,17'd10375,17'd9928,17'd10376,17'd10223,17'd10222,17'd10222,17'd10223,17'd10377,17'd10225,17'd10226,17'd9384,17'd9780,17'd9517,17'd9652,17'd10228,17'd9519,17'd9389,17'd10378,17'd10232,17'd10233,17'd10233,17'd10233,17'd10233,17'd7010,17'd9522,17'd6849,17'd6849,17'd7329,17'd7329,17'd8147,17'd8147,17'd7169,17'd7169,17'd6550,17'd6386,17'd6850,17'd6850,17'd8932,17'd10379,17'd8000,17'd10236,17'd9394,17'd9090,17'd8154,17'd9394,17'd8780,17'd8780,17'd9933,17'd10380,17'd8001,17'd8001,17'd6559,17'd7501,17'd8156,17'd8157,17'd10381,17'd10239,17'd8004,17'd10382,17'd10240,17'd10383,17'd10384,17'd10242,17'd10243,17'd10385,17'd10386,17'd10387,17'd10388,17'd4398,17'd623,17'd1678,17'd3097,17'd3096,17'd8642,17'd10389,17'd3238,17'd4076,17'd6874,17'd4412,17'd10390,17'd8803,17'd7687,17'd7687,17'd8020,17'd7857,17'd10076,17'd9405,17'd9405,17'd9405,17'd10391,17'd9536,17'd9947,17'd10249,17'd9949,17'd9113,17'd9408,17'd8495,17'd7347,17'd7347,17'd6873,17'd6873,17'd7348,17'd7347,17'd9409,17'd8648,17'd10250,17'd10250,17'd10250,17'd8959,17'd8650,17'd7350,17'd9542,17'd9542,17'd7867,17'd8653,17'd10253,17'd10392,17'd9119,17'd10252,17'd8500,17'd10255,17'd7867,17'd7867,17'd8809,17'd8809,17'd9799,17'd9120,17'd7876,17'd10393,17'd10394,17'd10395,17'd7705,17'd9124,17'd9261,17'd7537,17'd8187,17'd10258,17'd6416,17'd6416,17'd8187,17'd8187,17'd6889,17'd3073,17'd4728,17'd4728,17'd4422,17'd3742,17'd1667,17'd1396,17'd775,17'd1272,17'd422,17'd10396
},
'{
17'd10397,17'd5198,17'd5200,17'd10398,17'd4245,17'd4887,17'd3250,17'd1689,17'd14,17'd14,17'd0,17'd1,17'd1,17'd0,17'd0,17'd2,17'd466,17'd466,17'd1127,17'd1689,17'd3250,17'd2422,17'd1831,17'd1127,17'd2,17'd806,17'd2591,17'd2421,17'd6,17'd5205,17'd8190,17'd8190,17'd8190,17'd8190,17'd8340,17'd8339,17'd8338,17'd8190,17'd9961,17'd6588,17'd6434,17'd9415,17'd10399,17'd7715,17'd6738,17'd7549,17'd9264,17'd7220,17'd8818,17'd9128,17'd10400,17'd9548,17'd9418,17'd8980,17'd7055,17'd10401,17'd10263,17'd9551,17'd10402,17'd10403,17'd10399,17'd7055,17'd7714,17'd6271,17'd10404,17'd10405,17'd10268,17'd10268,17'd10406,17'd10407,17'd3752,17'd3429,17'd982,17'd469,17'd3254,17'd3255,17'd3755,17'd3907,17'd6598,17'd10093,17'd9555,17'd7556,17'd10408,17'd10409,17'd7392,17'd6282,17'd6282,17'd7065,17'd7065,17'd5979,17'd5979,17'd7066,17'd10410,17'd9818,17'd10270,17'd10411,17'd6911,17'd9558,17'd10412,17'd9688,17'd10413,17'd10414,17'd10415,17'd10416,17'd10417,17'd10418,17'd10419,17'd8681,17'd10420,17'd10421,17'd10422,17'd10423,17'd10424,17'd10425,17'd10109,17'd10109,17'd10109,17'd10109,17'd9568,17'd9841,17'd9841,17'd9568,17'd10426,17'd8064,17'd10285,17'd10427,17'd10286,17'd10286,17'd9574,17'd9574,17'd10428,17'd10428,17'd10429,17'd10429,17'd9703,17'd9703,17'd9703,17'd9703,17'd10430,17'd7750,17'd5255,17'd5689,17'd5689,17'd5689,17'd6139,17'd6139,17'd6138,17'd6304,17'd9008,17'd9842,17'd9986,17'd10431,17'd10432,17'd10432,17'd8844,17'd10119,17'd9844,17'd9844,17'd9988,17'd9989,17'd10122,17'd10122,17'd10433,17'd10434,17'd10291,17'd10126,17'd10292,17'd9708,17'd9447,17'd10129,17'd9169,17'd10435,17'd9710,17'd10436,17'd10437,17'd10438,17'd10439,17'd10440,17'd10441,17'd10442,17'd10443,17'd10444,17'd10445,17'd10446,17'd10447,17'd10448,17'd10449,17'd10450,17'd10451,17'd10452,17'd10453,17'd10454,17'd10455,17'd10456,17'd10457,17'd10458,17'd10459,17'd10460,17'd10461,17'd10462,17'd10463,17'd10155,17'd10464,17'd10464,17'd10465,17'd10465,17'd10156,17'd10466,17'd10467,17'd10468,17'd10323,17'd10469,17'd10470,17'd10471,17'd10472,17'd10472,17'd10473,17'd10474,17'd10475,17'd10476,17'd10477,17'd10478,17'd10479,17'd9884,17'd9479,17'd9345,17'd9346,17'd9743,17'd9743,17'd10175,17'd8879,17'd9744,17'd8101,17'd10480,17'd8424,17'd10481,17'd10482,17'd10483,17'd10484,17'd10485,17'd10486,17'd8592,17'd10487,17'd10488,17'd10489,17'd10490,17'd10037,17'd10491,17'd7978,17'd7812,17'd6529,17'd719,17'd356,17'd1481,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd542,17'd133,17'd132,17'd357,17'd10492,17'd10493,17'd10494,17'd8905,17'd10495,17'd10496,17'd10497,17'd10498,17'd8911,17'd8608,17'd10359,17'd10359,17'd10499,17'd10500,17'd8759,17'd9069,17'd10362,17'd10501,17'd9640,17'd9767,17'd10204,17'd10049,17'd10049,17'd9643,17'd10365,17'd10366,17'd9644,17'd10502,17'd10503,17'd10367,17'd10504,17'd10210,17'd9923,17'd10056,17'd10505,17'd10506,17'd10374,17'd10215,17'd10507,17'd10507,17'd8928,17'd8928,17'd10508,17'd10509,17'd10508,17'd10064,17'd9517,17'd10063,17'd10221,17'd10221,17'd10063,17'd9517,17'd10377,17'd10510,17'd10227,17'd10226,17'd9518,17'd9652,17'd9653,17'd9388,17'd9389,17'd10511,17'd10232,17'd10232,17'd10232,17'd10232,17'd10233,17'd10235,17'd6849,17'd6849,17'd6849,17'd7329,17'd8146,17'd8146,17'd8146,17'd6848,17'd6550,17'd6550,17'd6216,17'd6217,17'd10512,17'd10512,17'd8000,17'd8000,17'd9394,17'd9090,17'd8154,17'd8154,17'd10513,17'd10514,17'd10515,17'd10516,17'd10517,17'd8001,17'd6709,17'd6710,17'd6711,17'd6712,17'd8157,17'd10518,17'd8635,17'd8004,17'd10382,17'd10240,17'd9242,17'd10519,17'd10520,17'd10521,17'd10245,17'd10522,17'd10523,17'd10524,17'd4398,17'd626,17'd10525,17'd2930,17'd3089,17'd3239,17'd3584,17'd3888,17'd5504,17'd3883,17'd7861,17'd9250,17'd8490,17'd7687,17'd7858,17'd8020,17'd9405,17'd10076,17'd9405,17'd8172,17'd8798,17'd10526,17'd9255,17'd10527,17'd9256,17'd9538,17'd9407,17'd9408,17'd8174,17'd7347,17'd8490,17'd7688,17'd7348,17'd7347,17'd9108,17'd8496,17'd10528,17'd10528,17'd10250,17'd9410,17'd8962,17'd7690,17'd9542,17'd8652,17'd10529,17'd8653,17'd10253,17'd10253,17'd10252,17'd10252,17'd7867,17'd8326,17'd8326,17'd7867,17'd8809,17'd8809,17'd9799,17'd10256,17'd8810,17'd10081,17'd10530,17'd10531,17'd7705,17'd7705,17'd9261,17'd7705,17'd8187,17'd8187,17'd6416,17'd8187,17'd8187,17'd8187,17'd4559,17'd6889,17'd7211,17'd4728,17'd4422,17'd1810,17'd1667,17'd605,17'd204,17'd1244,17'd1527,17'd10396
},
'{
17'd10532,17'd5053,17'd10533,17'd10534,17'd4887,17'd7711,17'd1689,17'd1127,17'd14,17'd15,17'd0,17'd1,17'd1,17'd0,17'd2,17'd2,17'd1127,17'd1127,17'd1689,17'd1689,17'd2422,17'd10535,17'd1688,17'd14,17'd12,17'd1275,17'd2421,17'd7215,17'd3753,17'd5205,17'd8190,17'd8190,17'd10536,17'd8190,17'd8040,17'd8338,17'd8338,17'd10537,17'd10538,17'd6435,17'd6104,17'd7546,17'd8666,17'd7221,17'd6895,17'd7550,17'd7377,17'd7220,17'd9678,17'd10539,17'd8819,17'd10540,17'd9549,17'd6898,17'd10401,17'd10541,17'd10542,17'd6103,17'd6734,17'd9962,17'd9416,17'd8822,17'd6741,17'd7056,17'd10543,17'd10544,17'd3429,17'd10268,17'd10545,17'd10546,17'd3429,17'd10547,17'd2259,17'd982,17'd3254,17'd3255,17'd3755,17'd9554,17'd6598,17'd6903,17'd7556,17'd7556,17'd10408,17'd7730,17'd6282,17'd6282,17'd7393,17'd10548,17'd10548,17'd5814,17'd5814,17'd10410,17'd9818,17'd10270,17'd6752,17'd8990,17'd8526,17'd10549,17'd10550,17'd9824,17'd10551,17'd10415,17'd10552,17'd10553,17'd10418,17'd10554,17'd10555,17'd10556,17'd10557,17'd10558,17'd10559,17'd10560,17'd10561,17'd10425,17'd10109,17'd10109,17'd10109,17'd10281,17'd9841,17'd9841,17'd9841,17'd9571,17'd8064,17'd10562,17'd10427,17'd10563,17'd10112,17'd10564,17'd9574,17'd9574,17'd10428,17'd10428,17'd10565,17'd10429,17'd9703,17'd9703,17'd9703,17'd8538,17'd7750,17'd5409,17'd5689,17'd5689,17'd5689,17'd5689,17'd5253,17'd6139,17'd6138,17'd6304,17'd9842,17'd9842,17'd9441,17'd10116,17'd7581,17'd10432,17'd10119,17'd10119,17'd9844,17'd10566,17'd9989,17'd10567,17'd10568,17'd10569,17'd10434,17'd10291,17'd10570,17'd9585,17'd9586,17'd10571,17'd10293,17'd9020,17'd10435,17'd9319,17'd9451,17'd10572,17'd10438,17'd10573,17'd10574,17'd10575,17'd10576,17'd10577,17'd10578,17'd10579,17'd10580,17'd10581,17'd10582,17'd10583,17'd10584,17'd10585,17'd10586,17'd10587,17'd10588,17'd10589,17'd10590,17'd10591,17'd10592,17'd10152,17'd10016,17'd10462,17'd10463,17'd10156,17'd10465,17'd10465,17'd10465,17'd10465,17'd10593,17'd10594,17'd10595,17'd10596,17'd10597,17'd10468,17'd10598,17'd10599,17'd10600,17'd10601,17'd10602,17'd10603,17'd10604,17'd10604,17'd10604,17'd10604,17'd10605,17'd10477,17'd10606,17'd10479,17'd9885,17'd9480,17'd9620,17'd9346,17'd9339,17'd9190,17'd9045,17'd10607,17'd10608,17'd7785,17'd10609,17'd10610,17'd10611,17'd10612,17'd7633,17'd10346,17'd10613,17'd10614,17'd10615,17'd10616,17'd10617,17'd10618,17'd10619,17'd10620,17'd10621,17'd9359,17'd6529,17'd3025,17'd134,17'd134,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd132,17'd131,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd357,17'd9060,17'd10622,17'd10623,17'd10624,17'd10495,17'd10625,17'd10626,17'd9764,17'd6543,17'd9503,17'd10627,17'd10628,17'd10499,17'd8454,17'd9372,17'd10362,17'd7828,17'd10629,17'd10630,17'd10631,17'd10632,17'd10633,17'd10633,17'd9643,17'd10365,17'd10366,17'd9644,17'd9645,17'd10634,17'd10208,17'd10635,17'd10209,17'd9923,17'd10057,17'd10636,17'd10637,17'd8925,17'd10638,17'd10639,17'd10640,17'd10217,17'd10217,17'd10508,17'd10509,17'd10509,17'd10508,17'd9384,17'd9780,17'd9517,17'd10063,17'd10063,17'd10063,17'd10377,17'd10225,17'd10226,17'd10227,17'd10226,17'd9518,17'd9652,17'd9653,17'd9388,17'd9389,17'd10511,17'd10232,17'd10232,17'd10231,17'd10378,17'd10378,17'd7010,17'd6849,17'd7329,17'd7329,17'd6848,17'd6848,17'd8146,17'd8146,17'd7168,17'd7168,17'd6550,17'd6217,17'd10512,17'd10512,17'd8000,17'd7999,17'd9394,17'd9394,17'd9090,17'd8154,17'd9657,17'd10641,17'd10642,17'd10515,17'd10516,17'd10517,17'd6557,17'd6559,17'd7501,17'd6711,17'd8156,17'd7331,17'd7017,17'd8308,17'd9935,17'd10643,17'd10644,17'd10645,17'd10646,17'd10243,17'd9939,17'd10647,17'd10648,17'd10649,17'd5495,17'd4398,17'd3072,17'd10525,17'd4241,17'd3089,17'd9532,17'd3238,17'd3887,17'd5505,17'd3408,17'd9108,17'd8490,17'd7687,17'd7858,17'd7858,17'd8019,17'd10076,17'd10076,17'd8019,17'd8955,17'd10526,17'd10650,17'd9110,17'd10249,17'd9949,17'd9538,17'd9539,17'd8495,17'd7347,17'd8490,17'd8490,17'd7347,17'd7347,17'd9108,17'd8496,17'd9115,17'd10528,17'd8801,17'd8801,17'd9541,17'd8650,17'd9411,17'd9411,17'd8027,17'd10651,17'd10652,17'd10652,17'd10252,17'd9119,17'd8809,17'd7867,17'd9259,17'd8809,17'd8809,17'd7867,17'd9955,17'd10653,17'd10654,17'd8656,17'd10655,17'd10394,17'd9414,17'd7705,17'd7705,17'd7705,17'd8187,17'd8187,17'd6416,17'd8187,17'd8187,17'd8187,17'd5183,17'd6889,17'd4882,17'd4728,17'd4422,17'd1810,17'd1667,17'd1394,17'd424,17'd202,17'd1527,17'd10396
},
'{
17'd4734,17'd4426,17'd4428,17'd6584,17'd3250,17'd1689,17'd1127,17'd2,17'd2,17'd0,17'd1,17'd1,17'd1,17'd0,17'd2,17'd14,17'd1689,17'd1689,17'd2781,17'd3250,17'd1831,17'd1831,17'd1127,17'd0,17'd806,17'd2591,17'd8,17'd6,17'd3753,17'd5205,17'd10656,17'd7884,17'd10536,17'd7374,17'd8338,17'd10657,17'd8339,17'd10658,17'd10659,17'd8518,17'd9680,17'd7889,17'd7550,17'd7053,17'd8974,17'd8974,17'd10660,17'd9548,17'd10262,17'd8665,17'd7719,17'd8980,17'd8666,17'd7714,17'd9133,17'd10661,17'd9137,17'd10662,17'd10663,17'd10664,17'd10665,17'd7722,17'd10666,17'd10667,17'd10668,17'd2781,17'd10545,17'd10407,17'd3593,17'd10669,17'd10669,17'd10670,17'd10671,17'd2259,17'd3254,17'd3754,17'd6278,17'd5971,17'd6437,17'd6903,17'd6904,17'd6904,17'd10672,17'd10672,17'd10673,17'd10674,17'd5814,17'd5813,17'd5813,17'd5386,17'd9818,17'd10270,17'd6910,17'd9686,17'd8990,17'd9557,17'd10675,17'd9974,17'd10676,17'd9826,17'd10677,17'd10678,17'd10679,17'd10680,17'd10554,17'd10681,17'd10682,17'd10683,17'd10684,17'd10685,17'd10686,17'd10687,17'd10688,17'd10689,17'd10109,17'd10281,17'd10281,17'd10281,17'd9841,17'd9841,17'd9571,17'd10690,17'd10111,17'd10691,17'd10286,17'd10564,17'd10692,17'd10692,17'd10428,17'd10428,17'd10428,17'd10693,17'd10428,17'd10428,17'd10694,17'd9159,17'd10430,17'd7750,17'd5409,17'd5689,17'd6140,17'd6140,17'd6305,17'd6305,17'd5253,17'd6139,17'd10695,17'd10114,17'd9986,17'd9441,17'd9987,17'd9987,17'd10696,17'd8844,17'd10697,17'd9844,17'd10566,17'd10698,17'd10288,17'd10122,17'd10699,17'd10700,17'd9444,17'd9311,17'd9446,17'd10701,17'd9708,17'd9447,17'd8856,17'd10702,17'd9319,17'd10703,17'd9592,17'd9854,17'd10704,17'd10705,17'd10575,17'd10706,17'd10707,17'd10708,17'd10709,17'd10710,17'd10711,17'd10712,17'd10713,17'd10714,17'd10715,17'd10716,17'd10717,17'd10718,17'd10719,17'd10720,17'd10721,17'd10722,17'd10723,17'd10724,17'd10155,17'd10725,17'd10726,17'd10726,17'd10726,17'd10725,17'd10155,17'd10463,17'd10595,17'd10727,17'd10728,17'd10159,17'd10729,17'd10730,17'd10468,17'd10731,17'd10323,17'd10732,17'd10733,17'd10734,17'd10735,17'd10736,17'd10737,17'd10738,17'd10739,17'd10740,17'd10325,17'd10741,17'd9473,17'd10742,17'd10743,17'd9341,17'd10744,17'd9191,17'd8720,17'd8723,17'd8416,17'd10745,17'd10746,17'd10747,17'd10748,17'd10749,17'd10750,17'd10751,17'd10752,17'd10753,17'd10754,17'd10616,17'd10755,17'd10756,17'd9631,17'd10757,17'd10758,17'd10351,17'd8131,17'd8132,17'd1197,17'd134,17'd1045,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd131,17'd357,17'd10759,17'd10760,17'd10761,17'd10762,17'd10763,17'd10764,17'd10765,17'd6542,17'd7658,17'd9503,17'd10627,17'd10766,17'd10499,17'd8759,17'd7496,17'd7497,17'd7828,17'd10629,17'd10630,17'd10767,17'd10768,17'd10633,17'd9643,17'd10769,17'd9508,17'd9508,17'd9644,17'd9644,17'd9645,17'd9770,17'd8921,17'd10770,17'd9922,17'd10771,17'd10772,17'd10059,17'd8925,17'd10217,17'd10640,17'd10509,17'd10508,17'd10064,17'd10064,17'd10508,17'd10508,17'd10508,17'd10508,17'd10508,17'd10064,17'd9928,17'd10376,17'd10219,17'd10224,17'd10224,17'd10225,17'd10226,17'd10227,17'd10773,17'd9518,17'd9781,17'd10774,17'd9388,17'd9519,17'd10230,17'd10775,17'd10776,17'd10511,17'd10230,17'd10231,17'd10233,17'd6849,17'd7329,17'd7329,17'd7329,17'd8146,17'd8147,17'd7329,17'd7168,17'd6550,17'd6386,17'd10512,17'd10512,17'd6850,17'd6704,17'd6707,17'd10237,17'd9394,17'd8154,17'd8304,17'd10777,17'd10642,17'd10642,17'd10778,17'd10779,17'd8001,17'd7836,17'd6559,17'd7501,17'd7501,17'd6561,17'd6713,17'd10780,17'd10781,17'd10782,17'd10783,17'd10784,17'd10645,17'd10785,17'd10786,17'd10787,17'd10788,17'd10789,17'd10790,17'd5936,17'd2558,17'd1945,17'd2585,17'd3894,17'd3414,17'd9533,17'd3888,17'd5041,17'd3405,17'd3578,17'd8490,17'd7687,17'd7686,17'd7686,17'd7856,17'd9405,17'd10076,17'd10076,17'd9405,17'd9946,17'd9254,17'd9110,17'd10078,17'd9256,17'd9949,17'd9538,17'd8495,17'd8495,17'd7347,17'd7347,17'd7347,17'd7347,17'd7347,17'd8022,17'd9115,17'd9115,17'd9407,17'd9407,17'd9541,17'd8962,17'd7691,17'd8499,17'd10791,17'd10529,17'd8653,17'd8653,17'd8653,17'd9119,17'd8028,17'd7867,17'd8326,17'd8809,17'd7867,17'd7867,17'd8809,17'd10653,17'd10792,17'd8655,17'd10793,17'd10082,17'd10794,17'd9544,17'd7705,17'd7705,17'd7705,17'd7537,17'd8507,17'd7537,17'd7537,17'd8187,17'd4714,17'd3073,17'd5940,17'd6415,17'd2905,17'd6407,17'd604,17'd781,17'd424,17'd1382,17'd1528,17'd195
},
'{
17'd4891,17'd4244,17'd4733,17'd4577,17'd1689,17'd1127,17'd2,17'd2,17'd0,17'd0,17'd0,17'd1,17'd0,17'd0,17'd2,17'd1127,17'd1689,17'd3250,17'd3250,17'd3250,17'd1688,17'd4247,17'd2,17'd3,17'd2933,17'd2421,17'd6,17'd6,17'd5205,17'd5205,17'd10656,17'd7884,17'd7374,17'd7374,17'd8339,17'd8339,17'd10795,17'd10796,17'd9135,17'd6595,17'd6897,17'd7550,17'd7219,17'd7219,17'd9548,17'd8979,17'd8979,17'd10262,17'd10797,17'd10798,17'd9418,17'd8345,17'd10799,17'd10401,17'd10661,17'd10800,17'd6106,17'd9272,17'd7546,17'd7890,17'd7051,17'd7546,17'd8983,17'd10801,17'd2781,17'd3750,17'd10407,17'd10545,17'd10669,17'd10802,17'd10802,17'd10802,17'd32,17'd982,17'd3255,17'd3754,17'd6278,17'd6598,17'd6903,17'd6903,17'd6904,17'd6904,17'd10672,17'd6112,17'd10548,17'd10548,17'd5223,17'd5386,17'd5386,17'd6751,17'd9971,17'd9280,17'd8831,17'd9557,17'd8526,17'd9821,17'd10095,17'd10803,17'd10804,17'd9287,17'd10417,17'd10805,17'd10806,17'd10807,17'd9429,17'd10682,17'd10808,17'd10809,17'd10685,17'd10810,17'd10687,17'd10811,17'd10812,17'd10689,17'd10281,17'd10281,17'd10813,17'd10814,17'd9841,17'd9571,17'd10283,17'd10815,17'd10427,17'd10816,17'd10817,17'd10564,17'd10692,17'd10692,17'd10428,17'd10428,17'd10428,17'd10428,17'd10428,17'd9574,17'd9159,17'd9159,17'd7750,17'd5409,17'd5255,17'd5689,17'd6140,17'd6140,17'd6305,17'd6305,17'd6139,17'd6139,17'd10695,17'd10114,17'd9986,17'd9441,17'd9987,17'd10432,17'd8844,17'd10119,17'd9844,17'd10566,17'd10698,17'd9989,17'd10122,17'd10568,17'd10699,17'd9849,17'd9445,17'd10818,17'd10701,17'd9447,17'd9587,17'd10129,17'd9169,17'd9171,17'd10703,17'd10819,17'd10820,17'd10705,17'd10821,17'd10822,17'd10823,17'd10707,17'd10824,17'd10825,17'd10826,17'd10827,17'd10828,17'd10829,17'd10830,17'd10831,17'd10832,17'd10833,17'd10717,17'd10834,17'd10835,17'd10836,17'd10837,17'd10838,17'd10153,17'd10317,17'd10839,17'd10840,17'd10840,17'd10840,17'd10841,17'd10842,17'd10843,17'd10319,17'd10157,17'd10158,17'd10844,17'd10845,17'd10846,17'd10846,17'd10847,17'd10848,17'd10848,17'd10849,17'd10850,17'd10851,17'd10852,17'd10737,17'd10737,17'd10853,17'd10854,17'd10739,17'd10855,17'd10741,17'd10856,17'd9473,17'd10743,17'd9341,17'd10857,17'd10744,17'd9192,17'd9188,17'd10858,17'd10859,17'd10860,17'd10861,17'd10862,17'd10863,17'd10864,17'd10865,17'd10866,17'd10867,17'd10868,17'd10869,17'd10870,17'd10871,17'd10872,17'd10620,17'd10758,17'd10351,17'd10873,17'd10874,17'd1045,17'd134,17'd1045,17'd1045,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd135,17'd131,17'd7649,17'd8752,17'd10875,17'd10876,17'd10877,17'd10878,17'd10879,17'd10880,17'd10881,17'd8912,17'd10198,17'd10882,17'd10199,17'd10883,17'd8759,17'd7497,17'd7498,17'd8613,17'd10201,17'd10884,17'd10885,17'd10886,17'd10887,17'd9643,17'd9375,17'd9508,17'd9644,17'd9644,17'd9644,17'd9644,17'd10888,17'd9075,17'd9648,17'd9776,17'd8461,17'd10889,17'd10890,17'd10891,17'd10892,17'd10064,17'd10508,17'd10508,17'd10064,17'd10064,17'd10064,17'd10064,17'd10508,17'd10509,17'd10509,17'd10509,17'd10508,17'd10064,17'd10893,17'd10224,17'd10224,17'd10224,17'd10225,17'd10894,17'd10894,17'd10227,17'd10773,17'd9781,17'd9652,17'd10774,17'd10895,17'd10230,17'd10775,17'd10776,17'd10776,17'd10896,17'd9390,17'd10233,17'd6849,17'd7329,17'd9522,17'd8147,17'd8147,17'd7329,17'd7329,17'd7168,17'd6550,17'd6850,17'd10512,17'd6850,17'd6850,17'd8000,17'd6852,17'd9394,17'd9090,17'd8304,17'd9657,17'd10897,17'd10642,17'd10642,17'd10778,17'd10380,17'd8001,17'd6558,17'd6559,17'd6709,17'd6710,17'd10898,17'd10899,17'd7017,17'd10900,17'd10901,17'd10902,17'd10784,17'd10384,17'd10067,17'd10903,17'd10904,17'd10522,17'd10905,17'd10906,17'd5496,17'd10907,17'd3245,17'd2774,17'd5955,17'd9532,17'd3238,17'd3732,17'd2755,17'd3406,17'd7689,17'd8490,17'd7029,17'd7029,17'd8169,17'd8171,17'd9405,17'd10076,17'd9405,17'd10076,17'd10391,17'd9254,17'd9947,17'd10078,17'd9256,17'd9949,17'd9665,17'd8495,17'd8804,17'd7347,17'd7347,17'd7347,17'd7347,17'd7347,17'd9409,17'd9115,17'd9407,17'd9407,17'd9666,17'd9541,17'd8026,17'd7691,17'd10908,17'd10909,17'd10529,17'd10651,17'd8653,17'd10252,17'd8028,17'd8809,17'd7867,17'd7867,17'd7867,17'd7867,17'd8809,17'd8326,17'd7523,17'd7199,17'd10910,17'd10081,17'd9804,17'd9414,17'd7705,17'd7705,17'd7705,17'd7537,17'd8507,17'd7537,17'd7537,17'd7537,17'd5183,17'd9123,17'd5940,17'd5630,17'd6415,17'd6407,17'd604,17'd10911,17'd1408,17'd1669,17'd416,17'd195
},
'{
17'd4428,17'd4733,17'd2592,17'd2781,17'd1689,17'd14,17'd2,17'd12,17'd12,17'd12,17'd0,17'd0,17'd0,17'd2,17'd2,17'd1127,17'd6583,17'd4577,17'd7545,17'd7711,17'd1688,17'd1127,17'd12,17'd1275,17'd25,17'd8,17'd7,17'd5205,17'd10912,17'd10913,17'd10913,17'd10656,17'd10914,17'd7884,17'd8340,17'd10795,17'd10915,17'd10916,17'd8815,17'd6432,17'd8517,17'd7219,17'd9127,17'd8818,17'd8974,17'd8979,17'd8976,17'd10539,17'd7719,17'd8517,17'd7720,17'd7055,17'd8823,17'd10917,17'd10918,17'd10919,17'd9136,17'd10920,17'd7722,17'd10921,17'd7890,17'd10922,17'd10923,17'd3750,17'd10545,17'd10407,17'd10546,17'd10669,17'd10924,17'd10924,17'd10925,17'd10669,17'd292,17'd1693,17'd9816,17'd3907,17'd6598,17'd6598,17'd6903,17'd7556,17'd10408,17'd7730,17'd6281,17'd6281,17'd6443,17'd6443,17'd5223,17'd5386,17'd6751,17'd9971,17'd8990,17'd6911,17'd9558,17'd10412,17'd10926,17'd9974,17'd10803,17'd10927,17'd10928,17'd10929,17'd10930,17'd10931,17'd10807,17'd9429,17'd10932,17'd10933,17'd10934,17'd10935,17'd10936,17'd10937,17'd10938,17'd10939,17'd10688,17'd10940,17'd10941,17'd10941,17'd10108,17'd10814,17'd10942,17'd9572,17'd10285,17'd10427,17'd10563,17'd10816,17'd10817,17'd10943,17'd10944,17'd10943,17'd10945,17'd10945,17'd10428,17'd10428,17'd9574,17'd9574,17'd8537,17'd8537,17'd5409,17'd5409,17'd6140,17'd6140,17'd6305,17'd6305,17'd6305,17'd6305,17'd6465,17'd6465,17'd7085,17'd10946,17'd10431,17'd10431,17'd10432,17'd10696,17'd10697,17'd9844,17'd10947,17'd10948,17'd10949,17'd10288,17'd10122,17'd10700,17'd10433,17'd10434,17'd9310,17'd10818,17'd9313,17'd9587,17'd10129,17'd9448,17'd10435,17'd9711,17'd9592,17'd10132,17'd10950,17'd10951,17'd10952,17'd10953,17'd10954,17'd10955,17'd10956,17'd10957,17'd10958,17'd10959,17'd10960,17'd10961,17'd10962,17'd10831,17'd10963,17'd10964,17'd10965,17'd10966,17'd10967,17'd10968,17'd10969,17'd10970,17'd10839,17'd10971,17'd10972,17'd10973,17'd10973,17'd10974,17'd10975,17'd10976,17'd10977,17'd10978,17'd10979,17'd10980,17'd10980,17'd10981,17'd10982,17'd10983,17'd10983,17'd10984,17'd10985,17'd10985,17'd10986,17'd10987,17'd10988,17'd10737,17'd10989,17'd10853,17'd10990,17'd10739,17'd10991,17'd10164,17'd9739,17'd9885,17'd9341,17'd10743,17'd10992,17'd9341,17'd9339,17'd9038,17'd8727,17'd10993,17'd10994,17'd10995,17'd10996,17'd10997,17'd10998,17'd10999,17'd11000,17'd11001,17'd11002,17'd11003,17'd11004,17'd11005,17'd11006,17'd11007,17'd10491,17'd10621,17'd7812,17'd8132,17'd3025,17'd134,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd135,17'd131,17'd7649,17'd11008,17'd11009,17'd11010,17'd11011,17'd10878,17'd11012,17'd8451,17'd9066,17'd8143,17'd7824,17'd11013,17'd11014,17'd11015,17'd8611,17'd10362,17'd7498,17'd8613,17'd11016,17'd11017,17'd11018,17'd10886,17'd11019,17'd9375,17'd9508,17'd10888,17'd9227,17'd9227,17'd9227,17'd9644,17'd9770,17'd11020,17'd9648,17'd9776,17'd11021,17'd11022,17'd11023,17'd11024,17'd11025,17'd11026,17'd10893,17'd11027,17'd11027,17'd11027,17'd11027,17'd11027,17'd11027,17'd11028,17'd11028,17'd11029,17'd11029,17'd11028,17'd11028,17'd10893,17'd11030,17'd11026,17'd10893,17'd10225,17'd10227,17'd10894,17'd10894,17'd9384,17'd9518,17'd9651,17'd9652,17'd10228,17'd11031,17'd10511,17'd10776,17'd11032,17'd9389,17'd11033,17'd10231,17'd7010,17'd7329,17'd7329,17'd6849,17'd7329,17'd7329,17'd7168,17'd7168,17'd6550,17'd6385,17'd11034,17'd11035,17'd10236,17'd10236,17'd11036,17'd11036,17'd9932,17'd9394,17'd10513,17'd10514,17'd11037,17'd11038,17'd11038,17'd10779,17'd8001,17'd11039,17'd8001,17'd6709,17'd11040,17'd10898,17'd7016,17'd7184,17'd11041,17'd11042,17'd11043,17'd10784,17'd10384,17'd11044,17'd9939,17'd11045,17'd11046,17'd11047,17'd11048,17'd11049,17'd2739,17'd2765,17'd3894,17'd3889,17'd3584,17'd3888,17'd6252,17'd4565,17'd7196,17'd7195,17'd8490,17'd7687,17'd8794,17'd8794,17'd8171,17'd10076,17'd11050,17'd10076,17'd9946,17'd10526,17'd9255,17'd11051,17'd10249,17'd9256,17'd9538,17'd11052,17'd8495,17'd9409,17'd7347,17'd7347,17'd8490,17'd7347,17'd9409,17'd8495,17'd9665,17'd11053,17'd11054,17'd9541,17'd8026,17'd7691,17'd10908,17'd10908,17'd10909,17'd10529,17'd11055,17'd11056,17'd11057,17'd11058,17'd8809,17'd10653,17'd8326,17'd8809,17'd8809,17'd7867,17'd9799,17'd11059,17'd8655,17'd8656,17'd10082,17'd11060,17'd9414,17'd7705,17'd9124,17'd7538,17'd7537,17'd7537,17'd11061,17'd11061,17'd5183,17'd4714,17'd3073,17'd5940,17'd6415,17'd5372,17'd11062,17'd1408,17'd202,17'd421,17'd195,17'd1673
},
'{
17'd4246,17'd4887,17'd2781,17'd1967,17'd14,17'd2,17'd12,17'd3,17'd12,17'd12,17'd0,17'd2,17'd2,17'd2,17'd2,17'd1127,17'd6096,17'd4577,17'd7545,17'd4886,17'd1127,17'd2,17'd806,17'd2591,17'd4,17'd6,17'd5205,17'd5205,17'd10912,17'd10913,17'd10913,17'd10913,17'd7884,17'd7884,17'd8340,17'd10658,17'd11063,17'd9135,17'd9272,17'd11064,17'd7548,17'd8515,17'd9127,17'd8819,17'd8975,17'd8979,17'd8977,17'd10539,17'd7720,17'd11065,17'd7054,17'd10799,17'd6899,17'd11066,17'd11067,17'd11068,17'd7222,17'd10263,17'd7217,17'd11069,17'd11064,17'd11070,17'd9968,17'd2781,17'd10406,17'd10545,17'd10802,17'd10670,17'd11071,17'd10924,17'd10925,17'd11072,17'd1834,17'd655,17'd11073,17'd11073,17'd10269,17'd10093,17'd9555,17'd10409,17'd10672,17'd6281,17'd6282,17'd6281,17'd6443,17'd5813,17'd5386,17'd9818,17'd10270,17'd9280,17'd6911,17'd11074,17'd11075,17'd9689,17'd9824,17'd10414,17'd11076,17'd10928,17'd11077,17'd10680,17'd11078,17'd11079,17'd10681,17'd11080,17'd11081,17'd11082,17'd11083,17'd10936,17'd11084,17'd10938,17'd10938,17'd11085,17'd10940,17'd10940,17'd11086,17'd11086,17'd10108,17'd10814,17'd9572,17'd10690,17'd10427,17'd11087,17'd10816,17'd10816,17'd10943,17'd10944,17'd10944,17'd11088,17'd10945,17'd10945,17'd10428,17'd9574,17'd9574,17'd8537,17'd8537,17'd7750,17'd5837,17'd5837,17'd6140,17'd6140,17'd11089,17'd11089,17'd11089,17'd6305,17'd6465,17'd6465,17'd7085,17'd10946,17'd10431,17'd11090,17'd11091,17'd10696,17'd10697,17'd10566,17'd10948,17'd11092,17'd10288,17'd9990,17'd10569,17'd9992,17'd11093,17'd11094,17'd11095,17'd9019,17'd9447,17'd10129,17'd9448,17'd10435,17'd9319,17'd11096,17'd11097,17'd9713,17'd11098,17'd11099,17'd11100,17'd11101,17'd11102,17'd11103,17'd10957,17'd11104,17'd11105,17'd11106,17'd11107,17'd11108,17'd11109,17'd11110,17'd11111,17'd11112,17'd11113,17'd11114,17'd11115,17'd11116,17'd10971,17'd10971,17'd10972,17'd11117,17'd11118,17'd11118,17'd11119,17'd10971,17'd10975,17'd10976,17'd11120,17'd11121,17'd11122,17'd11123,17'd10983,17'd11124,17'd11125,17'd11126,17'd11127,17'd11128,17'd10596,17'd10159,17'd10322,17'd10469,17'd10988,17'd10853,17'd11129,17'd11130,17'd11131,17'd11132,17'd11133,17'd11134,17'd11135,17'd9741,17'd11136,17'd10992,17'd9885,17'd9885,17'd9340,17'd9192,17'd8722,17'd11137,17'd11138,17'd11139,17'd11140,17'd11141,17'd11142,17'd11143,17'd11144,17'd11145,17'd11146,17'd11147,17'd11148,17'd11149,17'd11150,17'd10188,17'd11151,17'd9495,17'd9359,17'd11152,17'd1045,17'd134,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd5593,17'd11153,17'd11154,17'd11155,17'd4348,17'd8906,17'd11156,17'd11157,17'd10881,17'd11158,17'd10198,17'd10882,17'd11159,17'd11160,17'd8611,17'd10362,17'd8613,17'd11161,17'd11016,17'd11162,17'd11163,17'd11164,17'd9643,17'd9375,17'd10888,17'd9227,17'd9227,17'd9227,17'd9227,17'd10502,17'd9770,17'd8921,17'd11165,17'd11166,17'd11167,17'd11168,17'd11169,17'd11170,17'd11170,17'd11171,17'd11172,17'd10893,17'd11027,17'd11027,17'd11027,17'd10893,17'd11027,17'd11027,17'd11027,17'd11028,17'd11028,17'd11029,17'd11029,17'd11173,17'd11174,17'd10893,17'd11026,17'd10224,17'd10377,17'd10226,17'd10894,17'd11175,17'd10226,17'd9780,17'd9651,17'd9651,17'd9652,17'd10229,17'd11032,17'd11176,17'd11032,17'd11177,17'd10896,17'd10232,17'd6849,17'd6849,17'd7010,17'd6849,17'd7329,17'd7168,17'd7991,17'd7168,17'd6386,17'd11034,17'd11178,17'd11035,17'd10236,17'd10236,17'd11179,17'd11180,17'd9932,17'd10513,17'd10777,17'd11181,17'd11037,17'd11037,17'd11038,17'd10380,17'd8001,17'd8001,17'd8001,17'd6709,17'd6561,17'd7330,17'd7016,17'd11182,17'd11183,17'd10901,17'd11184,17'd10784,17'd10384,17'd10243,17'd11185,17'd11186,17'd11187,17'd11188,17'd5356,17'd5497,17'd3245,17'd3422,17'd3585,17'd3414,17'd3238,17'd4075,17'd6578,17'd4070,17'd7196,17'd7688,17'd10248,17'd8794,17'd11189,17'd7856,17'd9405,17'd11190,17'd11191,17'd9405,17'd9946,17'd9254,17'd9110,17'd10078,17'd11192,17'd9949,17'd9538,17'd9665,17'd8495,17'd7347,17'd7347,17'd8490,17'd8490,17'd9250,17'd8495,17'd9665,17'd11053,17'd11054,17'd9666,17'd8026,17'd7691,17'd11193,17'd8964,17'd8964,17'd10529,17'd11055,17'd11055,17'd11056,17'd11194,17'd8809,17'd11195,17'd9259,17'd8809,17'd8809,17'd8809,17'd9955,17'd11195,17'd9668,17'd11196,17'd9957,17'd11197,17'd9414,17'd7705,17'd9124,17'd7538,17'd7705,17'd7705,17'd11061,17'd11061,17'd2906,17'd4714,17'd9123,17'd5940,17'd1946,17'd6415,17'd11062,17'd423,17'd1526,17'd419,17'd1813,17'd1530
},
'{
17'd3250,17'd1688,17'd1689,17'd1127,17'd2,17'd12,17'd12,17'd3,17'd0,17'd0,17'd0,17'd0,17'd14,17'd14,17'd1127,17'd1689,17'd4577,17'd4887,17'd7545,17'd5196,17'd2,17'd12,17'd2933,17'd978,17'd6,17'd3753,17'd5205,17'd8040,17'd10913,17'd10913,17'd10913,17'd10913,17'd10913,17'd10656,17'd8190,17'd11198,17'd6588,17'd9136,17'd11199,17'd8517,17'd7219,17'd7716,17'd9548,17'd10798,17'd10798,17'd10262,17'd9128,17'd8974,17'd8517,17'd11200,17'd6431,17'd10403,17'd10541,17'd11201,17'd11202,17'd11203,17'd11204,17'd7885,17'd7217,17'd11064,17'd11205,17'd11206,17'd2592,17'd2781,17'd10546,17'd3593,17'd10924,17'd10924,17'd10925,17'd10925,17'd292,17'd11207,17'd11208,17'd11209,17'd11210,17'd10269,17'd6746,17'd11211,17'd10408,17'd10408,17'd6112,17'd10548,17'd10548,17'd5811,17'd11212,17'd11213,17'd5386,17'd6751,17'd10411,17'd8831,17'd9972,17'd11075,17'd11214,17'd10414,17'd11215,17'd11216,17'd11217,17'd11218,17'd10680,17'd10931,17'd11219,17'd8681,17'd11220,17'd11221,17'd11222,17'd11223,17'd11224,17'd11225,17'd11226,17'd11227,17'd10688,17'd10561,17'd10940,17'd11228,17'd10941,17'd10941,17'd10108,17'd10814,17'd11229,17'd11230,17'd10563,17'd10816,17'd10817,17'd10943,17'd10943,17'd10944,17'd11231,17'd10944,17'd10945,17'd10692,17'd11232,17'd9158,17'd9159,17'd8537,17'd7418,17'd5837,17'd5837,17'd5689,17'd6140,17'd6626,17'd6626,17'd6626,17'd10695,17'd10114,17'd10946,17'd6625,17'd7251,17'd7251,17'd11233,17'd7581,17'd10119,17'd9844,17'd11234,17'd11235,17'd11236,17'd11237,17'd10568,17'd9991,17'd9991,17'd9849,17'd11238,17'd11239,17'd9585,17'd10571,17'd9587,17'd9315,17'd10435,17'd11240,17'd10703,17'd9452,17'd10297,17'd10705,17'd10822,17'd11099,17'd11241,17'd11242,17'd11243,17'd11103,17'd11244,17'd11245,17'd11246,17'd11247,17'd11248,17'd11249,17'd11250,17'd11251,17'd11252,17'd11253,17'd11254,17'd11255,17'd11256,17'd11119,17'd11119,17'd11119,17'd11118,17'd11257,17'd11258,17'd11259,17'd11260,17'd10971,17'd10840,17'd10725,17'd11261,17'd11262,17'd11263,17'd11264,17'd11265,17'd11266,17'd11267,17'd11268,17'd11269,17'd11270,17'd10157,17'd11271,17'd11272,17'd11273,17'd10852,17'd10736,17'd11274,17'd11275,17'd10854,17'd11132,17'd11133,17'd11134,17'd11276,17'd11277,17'd9885,17'd10992,17'd9885,17'd9741,17'd10743,17'd9347,17'd8721,17'd8727,17'd8413,17'd11278,17'd11279,17'd11280,17'd11281,17'd11282,17'd11283,17'd11284,17'd11285,17'd10868,17'd11286,17'd11287,17'd11288,17'd7809,17'd11007,17'd8750,17'd9359,17'd11289,17'd3025,17'd1197,17'd1197,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd5593,17'd5593,17'd6831,17'd11290,17'd11291,17'd11292,17'd11293,17'd9761,17'd7001,17'd8607,17'd11294,17'd10359,17'd10882,17'd11159,17'd11295,17'd8611,17'd11296,17'd8612,17'd11161,17'd10202,17'd11297,17'd11163,17'd11298,17'd10769,17'd9644,17'd10888,17'd11299,17'd11300,17'd11300,17'd11301,17'd11302,17'd9512,17'd8921,17'd8296,17'd9777,17'd11303,17'd11169,17'd11304,17'd11305,17'd11306,17'd11170,17'd11171,17'd11025,17'd11172,17'd10893,17'd11028,17'd11028,17'd11028,17'd11027,17'd11027,17'd10893,17'd11027,17'd11028,17'd11029,17'd11307,17'd11308,17'd11174,17'd11174,17'd10893,17'd10893,17'd11027,17'd11027,17'd11309,17'd10227,17'd10227,17'd10226,17'd9780,17'd10063,17'd11310,17'd10228,17'd9389,17'd10775,17'd10511,17'd9388,17'd9653,17'd10775,17'd7010,17'd6849,17'd6849,17'd6849,17'd6849,17'd6849,17'd6550,17'd6550,17'd6386,17'd11311,17'd11312,17'd10512,17'd10236,17'd11036,17'd11313,17'd11314,17'd11315,17'd10777,17'd11181,17'd11316,17'd11317,17'd11318,17'd11038,17'd10380,17'd9934,17'd11039,17'd6709,17'd6560,17'd6856,17'd8475,17'd11319,17'd11320,17'd11321,17'd11043,17'd9241,17'd11322,17'd11323,17'd11324,17'd11325,17'd11326,17'd11327,17'd11048,17'd11328,17'd2391,17'd1945,17'd3741,17'd3889,17'd9532,17'd3581,17'd4075,17'd2755,17'd3407,17'd4413,17'd8803,17'd10248,17'd10248,17'd8169,17'd7856,17'd11191,17'd11191,17'd9405,17'd8955,17'd9536,17'd9110,17'd11329,17'd10078,17'd11330,17'd9112,17'd9539,17'd9408,17'd8174,17'd7517,17'd7686,17'd7687,17'd8804,17'd8804,17'd8495,17'd11331,17'd9538,17'd8801,17'd8962,17'd9953,17'd7691,17'd8499,17'd10908,17'd8027,17'd10529,17'd10651,17'd11056,17'd11056,17'd8809,17'd7867,17'd7867,17'd7867,17'd8809,17'd8809,17'd9955,17'd9955,17'd10080,17'd11332,17'd11333,17'd10082,17'd11334,17'd7705,17'd7538,17'd9124,17'd11335,17'd11336,17'd11061,17'd11061,17'd11061,17'd5183,17'd9123,17'd5940,17'd5372,17'd5372,17'd11337,17'd423,17'd1529,17'd600,17'd1813,17'd2102
},
'{
17'd1688,17'd1689,17'd1127,17'd2,17'd13,17'd12,17'd12,17'd3,17'd0,17'd0,17'd0,17'd14,17'd14,17'd1127,17'd1127,17'd1688,17'd4577,17'd4887,17'd4886,17'd6419,17'd13,17'd2423,17'd4242,17'd7373,17'd3753,17'd5205,17'd8040,17'd8340,17'd10913,17'd10913,17'd10913,17'd10913,17'd10913,17'd11338,17'd10536,17'd5648,17'd6596,17'd7885,17'd7715,17'd7549,17'd7377,17'd7377,17'd10798,17'd10798,17'd11339,17'd10400,17'd9267,17'd9678,17'd11340,17'd10399,17'd9680,17'd7056,17'd8984,17'd11341,17'd11342,17'd11201,17'd9966,17'd9551,17'd7722,17'd10922,17'd11343,17'd11344,17'd7371,17'd2592,17'd3593,17'd10669,17'd10924,17'd10924,17'd10924,17'd10924,17'd292,17'd11207,17'd11209,17'd11209,17'd11210,17'd10269,17'd6746,17'd11211,17'd10408,17'd11345,17'd6111,17'd5662,17'd5662,17'd5385,17'd5523,17'd5523,17'd5387,17'd10411,17'd11346,17'd11347,17'd9822,17'd10413,17'd11348,17'd11216,17'd11349,17'd11218,17'd11350,17'd9428,17'd11351,17'd11079,17'd11352,17'd9152,17'd11353,17'd11354,17'd10809,17'd11355,17'd11356,17'd11357,17'd11358,17'd10811,17'd10424,17'd10279,17'd10941,17'd10941,17'd11086,17'd11359,17'd10814,17'd11360,17'd11361,17'd11362,17'd10816,17'd10816,17'd11088,17'd10943,17'd10944,17'd10944,17'd11231,17'd10944,17'd10564,17'd10564,17'd11232,17'd11232,17'd9159,17'd8537,17'd5409,17'd5837,17'd5689,17'd5689,17'd6626,17'd6626,17'd6626,17'd6140,17'd10695,17'd7085,17'd6625,17'd6625,17'd7251,17'd7251,17'd7581,17'd10696,17'd10697,17'd9844,17'd11363,17'd11235,17'd11236,17'd10568,17'd9991,17'd9848,17'd9848,17'd9583,17'd11239,17'd10818,17'd9312,17'd11364,17'd10129,17'd9590,17'd9319,17'd11365,17'd11366,17'd11097,17'd10573,17'd11367,17'd10822,17'd10953,17'd11368,17'd11369,17'd11370,17'd11371,17'd11245,17'd11372,17'd11373,17'd11247,17'd11374,17'd11375,17'd11376,17'd11377,17'd11378,17'd11379,17'd11380,17'd11381,17'd11382,17'd11383,17'd11384,17'd11385,17'd11385,17'd11382,17'd11382,17'd11259,17'd11260,17'd10971,17'd11386,17'd11387,17'd11388,17'd11389,17'd11390,17'd11390,17'd11390,17'd11391,17'd11392,17'd11388,17'd11393,17'd11269,17'd11128,17'd10985,17'd10986,17'd11394,17'd10735,17'd11395,17'd11396,17'd11397,17'd11398,17'd11399,17'd11400,17'd10329,17'd11401,17'd11276,17'd9884,17'd9885,17'd10169,17'd10024,17'd10992,17'd9339,17'd11402,17'd11403,17'd11404,17'd11405,17'd11406,17'd11407,17'd7457,17'd8112,17'd9894,17'd11408,17'd11409,17'd11410,17'd11411,17'd11412,17'd11288,17'd7809,17'd11007,17'd8750,17'd9359,17'd11152,17'd11413,17'd1197,17'd1197,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd5593,17'd5593,17'd11414,17'd11415,17'd11416,17'd11417,17'd11418,17'd11419,17'd11420,17'd10881,17'd11294,17'd10882,17'd11421,17'd11422,17'd11423,17'd9505,17'd8761,17'd10201,17'd11424,17'd10202,17'd11162,17'd11163,17'd10769,17'd11425,17'd10888,17'd9228,17'd11301,17'd11300,17'd11300,17'd9228,17'd9075,17'd8921,17'd9648,17'd9776,17'd11021,17'd11426,17'd11169,17'd11427,17'd11305,17'd11306,17'd11171,17'd11025,17'd11025,17'd11172,17'd11026,17'd10893,17'd11027,17'd11027,17'd11028,17'd11028,17'd11028,17'd11027,17'd11028,17'd11028,17'd11428,17'd11428,17'd11428,17'd11308,17'd11027,17'd11027,17'd11027,17'd11028,17'd11309,17'd11309,17'd10227,17'd10227,17'd10226,17'd9780,17'd9517,17'd10063,17'd10228,17'd9519,17'd10230,17'd10230,17'd9519,17'd9388,17'd10230,17'd10234,17'd7010,17'd6849,17'd7329,17'd6849,17'd6550,17'd6550,17'd6386,17'd6385,17'd11035,17'd11312,17'd11179,17'd11036,17'd11180,17'd11314,17'd11429,17'd11430,17'd11181,17'd11431,17'd11317,17'd11432,17'd11317,17'd11038,17'd9934,17'd10238,17'd6558,17'd7501,17'd6561,17'd8157,17'd11433,17'd11319,17'd11434,17'd11321,17'd11435,17'd11436,17'd11437,17'd11438,17'd11439,17'd11440,17'd11441,17'd11442,17'd4711,17'd4556,17'd2095,17'd11443,17'd3585,17'd9532,17'd3582,17'd3885,17'd6578,17'd3406,17'd4567,17'd10390,17'd7687,17'd10248,17'd8169,17'd7856,17'd11444,17'd11191,17'd9405,17'd9405,17'd10391,17'd10650,17'd9110,17'd10078,17'd9948,17'd11330,17'd9538,17'd9407,17'd8495,17'd8174,17'd7517,17'd7687,17'd8804,17'd9250,17'd8495,17'd11331,17'd9538,17'd9407,17'd9541,17'd8962,17'd7691,17'd7691,17'd11193,17'd8027,17'd9259,17'd10651,17'd11055,17'd11056,17'd8809,17'd7867,17'd7867,17'd7867,17'd7867,17'd8809,17'd9955,17'd9955,17'd10080,17'd9956,17'd10910,17'd9957,17'd9804,17'd9544,17'd7705,17'd9124,17'd11336,17'd11336,17'd11061,17'd11061,17'd11061,17'd11336,17'd9123,17'd9123,17'd5630,17'd6415,17'd11062,17'd11445,17'd1529,17'd417,17'd1947,17'd2102
},
'{
17'd1127,17'd1127,17'd2,17'd2,17'd12,17'd12,17'd12,17'd12,17'd0,17'd2,17'd14,17'd14,17'd14,17'd1689,17'd4886,17'd7214,17'd7545,17'd7545,17'd4247,17'd2,17'd806,17'd2933,17'd23,17'd6,17'd5205,17'd5205,17'd8040,17'd8340,17'd8340,17'd8340,17'd8339,17'd8339,17'd8340,17'd10537,17'd7375,17'd11446,17'd8669,17'd11199,17'd7889,17'd7053,17'd11447,17'd11447,17'd11448,17'd10540,17'd11449,17'd10539,17'd9678,17'd11450,17'd8667,17'd7376,17'd7056,17'd7379,17'd11451,17'd11452,17'd9681,17'd9133,17'd7885,17'd6429,17'd6429,17'd11453,17'd11454,17'd6424,17'd10407,17'd3593,17'd10669,17'd10924,17'd10925,17'd10924,17'd32,17'd292,17'd470,17'd1834,17'd11209,17'd11209,17'd11210,17'd6278,17'd6746,17'd11211,17'd6279,17'd6111,17'd5662,17'd5222,17'd5222,17'd5524,17'd11455,17'd6910,17'd11456,17'd11457,17'd11458,17'd9822,17'd10273,17'd11459,17'd11460,17'd11461,17'd11462,17'd11463,17'd11464,17'd11465,17'd11466,17'd11467,17'd11468,17'd11469,17'd11470,17'd11471,17'd11472,17'd11224,17'd11473,17'd11358,17'd11474,17'd10811,17'd10424,17'd11475,17'd11476,17'd10941,17'd11086,17'd11359,17'd11477,17'd11478,17'd11230,17'd11362,17'd10816,17'd10816,17'd11088,17'd10943,17'd10944,17'd10944,17'd10944,17'd10944,17'd9158,17'd11232,17'd11232,17'd11232,17'd9159,17'd8537,17'd5409,17'd5409,17'd5689,17'd5255,17'd11479,17'd6626,17'd6140,17'd7085,17'd6140,17'd6140,17'd7417,17'd8368,17'd7415,17'd7415,17'd8844,17'd10119,17'd11480,17'd11363,17'd11481,17'd11482,17'd11483,17'd10289,17'd11484,17'd11093,17'd9309,17'd9310,17'd10818,17'd10701,17'd9313,17'd8856,17'd9170,17'd9591,17'd10703,17'd11366,17'd11485,17'd10297,17'd11486,17'd11487,17'd11488,17'd11489,17'd11490,17'd11491,17'd11492,17'd11493,17'd11372,17'd11494,17'd11495,17'd11496,17'd11497,17'd11498,17'd11499,17'd11500,17'd11501,17'd11502,17'd11503,17'd11504,17'd11505,17'd11506,17'd11507,17'd11507,17'd11507,17'd11384,17'd11382,17'd11257,17'd11260,17'd10972,17'd11508,17'd11509,17'd11510,17'd11510,17'd11511,17'd11512,17'd11513,17'd11513,17'd11514,17'd11515,17'd10725,17'd11269,17'd11516,17'd10980,17'd11517,17'd11518,17'd11519,17'd11520,17'd11521,17'd11522,17'd11523,17'd11524,17'd11525,17'd11526,17'd11527,17'd11528,17'd11276,17'd9884,17'd9884,17'd9741,17'd10743,17'd9342,17'd11529,17'd11530,17'd9482,17'd11531,17'd11532,17'd11533,17'd11534,17'd7459,17'd11535,17'd11536,17'd11537,17'd11538,17'd10754,17'd11539,17'd11540,17'd9630,17'd7976,17'd8750,17'd9359,17'd6529,17'd6198,17'd3025,17'd889,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd11541,17'd5593,17'd6370,17'd11542,17'd11543,17'd11544,17'd3670,17'd11545,17'd11546,17'd10881,17'd11547,17'd11548,17'd11549,17'd11550,17'd11551,17'd9505,17'd9505,17'd9641,17'd10202,17'd10202,17'd9374,17'd11552,17'd11425,17'd10888,17'd10502,17'd9228,17'd9228,17'd11553,17'd11553,17'd11554,17'd11555,17'd9513,17'd11556,17'd11166,17'd11557,17'd11426,17'd11169,17'd11558,17'd11559,17'd11560,17'd11023,17'd11024,17'd11023,17'd11024,17'd11561,17'd11562,17'd10892,17'd10218,17'd11563,17'd11564,17'd11029,17'd11028,17'd11173,17'd11173,17'd11028,17'd11565,17'd11566,17'd11566,17'd11029,17'd11028,17'd11028,17'd11029,17'd11309,17'd11309,17'd11309,17'd11309,17'd11309,17'd10510,17'd10510,17'd10226,17'd9517,17'd9651,17'd10229,17'd11567,17'd11031,17'd9652,17'd10774,17'd10230,17'd11176,17'd11568,17'd11569,17'd11569,17'd6386,17'd6386,17'd6386,17'd6385,17'd6850,17'd11570,17'd11571,17'd11572,17'd11573,17'd11574,17'd11575,17'd11315,17'd10641,17'd11576,17'd11577,17'd11578,17'd11579,17'd11317,17'd10515,17'd10238,17'd7011,17'd6559,17'd7501,17'd6712,17'd7841,17'd7332,17'd11580,17'd11581,17'd11435,17'd9241,17'd11582,17'd11323,17'd11583,17'd11584,17'd11585,17'd11586,17'd11587,17'd11588,17'd11589,17'd11590,17'd5192,17'd11591,17'd3411,17'd3581,17'd4075,17'd4410,17'd4568,17'd4567,17'd8490,17'd7687,17'd8169,17'd7856,17'd8170,17'd8491,17'd8795,17'd9405,17'd11592,17'd11593,17'd9110,17'd11594,17'd10078,17'd10249,17'd11595,17'd9538,17'd9950,17'd8174,17'd7517,17'd11596,17'd8804,17'd9250,17'd9409,17'd9950,17'd9539,17'd9539,17'd9666,17'd9541,17'd8650,17'd9953,17'd9411,17'd8499,17'd8027,17'd10529,17'd10651,17'd8653,17'd9667,17'd8500,17'd7867,17'd7867,17'd9799,17'd9955,17'd8181,17'd8181,17'd9799,17'd10256,17'd11597,17'd11333,17'd11598,17'd11599,17'd7705,17'd7705,17'd11061,17'd11061,17'd11061,17'd11061,17'd11336,17'd11335,17'd9123,17'd9123,17'd5940,17'd5630,17'd11600,17'd11445,17'd415,17'd417,17'd1947,17'd11601
},
'{
17'd14,17'd14,17'd2,17'd0,17'd12,17'd12,17'd12,17'd0,17'd0,17'd14,17'd1127,17'd1689,17'd1967,17'd1689,17'd7214,17'd7372,17'd7372,17'd4886,17'd466,17'd12,17'd2933,17'd4242,17'd5,17'd6,17'd5205,17'd5205,17'd8040,17'd8340,17'd8340,17'd8340,17'd8339,17'd8339,17'd8040,17'd10536,17'd5648,17'd8042,17'd9551,17'd11602,17'd8517,17'd7053,17'd11448,17'd10798,17'd11447,17'd10262,17'd11603,17'd10539,17'd11339,17'd8345,17'd11604,17'd7885,17'd11605,17'd10541,17'd11606,17'd9545,17'd7056,17'd9680,17'd6590,17'd7376,17'd11607,17'd11608,17'd2782,17'd2592,17'd10407,17'd11072,17'd10924,17'd10925,17'd11609,17'd10924,17'd292,17'd470,17'd1834,17'd11207,17'd11209,17'd9816,17'd6278,17'd6278,17'd6746,17'd11211,17'd6279,17'd5976,17'd11610,17'd11611,17'd6284,17'd11612,17'd7394,17'd8674,17'd11613,17'd11614,17'd11615,17'd10273,17'd11459,17'd11616,17'd11617,17'd11462,17'd11618,17'd11466,17'd11619,17'd11620,17'd9563,17'd11468,17'd11621,17'd11622,17'd11082,17'd11623,17'd11624,17'd11356,17'd11357,17'd11226,17'd11227,17'd10938,17'd11625,17'd11475,17'd10941,17'd10941,17'd11359,17'd11626,17'd11627,17'd11628,17'd11362,17'd11629,17'd10816,17'd10816,17'd10943,17'd10944,17'd10944,17'd10944,17'd10944,17'd10943,17'd9158,17'd11232,17'd11232,17'd9006,17'd8537,17'd5409,17'd5409,17'd5409,17'd5255,17'd5255,17'd6626,17'd6626,17'd6140,17'd6140,17'd6140,17'd6468,17'd8368,17'd8368,17'd7415,17'd7579,17'd10119,17'd9844,17'd11235,17'd11235,17'd11482,17'd11483,17'd10289,17'd11484,17'd11630,17'd11094,17'd11631,17'd11095,17'd9446,17'd9313,17'd9167,17'd9170,17'd9171,17'd11632,17'd11366,17'd11633,17'd11634,17'd10573,17'd11487,17'd11635,17'd11636,17'd11101,17'd11637,17'd11638,17'd11639,17'd11640,17'd11372,17'd11641,17'd11495,17'd11642,17'd11643,17'd11644,17'd11645,17'd11646,17'd11647,17'd11648,17'd11649,17'd11650,17'd11651,17'd11652,17'd11653,17'd11653,17'd11654,17'd11505,17'd11384,17'd11118,17'd11655,17'd11655,17'd11655,17'd11656,17'd11657,17'd11658,17'd11659,17'd11660,17'd11661,17'd11662,17'd10973,17'd10840,17'd11268,17'd11127,17'd10982,17'd11663,17'd11664,17'd11665,17'd11666,17'd11667,17'd11667,17'd11521,17'd11522,17'd11523,17'd11668,17'd11669,17'd10476,17'd11527,17'd11670,17'd11276,17'd11671,17'd9884,17'd9885,17'd9344,17'd8720,17'd11530,17'd11672,17'd9886,17'd11673,17'd11674,17'd7786,17'd11675,17'd11676,17'd11677,17'd11678,17'd11679,17'd11680,17'd11681,17'd11682,17'd9630,17'd7976,17'd8750,17'd9359,17'd11152,17'd11413,17'd3025,17'd889,17'd1045,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd131,17'd11683,17'd11684,17'd11685,17'd11686,17'd11687,17'd11688,17'd11689,17'd11690,17'd9215,17'd11691,17'd11692,17'd11549,17'd11422,17'd9640,17'd8762,17'd11693,17'd9912,17'd9642,17'd11694,17'd11694,17'd9071,17'd11695,17'd10502,17'd9228,17'd9228,17'd11696,17'd11553,17'd11554,17'd8920,17'd11697,17'd9774,17'd11698,17'd11699,17'd11167,17'd11426,17'd11560,17'd11560,17'd11023,17'd11700,17'd11701,17'd11168,17'd11702,17'd11168,17'd11023,17'd11561,17'd11024,17'd11562,17'd11703,17'd11564,17'd11029,17'd11029,17'd11308,17'd11308,17'd11028,17'd11565,17'd11704,17'd11704,17'd11566,17'd11565,17'd11565,17'd11565,17'd11705,17'd11309,17'd11309,17'd11309,17'd11309,17'd11309,17'd11309,17'd11309,17'd11309,17'd10226,17'd9780,17'd10774,17'd10229,17'd10229,17'd10228,17'd10228,17'd11706,17'd10776,17'd11568,17'd11568,17'd6385,17'd6385,17'd6385,17'd6551,17'd6850,17'd11312,17'd11571,17'd11707,17'd11573,17'd11708,17'd11429,17'd11575,17'd10641,17'd11576,17'd11709,17'd11710,17'd11711,17'd11711,17'd11316,17'd10380,17'd6558,17'd6559,17'd7501,17'd6711,17'd7331,17'd11433,17'd11182,17'd11434,17'd11581,17'd11712,17'd11713,17'd11714,17'd11715,17'd11716,17'd11717,17'd11718,17'd11719,17'd11720,17'd5027,17'd11589,17'd11721,17'd5956,17'd3088,17'd3411,17'd3885,17'd6578,17'd3232,17'd4568,17'd7689,17'd8490,17'd8169,17'd7856,17'd8018,17'd8170,17'd8795,17'd8795,17'd9405,17'd11722,17'd11593,17'd11723,17'd10078,17'd10078,17'd11724,17'd9112,17'd11052,17'd8495,17'd11596,17'd8320,17'd8804,17'd9250,17'd8496,17'd8495,17'd9539,17'd9538,17'd11725,17'd9666,17'd8650,17'd8650,17'd8324,17'd9411,17'd10908,17'd8027,17'd10529,17'd11726,17'd11727,17'd8500,17'd7867,17'd7867,17'd9799,17'd9955,17'd8181,17'd8181,17'd9955,17'd10256,17'd10654,17'd11196,17'd11728,17'd11060,17'd9544,17'd7705,17'd11061,17'd11061,17'd11061,17'd11061,17'd11336,17'd11335,17'd9123,17'd9123,17'd5630,17'd5630,17'd11600,17'd11445,17'd776,17'd1813,17'd11729,17'd11601
},
'{
17'd2,17'd0,17'd0,17'd0,17'd12,17'd12,17'd0,17'd0,17'd2,17'd14,17'd1127,17'd1689,17'd5196,17'd7711,17'd7545,17'd7372,17'd1831,17'd1127,17'd12,17'd1275,17'd23,17'd5,17'd6,17'd5205,17'd5205,17'd5205,17'd5205,17'd8190,17'd8340,17'd8340,17'd8339,17'd8340,17'd8190,17'd5378,17'd11730,17'd9137,17'd11731,17'd8666,17'd7054,17'd7221,17'd11732,17'd10798,17'd10262,17'd11449,17'd10539,17'd11450,17'd8345,17'd11733,17'd11199,17'd10263,17'd10542,17'd9137,17'd6103,17'd9415,17'd6430,17'd6740,17'd11734,17'd11735,17'd11736,17'd6265,17'd10268,17'd10268,17'd3593,17'd11071,17'd656,17'd811,17'd984,17'd33,17'd470,17'd1834,17'd3431,17'd11208,17'd3756,17'd3756,17'd5656,17'd5804,17'd11737,17'd11737,17'd11738,17'd11739,17'd11740,17'd5062,17'd5063,17'd11741,17'd6912,17'd11742,17'd11743,17'd9824,17'd11744,17'd10927,17'd11745,17'd11746,17'd11747,17'd11748,17'd11749,17'd11750,17'd11751,17'd10932,17'd11752,17'd11753,17'd11754,17'd11755,17'd11756,17'd11757,17'd11758,17'd11759,17'd11760,17'd11357,17'd11761,17'd10687,17'd11762,17'd11625,17'd11086,17'd11476,17'd11477,17'd11763,17'd11478,17'd11764,17'd10815,17'd10815,17'd11087,17'd11087,17'd10944,17'd10944,17'd10692,17'd10564,17'd10564,17'd10564,17'd11232,17'd11232,17'd9159,17'd8537,17'd6143,17'd5837,17'd5409,17'd4927,17'd4927,17'd5255,17'd6626,17'd6626,17'd6468,17'd6468,17'd6141,17'd6141,17'd8368,17'd8218,17'd7748,17'd8065,17'd11480,17'd11765,17'd11766,17'd11482,17'd11483,17'd11483,17'd10289,17'd11484,17'd11630,17'd11094,17'd9310,17'd11095,17'd9019,17'd8703,17'd7266,17'd10435,17'd11767,17'd11768,17'd11769,17'd11770,17'd11771,17'd11486,17'd11487,17'd11772,17'd11773,17'd11490,17'd11774,17'd11775,17'd11776,17'd11777,17'd11778,17'd11779,17'd11780,17'd11642,17'd11781,17'd11782,17'd11783,17'd11784,17'd11785,17'd11786,17'd11787,17'd11788,17'd11789,17'd11790,17'd11791,17'd11791,17'd11792,17'd11793,17'd11507,17'd11794,17'd11795,17'd11796,17'd11795,17'd11797,17'd11798,17'd11799,17'd11800,17'd11506,17'd11660,17'd11662,17'd11510,17'd11801,17'd11802,17'd11124,17'd11803,17'd11804,17'd11805,17'd11806,17'd11806,17'd11806,17'd11806,17'd11807,17'd11807,17'd11522,17'd11396,17'd11808,17'd10854,17'd10476,17'd10991,17'd11670,17'd11276,17'd11277,17'd11809,17'd9344,17'd8873,17'd11810,17'd11530,17'd8412,17'd11811,17'd11812,17'd8254,17'd11813,17'd11814,17'd11815,17'd11816,17'd11817,17'd11818,17'd11819,17'd11820,17'd9898,17'd9358,17'd10037,17'd8597,17'd6529,17'd6198,17'd3025,17'd889,17'd889,17'd1197,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd131,17'd11821,17'd11822,17'd11823,17'd11824,17'd11825,17'd11826,17'd11827,17'd6540,17'd11828,17'd11829,17'd11830,17'd11549,17'd11831,17'd9505,17'd8762,17'd11017,17'd11162,17'd8917,17'd11832,17'd11832,17'd8918,17'd9075,17'd9228,17'd10502,17'd10502,17'd11833,17'd11695,17'd8920,17'd11834,17'd9774,17'd11835,17'd11166,17'd11699,17'd11167,17'd11836,17'd11701,17'd8776,17'd9927,17'd9778,17'd11836,17'd11837,17'd11837,17'd11167,17'd11836,17'd11022,17'd11022,17'd11838,17'd11562,17'd10218,17'd10064,17'd10509,17'd11565,17'd11565,17'd11839,17'd11839,17'd11566,17'd11566,17'd11704,17'd11840,17'd11841,17'd11842,17'd11843,17'd11843,17'd11844,17'd11844,17'd11845,17'd11845,17'd11846,17'd10510,17'd11309,17'd11309,17'd11309,17'd10226,17'd10063,17'd11847,17'd11847,17'd9652,17'd10774,17'd11706,17'd11176,17'd11848,17'd11849,17'd11849,17'd11850,17'd11851,17'd11850,17'd11851,17'd11707,17'd11571,17'd11707,17'd11572,17'd11313,17'd11852,17'd11576,17'd11576,17'd11853,17'd11854,17'd11579,17'd11855,17'd11579,17'd11856,17'd8001,17'd7836,17'd6559,17'd7501,17'd6712,17'd11433,17'd11319,17'd11580,17'd11857,17'd11858,17'd11859,17'd11860,17'd11861,17'd11862,17'd11863,17'd11864,17'd11865,17'd11866,17'd11867,17'd11868,17'd11869,17'd1810,17'd11870,17'd11871,17'd3412,17'd3727,17'd6725,17'd3406,17'd7518,17'd7688,17'd7029,17'd7858,17'd8794,17'd8954,17'd8491,17'd8795,17'd11191,17'd10076,17'd10077,17'd11872,17'd11051,17'd11329,17'd11873,17'd11874,17'd9538,17'd9408,17'd11875,17'd8320,17'd9797,17'd8804,17'd9409,17'd9409,17'd9408,17'd8800,17'd9538,17'd9407,17'd8649,17'd8650,17'd7690,17'd7864,17'd8499,17'd11876,17'd11877,17'd11877,17'd11878,17'd11727,17'd7867,17'd7867,17'd9799,17'd9799,17'd8181,17'd7698,17'd7698,17'd9955,17'd10080,17'd11879,17'd11880,17'd11881,17'd9414,17'd9544,17'd11882,17'd11061,17'd11061,17'd11061,17'd11336,17'd11335,17'd4714,17'd9123,17'd5630,17'd5630,17'd11600,17'd414,17'd1671,17'd1673,17'd11883,17'd11884
},
'{
17'd0,17'd0,17'd0,17'd1,17'd3,17'd12,17'd0,17'd2,17'd14,17'd1967,17'd1689,17'd1688,17'd7711,17'd7545,17'd7545,17'd7214,17'd4247,17'd2,17'd806,17'd2591,17'd4,17'd6,17'd5205,17'd5205,17'd5205,17'd5205,17'd8190,17'd8190,17'd8340,17'd8340,17'd8339,17'd8340,17'd7374,17'd5650,17'd5965,17'd6271,17'd9962,17'd7715,17'd6897,17'd6897,17'd11732,17'd11447,17'd9128,17'd9268,17'd9129,17'd8665,17'd11200,17'd8982,17'd6432,17'd10084,17'd9966,17'd8669,17'd6104,17'd6432,17'd6592,17'd11885,17'd10921,17'd11886,17'd11887,17'd2781,17'd2936,17'd2597,17'd10670,17'd11888,17'd471,17'd471,17'd294,17'd293,17'd1834,17'd1834,17'd3431,17'd11208,17'd3756,17'd3756,17'd5656,17'd11889,17'd11737,17'd11890,17'd5976,17'd11891,17'd11892,17'd5063,17'd11893,17'd11894,17'd6756,17'd11895,17'd11896,17'd9826,17'd11897,17'd11217,17'd11898,17'd11899,17'd11900,17'd11901,17'd11749,17'd11750,17'd11902,17'd11903,17'd11904,17'd11905,17'd11906,17'd11907,17'd11908,17'd11909,17'd11910,17'd11911,17'd11759,17'd11761,17'd11762,17'd11762,17'd11912,17'd10940,17'd11086,17'd11626,17'd11763,17'd11478,17'd11913,17'd11914,17'd10815,17'd10815,17'd11087,17'd11915,17'd10944,17'd10943,17'd10564,17'd10817,17'd10817,17'd10817,17'd11232,17'd9006,17'd8537,17'd5409,17'd5837,17'd5837,17'd5255,17'd4927,17'd9302,17'd4927,17'd6626,17'd6626,17'd8370,17'd8370,17'd6468,17'd6769,17'd7086,17'd8218,17'd8065,17'd11916,17'd11765,17'd11235,17'd11482,17'd11917,17'd11483,17'd11483,17'd11918,17'd11919,17'd11094,17'd11238,17'd11095,17'd10818,17'd11920,17'd7590,17'd10702,17'd11240,17'd11921,17'd11922,17'd11923,17'd9996,17'd10705,17'd11486,17'd11635,17'd11924,17'd11925,17'd11926,17'd11638,17'd11927,17'd11777,17'd11778,17'd11778,17'd11928,17'd11780,17'd11929,17'd11930,17'd11931,17'd11932,17'd11933,17'd11934,17'd11935,17'd11936,17'd11937,17'd11650,17'd11650,17'd11938,17'd11939,17'd11940,17'd11941,17'd11942,17'd11943,17'd11944,17'd11945,17'd11946,17'd11946,17'd11947,17'd11948,17'd11949,17'd11385,17'd11950,17'd11951,17'd11952,17'd11953,17'd11954,17'd11955,17'd11956,17'd11957,17'd11958,17'd11959,17'd11959,17'd11960,17'd11961,17'd11806,17'd11962,17'd11962,17'd11963,17'd11964,17'd11965,17'd10990,17'd10739,17'd11133,17'd11134,17'd11277,17'd11809,17'd9344,17'd8873,17'd8881,17'd10027,17'd11966,17'd11967,17'd11812,17'd11968,17'd8257,17'd11969,17'd11970,17'd8265,17'd11971,17'd11972,17'd11973,17'd11974,17'd11975,17'd11976,17'd10037,17'd11977,17'd8444,17'd11289,17'd11413,17'd7980,17'd7980,17'd1045,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd131,17'd11978,17'd3660,17'd11979,17'd11980,17'd11981,17'd11982,17'd10765,17'd11983,17'd9215,17'd11984,17'd11985,17'd11986,17'd9505,17'd10201,17'd11987,17'd11162,17'd10767,17'd11988,17'd11832,17'd11989,17'd11990,17'd11991,17'd9228,17'd10502,17'd10888,17'd11833,17'd11833,17'd11992,17'd11993,17'd11994,17'd11995,17'd11699,17'd11996,17'd11836,17'd11836,17'd8777,17'd11997,17'd11997,17'd11997,17'd11998,17'd11998,17'd11998,17'd11837,17'd11837,17'd11837,17'd11836,17'd11426,17'd11700,17'd11024,17'd10219,17'd9928,17'd11029,17'd11565,17'd11839,17'd11839,17'd11565,17'd11566,17'd11704,17'd11840,17'd11999,17'd11999,17'd12000,17'd12001,17'd12001,17'd11843,17'd11844,17'd11845,17'd11846,17'd11846,17'd10510,17'd11309,17'd11705,17'd11705,17'd10226,17'd9780,17'd10063,17'd11310,17'd9651,17'd10228,17'd12002,17'd11176,17'd11849,17'd11849,17'd11850,17'd11851,17'd12003,17'd11851,17'd11572,17'd12004,17'd12004,17'd11572,17'd11313,17'd11852,17'd11853,17'd11853,17'd11576,17'd11576,17'd11432,17'd11855,17'd11855,17'd12005,17'd10779,17'd8002,17'd8472,17'd8472,17'd6561,17'd7330,17'd7183,17'd12006,17'd12007,17'd12008,17'd12009,17'd12010,17'd12011,17'd12012,17'd12013,17'd12014,17'd12015,17'd12016,17'd11720,17'd11868,17'd11869,17'd3247,17'd5788,17'd11591,17'd12017,17'd3887,17'd5368,17'd6874,17'd4568,17'd7689,17'd7029,17'd7858,17'd9252,17'd9252,17'd8491,17'd8795,17'd11191,17'd11191,17'd12018,17'd12019,17'd9110,17'd12020,17'd12021,17'd11724,17'd9256,17'd9538,17'd11331,17'd12022,17'd12023,17'd12024,17'd8804,17'd9409,17'd9408,17'd11052,17'd9538,17'd9539,17'd9951,17'd8649,17'd8650,17'd7690,17'd9411,17'd8499,17'd11876,17'd11877,17'd12025,17'd11878,17'd7867,17'd8809,17'd9799,17'd9799,17'd9955,17'd8181,17'd7698,17'd8181,17'd9956,17'd11332,17'd8656,17'd10530,17'd9958,17'd9544,17'd11061,17'd11061,17'd11061,17'd11061,17'd11336,17'd11335,17'd4714,17'd9123,17'd5940,17'd5940,17'd12026,17'd421,17'd418,17'd1951,17'd12027,17'd12028
},
'{
17'd0,17'd0,17'd1,17'd1,17'd3,17'd12,17'd0,17'd2,17'd14,17'd1967,17'd5196,17'd7711,17'd7545,17'd7545,17'd12029,17'd4886,17'd466,17'd3,17'd465,17'd2421,17'd6,17'd5205,17'd8040,17'd8040,17'd8190,17'd8190,17'd8190,17'd8190,17'd8340,17'd8340,17'd8339,17'd8340,17'd7727,17'd8520,17'd9136,17'd10263,17'd7055,17'd6592,17'd12030,17'd12031,17'd12032,17'd8665,17'd9131,17'd8817,17'd7887,17'd7550,17'd10399,17'd11605,17'd10263,17'd10920,17'd9137,17'd6105,17'd9420,17'd10663,17'd12033,17'd8043,17'd12034,17'd12035,17'd6265,17'd1967,17'd2257,17'd2426,17'd10802,17'd11888,17'd471,17'd471,17'd34,17'd2427,17'd12036,17'd12036,17'd3431,17'd3754,17'd3910,17'd3910,17'd5804,17'd11737,17'd12037,17'd12037,17'd5975,17'd12038,17'd12039,17'd12040,17'd5390,17'd12041,17'd12042,17'd12043,17'd12044,17'd12045,17'd11461,17'd12046,17'd12047,17'd11748,17'd12048,17'd12049,17'd12050,17'd12051,17'd11751,17'd12052,17'd12053,17'd12054,17'd12055,17'd12056,17'd12057,17'd12058,17'd12059,17'd12060,17'd12061,17'd10937,17'd12062,17'd11761,17'd12063,17'd12064,17'd11476,17'd12065,17'd11763,17'd11478,17'd12066,17'd11914,17'd10815,17'd10816,17'd11087,17'd11087,17'd10564,17'd10564,17'd10817,17'd10817,17'd10286,17'd10564,17'd11232,17'd8537,17'd7418,17'd5409,17'd5409,17'd5255,17'd4927,17'd4927,17'd4927,17'd4927,17'd4927,17'd4927,17'd8370,17'd6468,17'd6142,17'd8368,17'd8218,17'd7414,17'd9570,17'd12067,17'd12068,17'd11766,17'd11917,17'd11917,17'd12069,17'd12069,17'd11918,17'd11484,17'd11094,17'd12070,17'd9311,17'd10818,17'd12071,17'd7590,17'd10435,17'd12072,17'd12073,17'd12074,17'd12075,17'd9855,17'd11486,17'd11487,17'd12076,17'd12077,17'd12078,17'd11491,17'd12079,17'd12080,17'd11778,17'd12081,17'd11778,17'd11928,17'd11780,17'd11929,17'd12082,17'd12083,17'd12084,17'd12085,17'd12086,17'd12087,17'd12088,17'd12089,17'd11649,17'd12090,17'd12091,17'd12092,17'd12093,17'd12094,17'd12095,17'd12096,17'd12097,17'd12097,17'd12097,17'd12098,17'd12099,17'd11948,17'd11794,17'd11655,17'd12100,17'd11952,17'd12101,17'd12102,17'd12103,17'd12104,17'd12105,17'd12106,17'd12107,17'd12107,17'd12108,17'd12109,17'd12110,17'd12111,17'd12112,17'd12112,17'd12113,17'd12114,17'd12115,17'd10989,17'd10988,17'd10740,17'd11134,17'd12116,17'd9479,17'd12117,17'd9188,17'd12118,17'd8726,17'd11966,17'd11967,17'd12119,17'd12120,17'd9351,17'd9891,17'd12121,17'd12122,17'd12123,17'd12124,17'd12125,17'd11681,17'd11287,17'd11976,17'd12126,17'd11977,17'd8444,17'd11289,17'd8132,17'd888,17'd7980,17'd1045,17'd1197,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd131,17'd12127,17'd5747,17'd12128,17'd12129,17'd12130,17'd12131,17'd12132,17'd12133,17'd12134,17'd12135,17'd12136,17'd11986,17'd9505,17'd12137,17'd12138,17'd12139,17'd11297,17'd12140,17'd8616,17'd12141,17'd12142,17'd11553,17'd11300,17'd10888,17'd10888,17'd12143,17'd12144,17'd8617,17'd9648,17'd12145,17'd9650,17'd11998,17'd11167,17'd11997,17'd11998,17'd12146,17'd12147,17'd12147,17'd12148,17'd12148,17'd12148,17'd12148,17'd12148,17'd12148,17'd12149,17'd11997,17'd11167,17'd12150,17'd12151,17'd12152,17'd9516,17'd9928,17'd10064,17'd11839,17'd11839,17'd11839,17'd12153,17'd11704,17'd11840,17'd11999,17'd11999,17'd12154,17'd12154,17'd12000,17'd12000,17'd12001,17'd11843,17'd11844,17'd11845,17'd11845,17'd11845,17'd11309,17'd11705,17'd12155,17'd12155,17'd10227,17'd9517,17'd9384,17'd9651,17'd12156,17'd12157,17'd12003,17'd11850,17'd11850,17'd12003,17'd12158,17'd12003,17'd12003,17'd12159,17'd12004,17'd12004,17'd11314,17'd11314,17'd11852,17'd11852,17'd11576,17'd10641,17'd12160,17'd12161,17'd12162,17'd12163,17'd12164,17'd12165,17'd6558,17'd6559,17'd11040,17'd6712,17'd7016,17'd12006,17'd12166,17'd12167,17'd12009,17'd12168,17'd12169,17'd12170,17'd12171,17'd12172,17'd12173,17'd12174,17'd12175,17'd12176,17'd11869,17'd1810,17'd2922,17'd12177,17'd3088,17'd3583,17'd3727,17'd2755,17'd6248,17'd7518,17'd6873,17'd7686,17'd9252,17'd9252,17'd8170,17'd8795,17'd11191,17'd11191,17'd12018,17'd12019,17'd11723,17'd12178,17'd12021,17'd11873,17'd11724,17'd11595,17'd8800,17'd11331,17'd12023,17'd12023,17'd9950,17'd8495,17'd9115,17'd11052,17'd9538,17'd9538,17'd9665,17'd8648,17'd12179,17'd7690,17'd7864,17'd12180,17'd11876,17'd12181,17'd11877,17'd11878,17'd8809,17'd8809,17'd9799,17'd10256,17'd9956,17'd9120,17'd7698,17'd7698,17'd9120,17'd12182,17'd11196,17'd12183,17'd12184,17'd9544,17'd11061,17'd11061,17'd11061,17'd11061,17'd11061,17'd11336,17'd4714,17'd9123,17'd5940,17'd2393,17'd11445,17'd421,17'd418,17'd1951,17'd12027,17'd11884
},
'{
17'd0,17'd0,17'd1,17'd1,17'd3,17'd12,17'd2,17'd14,17'd1689,17'd3750,17'd6096,17'd7711,17'd7545,17'd5508,17'd7214,17'd6419,17'd13,17'd1275,17'd2591,17'd2421,17'd6,17'd5205,17'd8190,17'd8040,17'd8340,17'd8190,17'd8190,17'd8340,17'd8340,17'd8340,17'd8340,17'd8190,17'd7375,17'd12185,17'd9137,17'd6271,17'd6741,17'd8342,17'd12186,17'd12187,17'd12188,17'd10262,17'd12189,17'd8978,17'd9264,17'd7054,17'd6899,17'd10917,17'd12190,17'd9420,17'd6105,17'd6595,17'd11199,17'd10665,17'd12191,17'd8191,17'd12192,17'd12193,17'd2781,17'd3249,17'd12194,17'd12195,17'd11072,17'd12196,17'd471,17'd294,17'd2119,17'd12197,17'd12198,17'd12036,17'd3431,17'd11210,17'd6278,17'd5804,17'd6110,17'd5976,17'd12037,17'd12199,17'd12200,17'd4898,17'd12201,17'd4099,17'd5391,17'd12202,17'd6758,17'd12203,17'd10552,17'd12204,17'd12205,17'd11463,17'd11901,17'd12206,17'd12050,17'd12207,17'd12207,17'd12051,17'd11752,17'd12053,17'd12208,17'd12209,17'd12210,17'd12211,17'd12212,17'd12059,17'd12213,17'd12060,17'd12214,17'd12215,17'd10937,17'd11761,17'd12063,17'd12216,17'd12217,17'd12218,17'd11627,17'd11913,17'd12066,17'd10815,17'd10427,17'd11087,17'd11087,17'd11087,17'd10564,17'd10817,17'd10817,17'd10817,17'd10112,17'd11232,17'd12219,17'd5409,17'd5837,17'd5409,17'd4927,17'd4927,17'd4927,17'd4927,17'd5255,17'd4927,17'd9302,17'd10430,17'd6468,17'd6142,17'd6142,17'd12220,17'd7414,17'd8065,17'd11916,17'd11765,17'd11766,17'd11482,17'd11917,17'd11917,17'd12069,17'd11918,17'd11919,17'd11094,17'd12070,17'd9311,17'd10818,17'd9166,17'd7923,17'd7925,17'd12221,17'd12222,17'd12223,17'd12224,17'd11098,17'd11367,17'd12225,17'd11487,17'd11924,17'd12226,17'd12227,17'd11638,17'd11639,17'd11640,17'd12228,17'd12081,17'd11778,17'd11779,17'd12229,17'd12230,17'd12231,17'd12232,17'd12233,17'd12234,17'd12235,17'd12236,17'd12088,17'd12237,17'd12238,17'd12239,17'd12240,17'd12241,17'd12242,17'd12243,17'd12094,17'd12095,17'd12244,17'd12244,17'd12244,17'd12096,17'd12245,17'd12246,17'd11795,17'd12247,17'd11801,17'd11268,17'd12248,17'd12249,17'd12250,17'd12251,17'd12252,17'd12253,17'd12254,17'd12255,17'd12108,17'd12253,17'd12256,17'd12257,17'd12258,17'd12258,17'd12259,17'd12260,17'd12261,17'd12262,17'd10737,17'd10475,17'd10330,17'd9741,17'd9480,17'd10174,17'd12263,17'd12264,17'd8412,17'd8412,17'd11967,17'd12119,17'd12265,17'd12266,17'd9891,17'd12267,17'd12268,17'd12269,17'd12270,17'd12271,17'd12272,17'd11412,17'd11976,17'd12273,17'd12274,17'd12275,17'd11152,17'd10874,17'd7980,17'd7980,17'd1045,17'd1197,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd6369,17'd4500,17'd12276,17'd3822,17'd12277,17'd12278,17'd6699,17'd12279,17'd12280,17'd11984,17'd12281,17'd11160,17'd9640,17'd12282,17'd12283,17'd12284,17'd12285,17'd8617,17'd8618,17'd9513,17'd12286,17'd11696,17'd9227,17'd10888,17'd11425,17'd12287,17'd12288,17'd8767,17'd9648,17'd11835,17'd12148,17'd12149,17'd12149,17'd9650,17'd8464,17'd8464,17'd8464,17'd9379,17'd8151,17'd8151,17'd12289,17'd12289,17'd12290,17'd12146,17'd11998,17'd11837,17'd12291,17'd12291,17'd12292,17'd10061,17'd10060,17'd10220,17'd10376,17'd10509,17'd11839,17'd12293,17'd11704,17'd11566,17'd11566,17'd11841,17'd12294,17'd12295,17'd12154,17'd12154,17'd12154,17'd12000,17'd12001,17'd11843,17'd11843,17'd12001,17'd11844,17'd11309,17'd12155,17'd12296,17'd12297,17'd11705,17'd11705,17'd11309,17'd10226,17'd12298,17'd12299,17'd12300,17'd12301,17'd12301,17'd12158,17'd12158,17'd12158,17'd12302,17'd12158,17'd12303,17'd12304,17'd12305,17'd11313,17'd11852,17'd12306,17'd11853,17'd10641,17'd11576,17'd12307,17'd12162,17'd12162,17'd12308,17'd12309,17'd8471,17'd6559,17'd7501,17'd8156,17'd11433,17'd7332,17'd12310,17'd12166,17'd12167,17'd12168,17'd12311,17'd12312,17'd12313,17'd12314,17'd12315,17'd12316,17'd12317,17'd12318,17'd5028,17'd2240,17'd6885,17'd5192,17'd11591,17'd3237,17'd3886,17'd6578,17'd4409,17'd6577,17'd7030,17'd7686,17'd8171,17'd9252,17'd8170,17'd8795,17'd11050,17'd11191,17'd10076,17'd12319,17'd12320,17'd11723,17'd12020,17'd12021,17'd11873,17'd11874,17'd9538,17'd9408,17'd12321,17'd12321,17'd11331,17'd8495,17'd9114,17'd9408,17'd9538,17'd9949,17'd11053,17'd9540,17'd8649,17'd7690,17'd7690,17'd7864,17'd8652,17'd12181,17'd12181,17'd11878,17'd8809,17'd8809,17'd9799,17'd10256,17'd10256,17'd9956,17'd8181,17'd12322,17'd12322,17'd12182,17'd12323,17'd12324,17'd12325,17'd9670,17'd2906,17'd11061,17'd11882,17'd11061,17'd11061,17'd11336,17'd4714,17'd9123,17'd5940,17'd5630,17'd11600,17'd1669,17'd417,17'd2102,17'd11601,17'd12326
},
'{
17'd15,17'd15,17'd1,17'd1,17'd3,17'd12,17'd2590,17'd6419,17'd5196,17'd7711,17'd7545,17'd5508,17'd3252,17'd1831,17'd4247,17'd466,17'd8814,17'd22,17'd4,17'd6,17'd6,17'd3753,17'd5205,17'd8040,17'd8040,17'd8339,17'd8339,17'd8340,17'd8340,17'd5205,17'd5205,17'd5206,17'd11730,17'd9136,17'd9420,17'd10920,17'd10541,17'd9681,17'd8341,17'd8342,17'd7720,17'd7548,17'd9264,17'd7549,17'd6898,17'd7056,17'd9133,17'd12327,17'd12328,17'd9136,17'd8669,17'd6271,17'd11069,17'd12329,17'd12330,17'd12331,17'd12332,17'd3750,17'd1688,17'd1831,17'd10669,17'd10924,17'd11888,17'd11888,17'd32,17'd292,17'd470,17'd12197,17'd12197,17'd12333,17'd12334,17'd12335,17'd12336,17'd6110,17'd12337,17'd5384,17'd12038,17'd4899,17'd12338,17'd12339,17'd3270,17'd12340,17'd4905,17'd12341,17'd12342,17'd12343,17'd11218,17'd12344,17'd11618,17'd12345,17'd12346,17'd12347,17'd12050,17'd12049,17'd11749,17'd11750,17'd12052,17'd12348,17'd12349,17'd12350,17'd12351,17'd12352,17'd12353,17'd12213,17'd12059,17'd12354,17'd12355,17'd12356,17'd12062,17'd12357,17'd12358,17'd12359,17'd12360,17'd12361,17'd12362,17'd12362,17'd11913,17'd11629,17'd10563,17'd10563,17'd10692,17'd10692,17'd10564,17'd10817,17'd10817,17'd10817,17'd10817,17'd11232,17'd6468,17'd6140,17'd6140,17'd6626,17'd4927,17'd9302,17'd8538,17'd7582,17'd8538,17'd10430,17'd10430,17'd12219,17'd12220,17'd8536,17'd7086,17'd7414,17'd12363,17'd11234,17'd12364,17'd12365,17'd12366,17'd12367,17'd12368,17'd12369,17'd11918,17'd11919,17'd11094,17'd9310,17'd9311,17'd9019,17'd12370,17'd12371,17'd12372,17'd12373,17'd12374,17'd12375,17'd12376,17'd12377,17'd12378,17'd12379,17'd12380,17'd11635,17'd11773,17'd12381,17'd12382,17'd12383,17'd11927,17'd11640,17'd12384,17'd12385,17'd12386,17'd12387,17'd12388,17'd12389,17'd12390,17'd12391,17'd12392,17'd12393,17'd12087,17'd12394,17'd12395,17'd11647,17'd12396,17'd12397,17'd12398,17'd12399,17'd12400,17'd12242,17'd12401,17'd12402,17'd12245,17'd12403,17'd12404,17'd12405,17'd12406,17'd12407,17'd11799,17'd12247,17'd11389,17'd12408,17'd12409,17'd12410,17'd12411,17'd12412,17'd12413,17'd12414,17'd12253,17'd12253,17'd12415,17'd12416,17'd12417,17'd12418,17'd12414,17'd12109,17'd12419,17'd12420,17'd12421,17'd12422,17'd11808,17'd12423,17'd10330,17'd10024,17'd9620,17'd8874,17'd8877,17'd12424,17'd12425,17'd9886,17'd11811,17'd12426,17'd12427,17'd12428,17'd12429,17'd12430,17'd10612,17'd12431,17'd12432,17'd11409,17'd12433,17'd11974,17'd11288,17'd12434,17'd12435,17'd7812,17'd7813,17'd8132,17'd889,17'd1045,17'd11413,17'd1045,17'd1045,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd135,17'd357,17'd6199,17'd12436,17'd12437,17'd12438,17'd12439,17'd12440,17'd11420,17'd12441,17'd12442,17'd12443,17'd12444,17'd12445,17'd9222,17'd12446,17'd12447,17'd12447,17'd9078,17'd9920,17'd9921,17'd12448,17'd11992,17'd9644,17'd9376,17'd9375,17'd9224,17'd12288,17'd11834,17'd12449,17'd12449,17'd11994,17'd12145,17'd12450,17'd12451,17'd12451,17'd12451,17'd12452,17'd12452,17'd12147,17'd12147,17'd12147,17'd12146,17'd11998,17'd12291,17'd12453,17'd12453,17'd12453,17'd12454,17'd12454,17'd12455,17'd12456,17'd12457,17'd12152,17'd12152,17'd10219,17'd10064,17'd11565,17'd11704,17'd11566,17'd11307,17'd12458,17'd11842,17'd11999,17'd12294,17'd12459,17'd12459,17'd12460,17'd12154,17'd12001,17'd11844,17'd12000,17'd11845,17'd11846,17'd11844,17'd12001,17'd12001,17'd12001,17'd12000,17'd12000,17'd11705,17'd11309,17'd10226,17'd10221,17'd12461,17'd12462,17'd11567,17'd12300,17'd12300,17'd12300,17'd12300,17'd12300,17'd12303,17'd12303,17'd11571,17'd12463,17'd12464,17'd11852,17'd12465,17'd12466,17'd12465,17'd12467,17'd12468,17'd12469,17'd12470,17'd12471,17'd6709,17'd6710,17'd6856,17'd8634,17'd7672,17'd12006,17'd12472,17'd12473,17'd12474,17'd12475,17'd12476,17'd12477,17'd12478,17'd12479,17'd12480,17'd12481,17'd12482,17'd12483,17'd12484,17'd12485,17'd2096,17'd6886,17'd7363,17'd3580,17'd12486,17'd2569,17'd6244,17'd6576,17'd7346,17'd8169,17'd7856,17'd8170,17'd8491,17'd8491,17'd8795,17'd10076,17'd11592,17'd12487,17'd12488,17'd12489,17'd12178,17'd11873,17'd11874,17'd11595,17'd9949,17'd8646,17'd8646,17'd11331,17'd9950,17'd9540,17'd9665,17'd9539,17'd9539,17'd9795,17'd11054,17'd8962,17'd7690,17'd8324,17'd8324,17'd9411,17'd9542,17'd8027,17'd8027,17'd8326,17'd8809,17'd8809,17'd9799,17'd9799,17'd9955,17'd12322,17'd12490,17'd12491,17'd12492,17'd11597,17'd12493,17'd9802,17'd12494,17'd4559,17'd12495,17'd11882,17'd11061,17'd11061,17'd11336,17'd4714,17'd5183,17'd5630,17'd12496,17'd414,17'd421,17'd417,17'd2104,17'd12497,17'd12498
},
'{
17'd15,17'd15,17'd0,17'd0,17'd12,17'd13,17'd2590,17'd6419,17'd6583,17'd7711,17'd4887,17'd4887,17'd2422,17'd4247,17'd466,17'd13,17'd22,17'd24,17'd5,17'd6,17'd7,17'd7,17'd5205,17'd8040,17'd8339,17'd8339,17'd8339,17'd8340,17'd8190,17'd7374,17'd10536,17'd5513,17'd6732,17'd8511,17'd7222,17'd9682,17'd11341,17'd11341,17'd8984,17'd10399,17'd7889,17'd7550,17'd7889,17'd7715,17'd6741,17'd8984,17'd10917,17'd12499,17'd8670,17'd8042,17'd9272,17'd7546,17'd12500,17'd12501,17'd12329,17'd12502,17'd12503,17'd1689,17'd1831,17'd3252,17'd11071,17'd11888,17'd12504,17'd12505,17'd32,17'd982,17'd470,17'd2427,17'd12197,17'd12333,17'd12506,17'd5658,17'd12507,17'd11737,17'd11738,17'd11891,17'd4899,17'd12508,17'd12509,17'd3604,17'd3606,17'd12510,17'd12511,17'd12512,17'd12513,17'd9288,17'd12514,17'd12515,17'd12345,17'd12516,17'd12346,17'd11750,17'd12517,17'd12347,17'd12347,17'd12518,17'd12519,17'd12520,17'd12521,17'd12522,17'd12523,17'd12524,17'd12060,17'd12525,17'd12354,17'd12526,17'd11084,17'd12062,17'd12062,17'd12527,17'd12528,17'd12529,17'd12530,17'd12362,17'd12362,17'd12362,17'd12531,17'd12532,17'd11362,17'd10563,17'd10692,17'd10817,17'd12533,17'd10817,17'd10564,17'd10564,17'd10564,17'd9158,17'd6468,17'd6626,17'd6626,17'd4927,17'd4927,17'd9302,17'd8538,17'd8538,17'd9007,17'd12534,17'd9006,17'd12219,17'd12535,17'd8536,17'd8218,17'd8065,17'd12536,17'd12537,17'd12365,17'd12366,17'd12367,17'd12538,17'd12368,17'd12369,17'd11918,17'd11093,17'd9310,17'd9165,17'd12370,17'd12071,17'd12071,17'd8857,17'd12539,17'd12540,17'd12541,17'd12542,17'd12543,17'd12544,17'd12545,17'd12546,17'd12547,17'd12548,17'd12549,17'd12550,17'd11244,17'd12080,17'd11776,17'd12551,17'd11777,17'd11372,17'd12552,17'd12553,17'd12554,17'd12555,17'd12556,17'd12557,17'd12558,17'd12559,17'd12560,17'd12395,17'd12561,17'd12562,17'd12563,17'd12564,17'd12565,17'd12566,17'd12567,17'd12568,17'd12569,17'd12570,17'd12571,17'd12245,17'd12572,17'd12406,17'd12406,17'd12572,17'd11949,17'd11510,17'd11264,17'd12573,17'd12574,17'd12575,17'd12576,17'd12576,17'd12577,17'd12577,17'd12414,17'd12578,17'd12418,17'd12416,17'd12416,17'd12416,17'd12253,17'd12579,17'd12580,17'd12419,17'd12581,17'd12582,17'd12583,17'd12584,17'd12585,17'd10024,17'd9620,17'd9038,17'd8723,17'd8728,17'd11404,17'd12586,17'd12587,17'd12588,17'd12589,17'd12590,17'd12591,17'd12592,17'd12593,17'd12594,17'd12595,17'd12596,17'd12597,17'd11974,17'd11975,17'd10036,17'd10620,17'd9756,17'd10873,17'd10874,17'd11413,17'd1197,17'd11413,17'd1045,17'd1045,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd134,17'd2861,17'd4816,17'd12598,17'd12599,17'd12600,17'd6697,17'd10765,17'd12601,17'd12602,17'd12603,17'd11692,17'd11160,17'd12604,17'd12605,17'd12446,17'd9078,17'd9230,17'd8770,17'd10053,17'd10053,17'd12606,17'd11020,17'd12607,17'd10205,17'd9224,17'd12608,17'd8920,17'd12609,17'd12610,17'd12610,17'd11994,17'd11994,17'd12611,17'd12611,17'd12611,17'd12145,17'd12452,17'd9650,17'd12147,17'd12146,17'd12146,17'd12612,17'd12291,17'd12453,17'd12455,17'd12455,17'd12613,17'd12613,17'd12455,17'd12455,17'd12613,17'd12456,17'd12152,17'd9779,17'd12614,17'd10219,17'd11027,17'd11565,17'd12458,17'd11842,17'd11842,17'd11841,17'd11841,17'd11999,17'd12615,17'd12459,17'd12460,17'd12295,17'd12154,17'd12000,17'd11844,17'd11843,17'd11843,17'd11844,17'd12616,17'd12617,17'd12618,17'd12618,17'd12001,17'd11843,17'd12297,17'd12296,17'd11309,17'd10222,17'd12619,17'd12620,17'd12300,17'd12157,17'd12157,17'd12157,17'd12157,17'd12621,17'd12304,17'd12303,17'd12463,17'd12464,17'd11852,17'd11852,17'd12465,17'd12465,17'd11854,17'd12622,17'd12623,17'd11855,17'd12624,17'd12625,17'd7501,17'd7838,17'd7330,17'd11433,17'd12626,17'd12006,17'd12473,17'd12627,17'd12475,17'd12628,17'd12629,17'd12630,17'd12631,17'd12632,17'd12633,17'd12634,17'd12635,17'd12483,17'd12636,17'd12485,17'd12637,17'd7704,17'd12638,17'd3085,17'd12639,17'd6245,17'd4718,17'd9116,17'd7685,17'd8169,17'd8018,17'd8170,17'd8491,17'd8795,17'd10076,17'd12018,17'd10077,17'd12487,17'd11723,17'd12178,17'd11873,17'd11724,17'd12640,17'd11192,17'd9796,17'd8646,17'd8646,17'd11331,17'd9665,17'd9665,17'd9539,17'd9949,17'd9795,17'd11725,17'd9666,17'd8650,17'd8324,17'd8324,17'd8324,17'd8324,17'd12641,17'd8027,17'd9259,17'd7867,17'd8809,17'd8809,17'd9955,17'd9955,17'd9956,17'd12322,17'd12642,17'd12492,17'd11597,17'd11597,17'd11333,17'd12643,17'd9670,17'd2906,17'd11882,17'd11882,17'd11061,17'd11336,17'd5183,17'd4714,17'd5940,17'd5940,17'd12496,17'd12644,17'd2560,17'd12645,17'd2395,17'd12646
},
'{
17'd15,17'd15,17'd0,17'd0,17'd13,17'd13,17'd12647,17'd6419,17'd6583,17'd4577,17'd2784,17'd2422,17'd1831,17'd1127,17'd0,17'd806,17'd23,17'd5,17'd6,17'd7,17'd5205,17'd8190,17'd8340,17'd8340,17'd8339,17'd8339,17'd8340,17'd8340,17'd5205,17'd10536,17'd12648,17'd12649,17'd8670,17'd7057,17'd7222,17'd9137,17'd12650,17'd12651,17'd10666,17'd10399,17'd7055,17'd7715,17'd7715,17'd6431,17'd10401,17'd9133,17'd7222,17'd8824,17'd6596,17'd6434,17'd10263,17'd7051,17'd12034,17'd7721,17'd6590,17'd12652,17'd2781,17'd1688,17'd3252,17'd3101,17'd10925,17'd11888,17'd12653,17'd12196,17'd293,17'd2943,17'd12654,17'd12654,17'd12654,17'd3258,17'd12335,17'd12655,17'd6110,17'd5976,17'd12656,17'd12657,17'd12508,17'd12658,17'd3441,17'd12659,17'd12660,17'd12661,17'd12662,17'd12663,17'd9150,17'd9829,17'd12664,17'd12665,17'd12666,17'd12667,17'd12051,17'd12517,17'd12668,17'd12669,17'd12670,17'd12671,17'd12054,17'd12672,17'd12673,17'd11908,17'd12674,17'd12675,17'd12059,17'd12525,17'd12676,17'd12526,17'd10937,17'd12677,17'd12678,17'd12679,17'd12529,17'd12360,17'd12218,17'd12362,17'd12680,17'd11913,17'd12532,17'd12681,17'd11362,17'd11362,17'd10427,17'd10691,17'd12533,17'd10817,17'd11232,17'd12682,17'd9158,17'd8369,17'd5837,17'd5255,17'd4927,17'd9302,17'd10430,17'd8538,17'd9007,17'd9007,17'd10694,17'd10694,17'd12219,17'd12219,17'd8687,17'd8218,17'd8686,17'd9569,17'd12683,17'd12684,17'd12367,17'd12538,17'd12538,17'd12368,17'd12368,17'd12369,17'd11918,17'd11093,17'd9444,17'd9165,17'd12685,17'd12686,17'd8855,17'd10702,17'd9023,17'd9173,17'd11769,17'd12687,17'd12688,17'd12379,17'd12546,17'd12546,17'd12689,17'd12077,17'd12690,17'd12691,17'd12692,17'd12693,17'd12694,17'd12694,17'd12695,17'd11928,17'd12387,17'd12696,17'd11781,17'd12697,17'd12698,17'd12699,17'd12235,17'd12700,17'd12701,17'd12702,17'd12703,17'd12704,17'd12705,17'd12706,17'd12707,17'd12708,17'd12709,17'd12568,17'd12569,17'd12710,17'd12711,17'd12712,17'd12407,17'd12403,17'd12245,17'd12099,17'd12713,17'd12714,17'd12715,17'd12716,17'd12717,17'd12575,17'd12577,17'd12577,17'd12718,17'd12420,17'd12109,17'd12578,17'd12418,17'd12418,17'd12415,17'd12416,17'd12253,17'd12109,17'd12110,17'd12110,17'd12719,17'd11962,17'd12720,17'd12721,17'd11401,17'd12116,17'd9344,17'd9188,17'd12722,17'd12723,17'd12724,17'd12725,17'd10339,17'd8580,17'd12726,17'd12727,17'd12728,17'd12729,17'd10612,17'd12730,17'd12731,17'd12732,17'd12733,17'd11974,17'd11287,17'd10872,17'd10037,17'd11977,17'd12275,17'd11152,17'd11413,17'd1045,17'd11413,17'd1045,17'd1045,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd10492,17'd12734,17'd9362,17'd12735,17'd12736,17'd12737,17'd8450,17'd12738,17'd12739,17'd12740,17'd12741,17'd12742,17'd9070,17'd12743,17'd12744,17'd12745,17'd12746,17'd8923,17'd12747,17'd12748,17'd12749,17'd9772,17'd12750,17'd10205,17'd11425,17'd11695,17'd8920,17'd11993,17'd11994,17'd12450,17'd12611,17'd12611,17'd12611,17'd12611,17'd12452,17'd12452,17'd8151,17'd9650,17'd12147,17'd12146,17'd12751,17'd12291,17'd9520,17'd12752,17'd12455,17'd12455,17'd12753,17'd12753,17'd12754,17'd12754,17'd12455,17'd12613,17'd12457,17'd10062,17'd12755,17'd11310,17'd11025,17'd10893,17'd11428,17'd12458,17'd11842,17'd11841,17'd11841,17'd11841,17'd12756,17'd12757,17'd12460,17'd12460,17'd12460,17'd12460,17'd11843,17'd12001,17'd12001,17'd11844,17'd11845,17'd11843,17'd12618,17'd12617,17'd12001,17'd12001,17'd12000,17'd12295,17'd12757,17'd11705,17'd10221,17'd12619,17'd12002,17'd11706,17'd12621,17'd12157,17'd12621,17'd12758,17'd12759,17'd12759,17'd12305,17'd12305,17'd11852,17'd12306,17'd11852,17'd11314,17'd11853,17'd12760,17'd12761,17'd12469,17'd12762,17'd12763,17'd7501,17'd7838,17'd6856,17'd8634,17'd12626,17'd12006,17'd12473,17'd12627,17'd12764,17'd12765,17'd12766,17'd12767,17'd12768,17'd12769,17'd12770,17'd12771,17'd12772,17'd12773,17'd5373,17'd4575,17'd4422,17'd6887,17'd3087,17'd12774,17'd12775,17'd5037,17'd4719,17'd4871,17'd6724,17'd7685,17'd8169,17'd7856,17'd8170,17'd8491,17'd10076,17'd11722,17'd11593,17'd12487,17'd11723,17'd12178,17'd12021,17'd11873,17'd12776,17'd11874,17'd8957,17'd8646,17'd8799,17'd8799,17'd9539,17'd8801,17'd9539,17'd9256,17'd9795,17'd12777,17'd11725,17'd9541,17'd12778,17'd8324,17'd8324,17'd9411,17'd8652,17'd8652,17'd8027,17'd8326,17'd8809,17'd8809,17'd9955,17'd9955,17'd10256,17'd9120,17'd12642,17'd12642,17'd8655,17'd11597,17'd11196,17'd12779,17'd12780,17'd5183,17'd11336,17'd11882,17'd11061,17'd11336,17'd5183,17'd9123,17'd3073,17'd2393,17'd2589,17'd1529,17'd418,17'd2103,17'd12498,17'd12646
},
'{
17'd15,17'd15,17'd0,17'd0,17'd13,17'd2,17'd6419,17'd5196,17'd7711,17'd4577,17'd2784,17'd2422,17'd1688,17'd14,17'd3,17'd1275,17'd4,17'd5,17'd7,17'd7,17'd8190,17'd8190,17'd8340,17'd8340,17'd8339,17'd8339,17'd8340,17'd5205,17'd7,17'd7216,17'd12781,17'd12782,17'd6900,17'd9682,17'd8824,17'd8518,17'd12650,17'd9681,17'd6741,17'd6741,17'd8982,17'd6741,17'd8342,17'd6734,17'd8823,17'd8984,17'd7222,17'd9136,17'd6100,17'd7057,17'd7217,17'd12331,17'd10921,17'd11734,17'd12783,17'd9815,17'd2422,17'd2422,17'd2935,17'd2934,17'd11888,17'd11888,17'd12784,17'd2119,17'd12785,17'd2430,17'd2430,17'd3105,17'd3105,17'd5658,17'd12655,17'd11889,17'd11890,17'd12786,17'd12787,17'd12788,17'd12789,17'd12790,17'd12791,17'd12792,17'd12793,17'd12794,17'd12795,17'd12513,17'd12796,17'd12797,17'd12798,17'd12799,17'd12800,17'd12801,17'd12051,17'd12802,17'd11904,17'd12803,17'd12671,17'd12804,17'd12805,17'd12806,17'd12807,17'd12808,17'd12809,17'd12675,17'd12213,17'd12810,17'd12811,17'd11761,17'd12677,17'd12812,17'd12813,17'd12065,17'd12814,17'd12530,17'd12815,17'd12362,17'd11913,17'd11764,17'd12681,17'd12681,17'd11362,17'd11629,17'd10691,17'd10691,17'd12533,17'd10817,17'd11232,17'd11232,17'd9158,17'd6142,17'd5409,17'd4927,17'd9302,17'd8066,17'd9007,17'd9007,17'd9301,17'd9301,17'd9159,17'd9159,17'd12219,17'd8368,17'd7414,17'd12816,17'd12817,17'd12818,17'd10280,17'd12819,17'd12820,17'd12538,17'd12368,17'd12069,17'd12821,17'd11918,17'd11484,17'd9849,17'd12822,17'd8387,17'd7265,17'd12823,17'd12824,17'd9319,17'd12825,17'd12826,17'd10132,17'd12827,17'd12828,17'd12829,17'd12546,17'd12830,17'd12831,17'd12832,17'd12227,17'd12833,17'd12834,17'd12693,17'd12694,17'd12835,17'd12836,17'd12837,17'd12838,17'd12839,17'd12840,17'd12841,17'd12842,17'd12564,17'd12843,17'd12701,17'd12844,17'd12845,17'd12846,17'd12847,17'd12706,17'd12707,17'd12708,17'd12848,17'd12848,17'd12849,17'd12242,17'd12850,17'd12710,17'd12712,17'd12572,17'd12099,17'd12851,17'd11656,17'd12852,17'd12853,17'd12854,17'd12717,17'd12855,17'd12856,17'd12419,17'd12110,17'd12857,17'd12858,17'd11958,17'd12414,17'd12418,17'd12859,17'd12860,17'd12415,17'd12253,17'd12579,17'd12109,17'd12110,17'd12113,17'd12861,17'd12862,17'd10605,17'd12863,17'd12116,17'd9344,17'd9188,17'd12864,17'd12865,17'd12725,17'd12866,17'd12867,17'd8251,17'd12726,17'd8258,17'd7791,17'd12868,17'd7629,17'd12869,17'd12870,17'd12871,17'd12872,17'd12873,17'd11287,17'd10872,17'd12126,17'd12874,17'd12275,17'd11152,17'd11413,17'd11413,17'd11413,17'd1045,17'd1045,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd12875,17'd12876,17'd12877,17'd12878,17'd12879,17'd12880,17'd12881,17'd12882,17'd12883,17'd10044,17'd12884,17'd12885,17'd12886,17'd12887,17'd12888,17'd12889,17'd8770,17'd12890,17'd12747,17'd12891,17'd10211,17'd12892,17'd12750,17'd9508,17'd12608,17'd12893,17'd8766,17'd12894,17'd12611,17'd12895,17'd12896,17'd12896,17'd12611,17'd12611,17'd12452,17'd12289,17'd9650,17'd12897,17'd12146,17'd12612,17'd12898,17'd12291,17'd12752,17'd12752,17'd12455,17'd12455,17'd12619,17'd12753,17'd12754,17'd12754,17'd12613,17'd12613,17'd12456,17'd12457,17'd10221,17'd10221,17'd11171,17'd11025,17'd11030,17'd11308,17'd11307,17'd11842,17'd11841,17'd11841,17'd12756,17'd12757,17'd12295,17'd12460,17'd12899,17'd12899,17'd12460,17'd12001,17'd11844,17'd11844,17'd11843,17'd11844,17'd12900,17'd12617,17'd12001,17'd12001,17'd12001,17'd12000,17'd12757,17'd12756,17'd10226,17'd11310,17'd12619,17'd11706,17'd12621,17'd12621,17'd12621,17'd12758,17'd12759,17'd12901,17'd12902,17'd12903,17'd12904,17'd12306,17'd12306,17'd11852,17'd11853,17'd11853,17'd12905,17'd12906,17'd12623,17'd12005,17'd12165,17'd6710,17'd6561,17'd8157,17'd8475,17'd12626,17'd12472,17'd12473,17'd12907,17'd12908,17'd12765,17'd12629,17'd12909,17'd12910,17'd12911,17'd12912,17'd12772,17'd12913,17'd12773,17'd12914,17'd2096,17'd7210,17'd12915,17'd12916,17'd12917,17'd4068,17'd4063,17'd4719,17'd6724,17'd7346,17'd8169,17'd7856,17'd8170,17'd8491,17'd9405,17'd10076,17'd10077,17'd11593,17'd9110,17'd11723,17'd12020,17'd12021,17'd12918,17'd11724,17'd9537,17'd8646,17'd8799,17'd12919,17'd9949,17'd9407,17'd9539,17'd9256,17'd9795,17'd9795,17'd12777,17'd11054,17'd12920,17'd8324,17'd12921,17'd8324,17'd9542,17'd8652,17'd10908,17'd9259,17'd7867,17'd8028,17'd8181,17'd9955,17'd9956,17'd9120,17'd12642,17'd12922,17'd8810,17'd8655,17'd11196,17'd12324,17'd10083,17'd5183,17'd11336,17'd12923,17'd11061,17'd11336,17'd5183,17'd5776,17'd5940,17'd5940,17'd2393,17'd1383,17'd777,17'd1248,17'd2397,17'd12924
},
'{
17'd0,17'd0,17'd0,17'd0,17'd2,17'd2,17'd6419,17'd5196,17'd7545,17'd4887,17'd2422,17'd2422,17'd4247,17'd2,17'd1275,17'd2591,17'd4,17'd6,17'd7,17'd7,17'd5205,17'd5205,17'd8340,17'd8339,17'd8339,17'd8339,17'd8040,17'd5205,17'd7374,17'd11198,17'd12925,17'd12926,17'd7380,17'd7057,17'd9136,17'd5965,17'd8194,17'd7885,17'd8342,17'd8342,17'd10920,17'd9682,17'd7057,17'd8511,17'd6272,17'd9682,17'd7892,17'd5965,17'd12927,17'd8984,17'd6735,17'd11885,17'd6737,17'd12928,17'd12929,17'd1689,17'd10535,17'd2935,17'd11071,17'd12505,17'd471,17'd294,17'd2119,17'd12930,17'd2260,17'd2260,17'd2264,17'd4739,17'd5379,17'd12931,17'd6110,17'd11737,17'd11890,17'd5807,17'd5218,17'd12339,17'd12790,17'd12932,17'd12933,17'd12934,17'd12935,17'd12936,17'd12937,17'd12938,17'd12939,17'd12940,17'd12941,17'd12942,17'd11468,17'd12518,17'd12943,17'd12944,17'd12803,17'd11905,17'd12945,17'd12946,17'd12947,17'd12948,17'd12949,17'd12950,17'd12951,17'd12058,17'd12952,17'd12953,17'd12526,17'd11084,17'd12677,17'd12954,17'd12955,17'd12218,17'd12218,17'd12956,17'd12957,17'd12680,17'd11764,17'd11628,17'd12681,17'd12681,17'd11629,17'd11629,17'd10562,17'd10691,17'd10112,17'd10112,17'd12535,17'd8687,17'd12220,17'd8369,17'd10430,17'd7582,17'd8538,17'd9007,17'd12958,17'd12959,17'd10113,17'd9703,17'd8537,17'd9159,17'd9158,17'd7086,17'd9296,17'd12960,17'd12961,17'd12683,17'd10812,17'd12962,17'd12820,17'd12368,17'd12069,17'd12821,17'd11919,17'd11919,17'd10569,17'd9707,17'd9016,17'd8548,17'd8855,17'd10702,17'd9319,17'd12072,17'd12222,17'd11485,17'd9854,17'd12963,17'd12964,17'd12965,17'd12966,17'd12967,17'd12968,17'd12969,17'd12970,17'd12971,17'd12972,17'd12973,17'd12974,17'd12975,17'd12976,17'd12977,17'd12978,17'd12979,17'd12980,17'd12981,17'd12240,17'd12238,17'd12982,17'd12983,17'd12984,17'd12985,17'd12558,17'd12986,17'd12707,17'd12987,17'd12988,17'd12567,17'd12567,17'd12400,17'd12849,17'd12243,17'd12989,17'd12402,17'd11789,17'd12990,17'd12713,17'd12991,17'd12992,17'd12993,17'd12994,17'd12257,17'd12256,17'd12995,17'd12419,17'd12419,17'd11961,17'd12996,17'd11958,17'd12109,17'd12859,17'd12997,17'd12860,17'd12415,17'd12418,17'd12856,17'd12419,17'd12110,17'd12998,17'd12999,17'd13000,17'd13001,17'd12863,17'd9741,17'd9346,17'd8875,17'd13002,17'd12865,17'd13003,17'd13004,17'd13005,17'd8252,17'd13006,17'd13007,17'd7791,17'd8428,17'd7629,17'd13008,17'd13009,17'd13010,17'd13011,17'd13012,17'd11287,17'd13013,17'd12273,17'd10621,17'd7812,17'd8131,17'd11289,17'd11413,17'd11413,17'd1045,17'd1045,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd133,17'd132,17'd132,17'd3169,17'd9361,17'd13014,17'd13015,17'd13016,17'd13017,17'd13018,17'd13019,17'd13020,17'd13021,17'd13022,17'd9069,17'd13023,17'd13024,17'd13025,17'd13025,17'd12746,17'd8923,17'd10054,17'd12748,17'd13026,17'd13027,17'd9224,17'd13028,17'd12608,17'd12893,17'd8766,17'd12611,17'd12611,17'd12896,17'd8456,17'd8456,17'd8456,17'd8294,17'd8153,17'd7996,17'd8464,17'd12290,17'd12751,17'd12898,17'd13029,17'd12752,17'd12752,17'd12752,17'd12619,17'd12619,17'd12619,17'd12619,17'd12754,17'd13030,17'd13031,17'd13032,17'd11306,17'd11305,17'd11310,17'd10221,17'd10222,17'd10223,17'd13033,17'd13034,17'd11308,17'd11307,17'd11842,17'd11841,17'd12756,17'd12756,17'd12295,17'd12295,17'd13035,17'd12899,17'd13036,17'd12756,17'd11843,17'd11843,17'd11843,17'd11844,17'd11844,17'd11843,17'd12001,17'd11843,17'd11844,17'd11844,17'd12296,17'd12757,17'd12296,17'd10226,17'd11847,17'd13037,17'd13038,17'd13039,17'd13038,17'd13040,17'd13041,17'd13042,17'd13043,17'd13044,17'd12904,17'd11852,17'd13045,17'd12306,17'd11575,17'd11429,17'd11577,17'd13046,17'd12623,17'd12762,17'd13047,17'd8155,17'd8473,17'd8156,17'd7331,17'd7841,17'd12626,17'd12310,17'd13048,17'd13049,17'd13050,17'd13051,17'd13052,17'd13053,17'd13054,17'd12633,17'd13055,17'd13056,17'd12773,17'd6582,17'd1810,17'd7210,17'd8165,17'd13057,17'd13058,17'd2753,17'd6249,17'd5033,17'd6576,17'd7346,17'd8169,17'd7856,17'd8171,17'd8019,17'd9405,17'd10076,17'd10077,17'd11593,17'd9110,17'd11723,17'd13059,17'd12020,17'd11873,17'd11873,17'd10527,17'd8957,17'd9538,17'd9949,17'd9256,17'd9538,17'd9539,17'd9538,17'd9795,17'd9795,17'd9795,17'd11725,17'd8962,17'd7690,17'd12921,17'd9411,17'd8652,17'd8652,17'd10908,17'd8027,17'd10653,17'd9955,17'd8181,17'd9955,17'd9120,17'd9120,17'd12322,17'd12490,17'd8810,17'd8810,17'd11196,17'd12324,17'd13060,17'd9670,17'd5183,17'd12495,17'd11061,17'd11336,17'd5183,17'd5776,17'd5940,17'd12496,17'd414,17'd415,17'd418,17'd2102,17'd13061,17'd12498
},
'{
17'd0,17'd0,17'd0,17'd0,17'd2,17'd1127,17'd5196,17'd6583,17'd4887,17'd4887,17'd2422,17'd1688,17'd466,17'd3,17'd2933,17'd2421,17'd5,17'd6,17'd7,17'd7,17'd5205,17'd8040,17'd8339,17'd8339,17'd8339,17'd8339,17'd8040,17'd5205,17'd7216,17'd13062,17'd13063,17'd6901,17'd7892,17'd8815,17'd5965,17'd5964,17'd6104,17'd6429,17'd7714,17'd6742,17'd7222,17'd6900,17'd8670,17'd8815,17'd9137,17'd7057,17'd9136,17'd6100,17'd11201,17'd10403,17'd13064,17'd6737,17'd6735,17'd13065,17'd1689,17'd2594,17'd10535,17'd2935,17'd12196,17'd12653,17'd294,17'd34,17'd2119,17'd2119,17'd2260,17'd13066,17'd2604,17'd5055,17'd13067,17'd6110,17'd11737,17'd11737,17'd13068,17'd13069,17'd13070,17'd13071,17'd13072,17'd13073,17'd13074,17'd13075,17'd13076,17'd13077,17'd13078,17'd13079,17'd13080,17'd13081,17'd13082,17'd13083,17'd11902,17'd12943,17'd12944,17'd12803,17'd13084,17'd13085,17'd12946,17'd13086,17'd13087,17'd13088,17'd13089,17'd13090,17'd13091,17'd12058,17'd12952,17'd12676,17'd11084,17'd12062,17'd13092,17'd13093,17'd13094,17'd13094,17'd11360,17'd11360,17'd12680,17'd11913,17'd11764,17'd11628,17'd12681,17'd12532,17'd10815,17'd10815,17'd10562,17'd10427,17'd10112,17'd10112,17'd8687,17'd8368,17'd12220,17'd12219,17'd9007,17'd8538,17'd8538,17'd9301,17'd13095,17'd13095,17'd10113,17'd9703,17'd9159,17'd9006,17'd8687,17'd7414,17'd13096,17'd13097,17'd13098,17'd13099,17'd13100,17'd12962,17'd13101,17'd13102,17'd12821,17'd13103,17'd11630,17'd9848,17'd13104,17'd13105,17'd13106,17'd8702,17'd9169,17'd9319,17'd12072,17'd12222,17'd11485,17'd9854,17'd13107,17'd13108,17'd13109,17'd13110,17'd12966,17'd13111,17'd13112,17'd13113,17'd13114,17'd12971,17'd13115,17'd12973,17'd12975,17'd12976,17'd13116,17'd13117,17'd13118,17'd13119,17'd13120,17'd13121,17'd12091,17'd13122,17'd13123,17'd13124,17'd13125,17'd13126,17'd13127,17'd13128,17'd12566,17'd12707,17'd13129,17'd12567,17'd12706,17'd13130,17'd12849,17'd13131,17'd12094,17'd12571,17'd12990,17'd12713,17'd12714,17'd13132,17'd13133,17'd13134,17'd12256,17'd12856,17'd12856,17'd12995,17'd12419,17'd12419,17'd11961,17'd13135,17'd11958,17'd12110,17'd12578,17'd12859,17'd12860,17'd12415,17'd12418,17'd12417,17'd12109,17'd12419,17'd13136,17'd12857,17'd13137,17'd13138,17'd11400,17'd10024,17'd9340,17'd8873,17'd10607,17'd8578,17'd12867,17'd13139,17'd13139,17'd8252,17'd13140,17'd13141,17'd7956,17'd8428,17'd13142,17'd13008,17'd13143,17'd13010,17'd11146,17'd11411,17'd13144,17'd13145,17'd12273,17'd10621,17'd7812,17'd10873,17'd11152,17'd11413,17'd11413,17'd11413,17'd1045,17'd1045,17'd133,17'd133,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd134,17'd131,17'd3512,17'd5470,17'd13146,17'd13147,17'd4009,17'd13148,17'd13149,17'd13150,17'd13151,17'd13152,17'd10500,17'd13153,17'd13154,17'd13024,17'd13155,17'd13156,17'd8459,17'd12890,17'd12747,17'd12747,17'd13157,17'd13158,17'd12608,17'd12608,17'd12893,17'd8765,17'd12611,17'd12611,17'd12611,17'd12896,17'd8456,17'd8456,17'd8456,17'd13159,17'd7997,17'd7996,17'd8465,17'd13160,17'd12898,17'd12291,17'd12752,17'd12752,17'd12752,17'd12752,17'd12619,17'd12619,17'd12753,17'd12753,17'd12754,17'd13031,17'd13161,17'd13161,17'd11170,17'd11306,17'd13037,17'd12755,17'd10223,17'd10224,17'd13034,17'd13034,17'd11174,17'd11173,17'd11307,17'd12458,17'd12296,17'd12756,17'd12154,17'd12154,17'd13162,17'd12295,17'd12757,17'd13163,17'd12460,17'd12001,17'd11844,17'd11844,17'd11843,17'd11843,17'd11843,17'd11843,17'd11843,17'd11843,17'd12296,17'd12757,17'd12756,17'd12297,17'd10224,17'd11310,17'd13040,17'd13038,17'd13038,17'd13040,17'd12902,17'd13041,17'd13164,17'd13042,17'd11852,17'd11852,17'd13045,17'd13165,17'd13166,17'd11575,17'd11709,17'd12905,17'd11855,17'd13167,17'd13168,17'd13169,17'd8630,17'd6394,17'd8157,17'd7331,17'd8475,17'd7332,17'd12472,17'd13170,17'd13049,17'd12765,17'd13171,17'd13172,17'd13173,17'd13174,17'd13175,17'd13056,17'd13176,17'd13177,17'd4575,17'd2905,17'd2576,17'd13178,17'd1391,17'd13179,17'd2247,17'd4563,17'd7193,17'd6724,17'd8169,17'd7856,17'd7856,17'd8171,17'd8019,17'd9405,17'd10077,17'd10077,17'd10650,17'd11723,17'd13059,17'd13059,17'd12021,17'd11873,17'd11594,17'd9537,17'd9538,17'd9949,17'd9256,17'd9949,17'd9538,17'd9539,17'd9795,17'd9795,17'd9795,17'd12777,17'd9666,17'd8650,17'd8324,17'd8324,17'd9542,17'd8652,17'd10908,17'd10908,17'd11195,17'd9799,17'd8181,17'd9955,17'd9956,17'd9956,17'd9956,17'd9120,17'd8810,17'd8655,17'd11196,17'd10910,17'd13180,17'd9804,17'd3570,17'd2906,17'd11336,17'd11336,17'd5183,17'd9123,17'd5630,17'd8185,17'd12496,17'd413,17'd1672,17'd599,17'd2102,17'd13061
},
'{
17'd2,17'd2,17'd14,17'd14,17'd14,17'd1689,17'd4886,17'd7545,17'd2935,17'd2784,17'd3250,17'd1127,17'd12,17'd1275,17'd4242,17'd7215,17'd6,17'd7,17'd8190,17'd8190,17'd8340,17'd8340,17'd8339,17'd8339,17'd8339,17'd8339,17'd8340,17'd10537,17'd11198,17'd10916,17'd13181,17'd6901,17'd6900,17'd8042,17'd5964,17'd6589,17'd9415,17'd7376,17'd6429,17'd10920,17'd7892,17'd8825,17'd13182,17'd13183,17'd7058,17'd9136,17'd8987,17'd6434,17'd9132,17'd13184,17'd6735,17'd6736,17'd13185,17'd13186,17'd4247,17'd2594,17'd10547,17'd11071,17'd12505,17'd12504,17'd35,17'd2120,17'd2260,17'd2939,17'd12785,17'd2264,17'd4739,17'd13067,17'd12337,17'd12337,17'd12337,17'd5807,17'd13187,17'd13188,17'd13189,17'd3438,17'd13190,17'd13191,17'd13192,17'd13193,17'd13194,17'd13195,17'd12939,17'd13196,17'd13197,17'd13198,17'd13199,17'd13200,17'd11752,17'd12943,17'd13201,17'd12804,17'd12945,17'd13202,17'd13203,17'd13204,17'd13205,17'd13089,17'd13090,17'd13206,17'd12058,17'd12058,17'd13207,17'd13208,17'd11084,17'd12357,17'd13209,17'd13210,17'd13211,17'd13094,17'd11360,17'd12956,17'd12066,17'd11361,17'd11230,17'd11230,17'd11764,17'd11913,17'd11914,17'd11914,17'd10691,17'd10427,17'd10286,17'd10286,17'd8536,17'd8368,17'd12219,17'd13212,17'd9007,17'd9704,17'd9575,17'd12959,17'd13095,17'd12959,17'd10113,17'd9703,17'd9574,17'd9573,17'd13213,17'd13214,17'd13215,17'd13216,17'd13217,17'd13218,17'd13219,17'd13220,17'd13101,17'd12368,17'd13221,17'd13103,17'd11094,17'd9310,17'd9016,17'd8853,17'd8702,17'd13222,17'd9171,17'd10703,17'd12222,17'd13223,17'd10820,17'd13224,17'd13108,17'd13109,17'd13110,17'd13225,17'd13226,17'd13227,17'd13228,17'd13229,17'd13230,17'd12971,17'd12972,17'd12973,17'd13231,17'd13232,17'd13233,17'd13234,17'd13235,17'd13236,17'd13237,17'd13238,17'd13239,17'd13240,17'd13124,17'd13241,17'd13242,17'd13243,17'd13244,17'd13245,17'd13246,17'd13246,17'd12567,17'd12400,17'd12706,17'd13130,17'd13247,17'd13131,17'd12094,17'd13248,17'd13249,17'd12991,17'd13250,17'd13251,17'd13134,17'd12860,17'd12859,17'd12417,17'd12580,17'd12580,17'd12420,17'd12113,17'd11962,17'd12861,17'd11961,17'd12110,17'd12578,17'd12578,17'd12859,17'd12859,17'd12859,17'd12418,17'd12109,17'd12109,17'd13252,17'd13136,17'd13253,17'd13254,17'd12423,17'd10167,17'd13255,17'd9189,17'd8730,17'd13256,17'd13257,17'd12426,17'd12588,17'd13258,17'd7786,17'd8257,17'd7956,17'd13259,17'd7629,17'd12730,17'd13009,17'd13010,17'd11146,17'd11411,17'd10488,17'd13260,17'd9631,17'd9495,17'd7812,17'd8131,17'd8132,17'd8132,17'd8132,17'd8132,17'd1045,17'd1045,17'd1197,17'd1197,17'd134,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd357,17'd3812,17'd13261,17'd13262,17'd13263,17'd4010,17'd13264,17'd13265,17'd13266,17'd13267,17'd13268,17'd8453,17'd13269,17'd13270,17'd13271,17'd13272,17'd13272,17'd12890,17'd13273,17'd12891,17'd12748,17'd13274,17'd13158,17'd13275,17'd8919,17'd12893,17'd8766,17'd12611,17'd12450,17'd8294,17'd8294,17'd12283,17'd12283,17'd8293,17'd8293,17'd7994,17'd7997,17'd8627,17'd8778,17'd9520,17'd12752,17'd12752,17'd12752,17'd11706,17'd11706,17'd11706,17'd12002,17'd11706,17'd11706,17'd12753,17'd13037,17'd13031,17'd13031,17'd11170,17'd11170,17'd13037,17'd10229,17'd11310,17'd10221,17'd10223,17'd10224,17'd10224,17'd10224,17'd10225,17'd11309,17'd12297,17'd12296,17'd12000,17'd12000,17'd12154,17'd12154,17'd12756,17'd13163,17'd13163,17'd12757,17'd12001,17'd11843,17'd11843,17'd11844,17'd11844,17'd11843,17'd12001,17'd11843,17'd11843,17'd12001,17'd12154,17'd12757,17'd12155,17'd10377,17'd13276,17'd13040,17'd13040,17'd13040,17'd13040,17'd13040,17'd13277,17'd13277,17'd13042,17'd13044,17'd13045,17'd13165,17'd13278,17'd13166,17'd11709,17'd11577,17'd11711,17'd13279,17'd13280,17'd13047,17'd13281,17'd7670,17'd8156,17'd8157,17'd11433,17'd13282,17'd13283,17'd13284,17'd13285,17'd12908,17'd13286,17'd13287,17'd13288,17'd13289,17'd12912,17'd12772,17'd12913,17'd13177,17'd4575,17'd6415,17'd412,17'd2762,17'd13290,17'd13058,17'd2401,17'd13291,17'd7031,17'd6576,17'd7346,17'd8169,17'd7856,17'd7856,17'd8019,17'd9405,17'd10391,17'd10391,17'd12487,17'd12488,17'd12489,17'd12489,17'd12021,17'd11873,17'd13292,17'd13293,17'd11595,17'd9112,17'd9112,17'd9112,17'd9949,17'd9538,17'd9795,17'd9795,17'd11192,17'd12777,17'd11054,17'd9541,17'd8650,17'd7690,17'd9542,17'd9542,17'd9411,17'd9411,17'd12641,17'd10653,17'd9955,17'd8181,17'd8181,17'd9955,17'd10256,17'd9120,17'd12492,17'd12492,17'd8655,17'd12493,17'd13294,17'd9803,17'd11334,17'd8187,17'd11336,17'd11061,17'd5183,17'd9123,17'd5630,17'd8185,17'd6868,17'd951,17'd778,17'd418,17'd1813,17'd1673
},
'{
17'd466,17'd466,17'd14,17'd14,17'd1689,17'd1688,17'd7545,17'd5508,17'd2935,17'd2422,17'd1688,17'd14,17'd3,17'd2591,17'd2421,17'd7373,17'd7,17'd7,17'd8190,17'd8190,17'd8340,17'd8340,17'd8339,17'd13295,17'd13295,17'd8340,17'd8190,17'd7727,17'd13296,17'd13063,17'd13297,17'd13298,17'd13183,17'd5962,17'd5964,17'd8511,17'd7885,17'd7885,17'd6271,17'd9271,17'd8973,17'd13182,17'd6427,17'd13299,17'd13300,17'd6435,17'd13301,17'd8511,17'd6734,17'd6740,17'd6431,17'd9550,17'd13302,17'd6583,17'd1831,17'd1689,17'd10547,17'd10924,17'd12505,17'd12504,17'd35,17'd2120,17'd2260,17'd13303,17'd2430,17'd3105,17'd5210,17'd12507,17'd12337,17'd5661,17'd5807,17'd13069,17'd13304,17'd13305,17'd13306,17'd13307,17'd13308,17'd13309,17'd13310,17'd13311,17'd13312,17'd12939,17'd13313,17'd13314,17'd13198,17'd13315,17'd13316,17'd13317,17'd11904,17'd11904,17'd13318,17'd13085,17'd13319,17'd13320,17'd13321,17'd12949,17'd13322,17'd13323,17'd13324,17'd13206,17'd13325,17'd13326,17'd12354,17'd12526,17'd12062,17'd13092,17'd13210,17'd12955,17'd13094,17'd13094,17'd12956,17'd11627,17'd12066,17'd11361,17'd11230,17'd11230,17'd11764,17'd11913,17'd11914,17'd11914,17'd10427,17'd10427,17'd13327,17'd8687,17'd12220,17'd6468,17'd13212,17'd12534,17'd13328,17'd9575,17'd12959,17'd13095,17'd12959,17'd12959,17'd10113,17'd10113,17'd9702,17'd7250,17'd13329,17'd13330,17'd13331,17'd13332,17'd13333,17'd13334,17'd13335,17'd13336,17'd13337,17'd12368,17'd13221,17'd11093,17'd9310,17'd9018,17'd8701,17'd8702,17'd8857,17'd10702,17'd11240,17'd11921,17'd11769,17'd9713,17'd13224,17'd13338,17'd13339,17'd13109,17'd13110,17'd12966,17'd13340,17'd13341,17'd13342,17'd13343,17'd13344,17'd13345,17'd12972,17'd12835,17'd13346,17'd13347,17'd11781,17'd11931,17'd13348,17'd12981,17'd13349,17'd13350,17'd13351,17'd11251,17'd12984,17'd13352,17'd13353,17'd13354,17'd12566,17'd12708,17'd13246,17'd13355,17'd13356,17'd12400,17'd13130,17'd13357,17'd13358,17'd13359,17'd12572,17'd11800,17'd13360,17'd13132,17'd13133,17'd13361,17'd12997,17'd12415,17'd12416,17'd12416,17'd12106,17'd12420,17'd12113,17'd12996,17'd13362,17'd11962,17'd13363,17'd13364,17'd12577,17'd12414,17'd12418,17'd12418,17'd12859,17'd12859,17'd12414,17'd12109,17'd12995,17'd13365,17'd13366,17'd13367,17'd13368,17'd13369,17'd13370,17'd10175,17'd13371,17'd13372,17'd13373,17'd13374,17'd13373,17'd13375,17'd13376,17'd13377,17'd13378,17'd13259,17'd10612,17'd13379,17'd13009,17'd13010,17'd11146,17'd13380,17'd13381,17'd13382,17'd9631,17'd9495,17'd7812,17'd10873,17'd10874,17'd8132,17'd8132,17'd8132,17'd11413,17'd1045,17'd1197,17'd1197,17'd134,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd357,17'd3812,17'd13383,17'd13384,17'd13385,17'd13386,17'd13387,17'd13388,17'd13389,17'd13390,17'd13391,17'd13392,17'd13393,17'd13394,17'd13395,17'd13396,17'd13396,17'd13397,17'd13398,17'd10505,17'd12891,17'd13157,17'd13399,17'd12893,17'd11834,17'd8766,17'd12894,17'd12450,17'd12145,17'd13400,17'd13400,17'd12283,17'd12283,17'd8293,17'd7832,17'd7831,17'd13401,17'd13402,17'd13402,17'd12752,17'd12752,17'd12752,17'd12752,17'd11706,17'd11706,17'd12002,17'd12002,17'd12002,17'd12002,17'd11706,17'd12619,17'd12619,17'd13403,17'd11305,17'd12457,17'd10228,17'd10229,17'd13404,17'd11847,17'd11310,17'd10223,17'd10224,17'd10224,17'd10224,17'd10225,17'd11705,17'd12297,17'd12000,17'd12000,17'd12000,17'd12154,17'd12757,17'd12756,17'd12757,17'd13163,17'd12899,17'd12000,17'd11844,17'd11845,17'd11844,17'd11843,17'd12001,17'd11843,17'd11845,17'd11844,17'd12000,17'd12460,17'd12757,17'd11309,17'd13405,17'd13276,17'd13276,17'd13276,17'd13040,17'd13040,17'd13043,17'd13164,17'd13164,17'd13041,17'd12306,17'd13165,17'd13406,17'd13407,17'd11431,17'd11431,17'd11579,17'd12623,17'd13168,17'd13408,17'd12164,17'd6559,17'd6394,17'd8156,17'd8634,17'd13409,17'd13410,17'd13411,17'd13412,17'd13413,17'd13414,17'd13415,17'd13416,17'd13417,17'd13418,17'd13419,17'd13056,17'd13420,17'd6259,17'd5372,17'd2409,17'd780,17'd949,17'd13421,17'd1953,17'd13422,17'd5946,17'd6243,17'd6724,17'd7685,17'd8169,17'd7856,17'd8019,17'd9405,17'd9946,17'd10391,17'd10077,17'd12320,17'd13423,17'd13424,17'd13425,17'd12021,17'd13292,17'd13426,17'd11724,17'd9112,17'd9112,17'd9112,17'd9949,17'd9949,17'd9795,17'd9795,17'd11192,17'd9795,17'd11725,17'd9666,17'd8962,17'd8650,17'd9411,17'd9542,17'd9542,17'd7691,17'd11193,17'd10653,17'd9955,17'd8181,17'd8181,17'd9955,17'd9956,17'd12322,17'd12642,17'd12492,17'd8655,17'd8655,17'd11196,17'd13427,17'd12494,17'd6727,17'd5183,17'd11061,17'd5183,17'd4714,17'd5630,17'd8185,17'd6868,17'd2575,17'd779,17'd778,17'd417,17'd1813
},
'{
17'd14,17'd14,17'd14,17'd14,17'd1689,17'd2422,17'd5508,17'd13428,17'd3250,17'd3250,17'd1127,17'd0,17'd1275,17'd4242,17'd6,17'd3753,17'd5205,17'd5205,17'd8190,17'd8190,17'd8340,17'd8340,17'd8339,17'd8339,17'd13295,17'd13429,17'd8340,17'd12648,17'd13062,17'd13430,17'd13431,17'd8825,17'd6099,17'd5798,17'd5965,17'd9272,17'd6733,17'd9551,17'd11204,17'd8815,17'd6435,17'd8661,17'd8347,17'd13432,17'd7724,17'd11730,17'd8815,17'd9415,17'd13433,17'd6740,17'd10401,17'd13434,17'd13435,17'd13436,17'd1831,17'd2422,17'd10670,17'd10925,17'd471,17'd471,17'd1968,17'd1968,17'd2939,17'd3103,17'd3253,17'd3435,17'd12336,17'd12786,17'd5384,17'd5383,17'd13437,17'd13438,17'd13439,17'd2437,17'd13440,17'd13441,17'd13442,17'd13443,17'd13311,17'd13444,17'd13445,17'd13446,17'd13447,17'd13448,17'd13449,17'd13450,17'd13451,17'd13452,17'd13453,17'd11905,17'd13084,17'd13454,17'd13455,17'd13456,17'd13457,17'd12950,17'd13090,17'd13458,17'd13206,17'd13459,17'd13459,17'd12212,17'd13460,17'd13461,17'd13462,17'd13463,17'd13210,17'd13210,17'd12955,17'd12065,17'd13464,17'd11627,17'd11361,17'd11230,17'd11230,17'd11230,17'd11361,17'd12066,17'd10815,17'd10815,17'd10563,17'd10427,17'd12533,17'd9158,17'd12219,17'd8370,17'd13212,17'd13465,17'd9575,17'd13466,17'd13467,17'd13468,17'd13469,17'd13470,17'd10565,17'd13471,17'd13472,17'd13473,17'd13474,17'd13475,17'd13476,17'd13477,17'd13478,17'd13479,17'd13337,17'd13480,17'd13481,17'd13482,17'd11918,17'd13483,17'd9445,17'd13484,17'd8702,17'd8224,17'd9021,17'd13485,17'd11632,17'd11366,17'd9713,17'd12827,17'd13486,17'd13487,17'd13488,17'd13488,17'd12965,17'd13226,17'd13489,17'd13490,17'd13229,17'd13491,17'd13344,17'd12079,17'd12834,17'd11778,17'd13492,17'd12978,17'd13493,17'd13494,17'd12847,17'd12240,17'd13495,17'd13496,17'd13123,17'd13124,17'd12846,17'd13497,17'd13498,17'd13499,17'd13500,17'd13501,17'd13502,17'd13502,17'd13502,17'd13503,17'd13504,17'd13505,17'd13506,17'd13507,17'd13508,17'd13509,17'd13510,17'd13511,17'd13512,17'd12417,17'd13513,17'd13514,17'd13515,17'd12416,17'd12580,17'd12581,17'd12996,17'd11806,17'd13362,17'd13516,17'd11963,17'd13363,17'd12577,17'd12109,17'd13517,17'd12417,17'd12997,17'd12859,17'd12109,17'd12856,17'd13518,17'd13519,17'd13520,17'd11522,17'd13521,17'd13522,17'd9620,17'd9194,17'd13523,17'd13524,17'd13525,17'd13526,17'd13527,17'd12427,17'd13376,17'd7620,17'd13528,17'd13529,17'd8739,17'd8740,17'd13530,17'd13531,17'd11285,17'd13532,17'd13381,17'd13382,17'd10036,17'd13533,17'd11977,17'd12275,17'd11152,17'd10874,17'd8132,17'd8132,17'd11413,17'd11413,17'd3025,17'd1197,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd132,17'd133,17'd133,17'd134,17'd131,17'd13534,17'd13535,17'd7816,17'd13536,17'd13537,17'd13538,17'd13539,17'd13540,17'd13541,17'd13542,17'd13543,17'd13544,17'd13545,17'd13395,17'd13396,17'd13546,17'd13397,17'd13547,17'd10505,17'd13548,17'd13274,17'd13399,17'd12141,17'd12141,17'd8765,17'd12449,17'd12145,17'd12451,17'd8294,17'd13400,17'd12282,17'd12283,17'd8293,17'd11296,17'd7828,17'd7830,17'd8627,17'd8778,17'd13549,17'd12454,17'd12752,17'd13550,17'd13551,17'd11567,17'd10511,17'd10775,17'd10511,17'd10511,17'd10775,17'd11567,17'd12454,17'd12752,17'd13552,17'd13552,17'd9654,17'd9654,17'd9654,17'd10061,17'd11847,17'd12755,17'd11310,17'd10221,17'd9780,17'd9780,17'd9780,17'd9384,17'd11705,17'd12297,17'd12000,17'd12154,17'd12296,17'd12155,17'd12155,17'd12757,17'd12899,17'd12295,17'd11843,17'd11844,17'd11844,17'd11843,17'd12001,17'd11843,17'd11844,17'd11844,17'd11843,17'd12000,17'd12756,17'd12296,17'd10510,17'd13161,17'd13553,17'd13554,17'd13405,17'd13555,17'd13041,17'd13043,17'd13277,17'd13043,17'd13556,17'd13556,17'd13557,17'd13558,17'd12760,17'd11853,17'd12160,17'd12161,17'd13559,17'd13280,17'd13560,17'd13561,17'd13562,17'd7502,17'd7330,17'd13563,17'd13410,17'd13411,17'd13284,17'd13564,17'd13565,17'd13566,17'd13567,17'd13568,17'd13569,17'd13570,17'd13571,17'd13572,17'd13177,17'd4728,17'd412,17'd951,17'd13573,17'd1108,17'd1953,17'd2401,17'd4064,17'd5946,17'd6576,17'd7685,17'd7858,17'd8020,17'd8171,17'd8019,17'd10076,17'd11722,17'd10391,17'd12487,17'd11723,17'd12489,17'd13425,17'd13425,17'd12021,17'd12021,17'd11873,17'd11595,17'd9112,17'd11595,17'd9256,17'd9949,17'd12777,17'd9795,17'd9795,17'd9795,17'd11725,17'd11054,17'd9541,17'd8962,17'd9411,17'd9411,17'd9542,17'd9542,17'd11193,17'd11193,17'd10653,17'd8181,17'd8181,17'd8181,17'd9956,17'd9956,17'd12322,17'd12491,17'd12492,17'd10654,17'd11196,17'd12324,17'd9803,17'd6727,17'd5183,17'd12495,17'd9123,17'd9123,17'd5630,17'd5630,17'd11062,17'd951,17'd601,17'd1246,17'd416,17'd416
},
'{
17'd14,17'd1127,17'd1127,17'd1689,17'd3250,17'd2422,17'd5508,17'd5508,17'd3250,17'd1689,17'd2,17'd12,17'd2933,17'd2421,17'd6,17'd5205,17'd5205,17'd5205,17'd8190,17'd8190,17'd8340,17'd8340,17'd8339,17'd8339,17'd13295,17'd8040,17'd10537,17'd10796,17'd13574,17'd13430,17'd6427,17'd8661,17'd5797,17'd11730,17'd6106,17'd8194,17'd6104,17'd9966,17'd8824,17'd6732,17'd6732,17'd8661,17'd6427,17'd13575,17'd8347,17'd6428,17'd9137,17'd6269,17'd13576,17'd6735,17'd9545,17'd13577,17'd12647,17'd13436,17'd2784,17'd2782,17'd11071,17'd11888,17'd471,17'd294,17'd1968,17'd2428,17'd13578,17'd3103,17'd3431,17'd3756,17'd12655,17'd5974,17'd13579,17'd5058,17'd4255,17'd13439,17'd13580,17'd835,17'd13581,17'd13582,17'd3767,17'd13583,17'd13584,17'd13585,17'd13586,17'd13587,17'd13588,17'd13589,17'd13590,17'd13591,17'd13451,17'd13451,17'd12945,17'd13085,17'd13592,17'd13593,17'd12947,17'd12056,17'd13594,17'd12809,17'd13091,17'd13091,17'd13206,17'd13595,17'd13595,17'd13596,17'd13461,17'd13597,17'd13598,17'd13463,17'd13599,17'd12955,17'd12065,17'd12814,17'd11763,17'd11627,17'd11361,17'd11361,17'd11361,17'd12066,17'd12066,17'd12066,17'd11629,17'd10427,17'd10427,17'd12533,17'd9573,17'd12219,17'd13212,17'd10430,17'd13600,17'd8067,17'd13095,17'd13466,17'd13468,17'd13468,17'd13601,17'd13601,17'd10429,17'd13602,17'd13603,17'd13604,17'd13605,17'd13606,17'd13477,17'd13607,17'd13334,17'd13608,17'd13609,17'd13610,17'd12368,17'd11483,17'd10289,17'd9849,17'd13611,17'd13612,17'd8224,17'd13613,17'd13614,17'd11632,17'd12072,17'd10819,17'd13615,17'd12963,17'd13487,17'd13616,17'd13617,17'd13618,17'd12830,17'd13619,17'd13620,17'd13113,17'd13621,17'd13230,17'd13622,17'd11639,17'd11640,17'd13623,17'd13624,17'd13625,17'd13626,17'd11785,17'd13627,17'd13238,17'd13628,17'd13629,17'd13630,17'd13631,17'd13632,17'd13354,17'd13633,17'd13499,17'd13634,17'd13635,17'd13636,17'd13636,17'd13636,17'd12236,17'd13637,17'd13638,17'd12405,17'd11944,17'd13639,17'd13640,17'd13641,17'd13642,17'd13643,17'd12418,17'd13644,17'd13514,17'd12417,17'd12418,17'd12109,17'd11958,17'd13135,17'd12996,17'd13516,17'd13645,17'd13362,17'd13135,17'd12110,17'd12109,17'd13517,17'd12417,17'd12997,17'd12859,17'd12109,17'd12856,17'd12856,17'd13136,17'd13646,17'd13254,17'd13647,17'd10169,17'd10174,17'd8728,17'd13648,17'd13649,17'd13650,17'd13651,17'd13652,17'd13649,17'd13653,17'd13654,17'd13528,17'd13529,17'd8739,17'd8740,17'd13530,17'd13655,17'd13656,17'd13532,17'd13381,17'd13657,17'd10036,17'd13533,17'd11977,17'd12275,17'd11152,17'd10874,17'd8132,17'd8132,17'd11413,17'd11413,17'd3025,17'd1197,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd132,17'd133,17'd133,17'd132,17'd131,17'd2865,17'd11822,17'd13658,17'd13659,17'd13660,17'd13265,17'd13661,17'd13267,17'd13662,17'd13663,17'd13664,17'd13665,17'd13666,17'd13667,17'd13546,17'd13668,17'd13273,17'd13669,17'd10505,17'd13670,17'd10211,17'd13671,17'd12141,17'd12141,17'd12894,17'd11994,17'd12452,17'd12451,17'd8294,17'd8294,17'd12282,17'd12282,17'd13672,17'd11296,17'd7832,17'd13673,17'd8627,17'd13402,17'd9783,17'd13550,17'd12454,17'd13549,17'd13674,17'd10775,17'd10511,17'd10230,17'd10775,17'd10511,17'd10230,17'd9656,17'd9656,17'd9783,17'd9783,17'd9656,17'd9236,17'd13675,17'd13675,17'd9655,17'd13404,17'd11847,17'd12755,17'd11310,17'd10063,17'd9517,17'd9780,17'd9384,17'd10226,17'd11705,17'd12297,17'd12296,17'd12155,17'd12297,17'd12296,17'd12297,17'd12000,17'd12295,17'd12154,17'd12001,17'd11844,17'd11843,17'd11843,17'd11843,17'd11844,17'd11844,17'd11843,17'd12001,17'd12757,17'd12757,17'd12297,17'd10224,17'd13554,17'd13676,17'd13555,17'd13405,17'd13043,17'd13042,17'd13043,17'd13277,17'd13677,17'd13556,17'd13556,17'd13677,17'd13278,17'd11854,17'd13678,17'd13679,17'd12163,17'd13559,17'd12308,17'd13047,17'd6709,17'd7670,17'd8157,17'd7331,17'd7505,17'd13680,17'd13681,17'd13564,17'd13682,17'd13683,17'd13684,17'd13685,17'd13686,17'd13687,17'd13688,17'd13689,17'd13176,17'd4728,17'd412,17'd602,17'd194,17'd1109,17'd7192,17'd1818,17'd4408,17'd4720,17'd7193,17'd7346,17'd7686,17'd7858,17'd8171,17'd8019,17'd9405,17'd10076,17'd13690,17'd10077,17'd11872,17'd13423,17'd13059,17'd13691,17'd13425,17'd12021,17'd11873,17'd11874,17'd11595,17'd11595,17'd9949,17'd9949,17'd12777,17'd9795,17'd11192,17'd9795,17'd12777,17'd11054,17'd9666,17'd9541,17'd9411,17'd9411,17'd9542,17'd9542,17'd11193,17'd13692,17'd11195,17'd9955,17'd8181,17'd8181,17'd9956,17'd10256,17'd9120,17'd12491,17'd12642,17'd11332,17'd12493,17'd10910,17'd10081,17'd8952,17'd4559,17'd2906,17'd4714,17'd4714,17'd8185,17'd8185,17'd11062,17'd2409,17'd193,17'd1382,17'd419,17'd600
},
'{
17'd1967,17'd1689,17'd1688,17'd2422,17'd7545,17'd7545,17'd2422,17'd2422,17'd1689,17'd14,17'd12,17'd806,17'd23,17'd5,17'd5205,17'd5205,17'd8040,17'd8040,17'd8340,17'd8340,17'd8340,17'd8340,17'd8340,17'd8340,17'd8340,17'd8340,17'd10537,17'd12648,17'd8195,17'd9673,17'd7713,17'd11730,17'd13693,17'd6099,17'd6106,17'd10662,17'd6272,17'd7057,17'd8973,17'd6435,17'd7223,17'd7223,17'd8825,17'd13182,17'd6266,17'd6435,17'd6595,17'd11205,17'd13576,17'd6740,17'd13694,17'd13695,17'd2595,17'd1688,17'd2782,17'd3751,17'd12196,17'd11888,17'd471,17'd294,17'd2261,17'd13696,17'd13578,17'd2430,17'd3756,17'd11210,17'd12336,17'd13579,17'd5058,17'd4255,17'd4094,17'd3262,17'd1710,17'd2442,17'd13697,17'd2276,17'd13698,17'd13699,17'd13700,17'd13701,17'd13702,17'd13703,17'd13704,17'd13589,17'd13705,17'd13706,17'd12804,17'd13707,17'd13708,17'd13709,17'd13710,17'd13711,17'd13712,17'd13713,17'd13714,17'd12951,17'd13091,17'd13206,17'd13715,17'd12212,17'd13596,17'd13716,17'd13717,17'd13718,17'd13463,17'd13598,17'd12954,17'd13093,17'd12814,17'd12360,17'd11763,17'd13719,17'd13720,17'd11764,17'd11914,17'd11914,17'd11914,17'd12066,17'd10427,17'd10563,17'd12533,17'd9701,17'd9573,17'd8537,17'd12534,17'd9007,17'd9301,17'd12959,17'd13467,17'd13466,17'd13721,17'd13721,17'd13470,17'd13469,17'd13722,17'd7578,17'd13723,17'd13724,17'd13725,17'd13726,17'd13727,17'd13478,17'd13728,17'd13729,17'd13730,17'd11483,17'd11483,17'd13731,17'd10433,17'd13732,17'd13733,17'd7265,17'd9021,17'd11240,17'd11365,17'd11366,17'd10819,17'd13734,17'd13735,17'd13736,17'd13737,17'd13738,17'd13739,17'd13740,17'd12967,17'd13741,17'd12969,17'd13621,17'd13742,17'd13344,17'd13743,17'd11776,17'd13744,17'd13745,17'd13746,17'd13747,17'd13748,17'd12394,17'd13238,17'd13495,17'd13123,17'd13749,17'd13631,17'd13242,17'd13243,17'd13750,17'd13751,17'd13500,17'd13634,17'd13635,17'd13752,17'd13753,17'd13754,17'd12088,17'd12242,17'd12402,17'd13755,17'd13756,17'd13757,17'd13758,17'd13759,17'd13760,17'd12417,17'd12859,17'd12997,17'd12256,17'd12856,17'd12575,17'd12110,17'd13761,17'd11806,17'd13362,17'd11129,17'd11965,17'd13762,17'd12996,17'd12419,17'd12580,17'd13517,17'd12418,17'd12997,17'd12859,17'd12856,17'd12856,17'd13763,17'd12111,17'd13764,17'd13138,17'd10330,17'd9480,17'd9040,17'd8415,17'd13765,17'd12266,17'd13766,17'd13767,17'd13768,17'd7954,17'd7619,17'd13769,17'd13770,17'd13771,17'd13772,17'd8740,17'd13009,17'd13773,17'd13774,17'd11819,17'd13381,17'd13775,17'd10036,17'd13533,17'd12874,17'd13776,17'd11152,17'd13777,17'd8132,17'd8132,17'd11413,17'd11413,17'd3025,17'd1197,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd133,17'd133,17'd132,17'd131,17'd6691,17'd11822,17'd13658,17'd13778,17'd13779,17'd13780,17'd13781,17'd13782,17'd13783,17'd13784,17'd13785,17'd13786,17'd13787,17'd13788,17'd13668,17'd13789,17'd13790,17'd13791,17'd10373,17'd13670,17'd13792,17'd13793,17'd8765,17'd8765,17'd12611,17'd11994,17'd12452,17'd12451,17'd13159,17'd8456,17'd12283,17'd12282,17'd12138,17'd11296,17'd7994,17'd7996,17'd8627,17'd8930,17'd8627,17'd8930,17'd9392,17'd9392,17'd9087,17'd9237,17'd9391,17'd9086,17'd9391,17'd9391,17'd9391,17'd9238,17'd9089,17'd7829,17'd7829,17'd7830,17'd13794,17'd13794,17'd13795,17'd9236,17'd9655,17'd9655,17'd9654,17'd9085,17'd9388,17'd9652,17'd9651,17'd9518,17'd9518,17'd9384,17'd10227,17'd12155,17'd12155,17'd12296,17'd12000,17'd11843,17'd11843,17'd12000,17'd12154,17'd12295,17'd11843,17'd11843,17'd11843,17'd11843,17'd11843,17'd11843,17'd11843,17'd11843,17'd12154,17'd12460,17'd12295,17'd11843,17'd13796,17'd13554,17'd13797,17'd13798,17'd13798,17'd13797,17'd13043,17'd13164,17'd13799,17'd13557,17'd13556,17'd13558,17'd12622,17'd12467,17'd13800,17'd13678,17'd13801,17'd13559,17'd13559,17'd13408,17'd13802,17'd7670,17'd8306,17'd7330,17'd7505,17'd13680,17'd13681,17'd13285,17'd13803,17'd13804,17'd13805,17'd13806,17'd13807,17'd13808,17'd13570,17'd13056,17'd13176,17'd4730,17'd6415,17'd602,17'd415,17'd13809,17'd1390,17'd1388,17'd3716,17'd3575,17'd6243,17'd6724,17'd7029,17'd7686,17'd7856,17'd8171,17'd8491,17'd9405,17'd13810,17'd10077,17'd11872,17'd13423,17'd13424,17'd13811,17'd13691,17'd12021,17'd11873,17'd11724,17'd11874,17'd11595,17'd9949,17'd9949,17'd12777,17'd9795,17'd11192,17'd9795,17'd12777,17'd11725,17'd9666,17'd9541,17'd12920,17'd12778,17'd9542,17'd9542,17'd13692,17'd13692,17'd8027,17'd7867,17'd8181,17'd7698,17'd8181,17'd9799,17'd9956,17'd12490,17'd12642,17'd12182,17'd11332,17'd10910,17'd10793,17'd9413,17'd3570,17'd2906,17'd5183,17'd4714,17'd5630,17'd5630,17'd11062,17'd603,17'd1381,17'd2256,17'd2932,17'd1528
},
'{
17'd1689,17'd3250,17'd2422,17'd3252,17'd5508,17'd7545,17'd2422,17'd1688,17'd14,17'd2,17'd12,17'd2933,17'd23,17'd6,17'd5205,17'd5205,17'd8040,17'd8340,17'd8340,17'd8340,17'd8340,17'd8340,17'd8340,17'd8340,17'd8040,17'd8340,17'd10658,17'd12648,17'd13812,17'd13813,17'd5796,17'd13814,17'd13814,17'd11730,17'd5965,17'd8669,17'd9137,17'd8518,17'd6596,17'd13182,17'd7223,17'd8973,17'd8973,17'd6596,17'd6596,17'd9136,17'd6733,17'd6594,17'd13815,17'd13816,17'd13817,17'd12647,17'd466,17'd1689,17'd2934,17'd4086,17'd12653,17'd12504,17'd471,17'd811,17'd13818,17'd13818,17'd2939,17'd12198,17'd3434,17'd12336,17'd5974,17'd13819,17'd13820,17'd13439,17'd3262,17'd996,17'd2792,17'd13821,17'd13822,17'd3610,17'd5986,17'd13823,17'd13824,17'd13825,17'd13826,17'd13827,17'd13828,17'd13449,17'd13829,17'd13830,17'd13085,17'd13831,17'd13832,17'd13202,17'd13833,17'd13834,17'd13835,17'd12674,17'd13836,17'd13091,17'd13206,17'd12212,17'd13595,17'd13837,17'd13838,17'd13718,17'd13839,17'd13598,17'd13463,17'd12954,17'd12813,17'd11626,17'd12814,17'd13840,17'd11478,17'd11478,17'd11764,17'd11913,17'd11914,17'd10690,17'd11914,17'd13841,17'd10427,17'd10286,17'd9701,17'd7418,17'd8537,17'd9300,17'd9007,17'd9575,17'd12959,17'd13466,17'd13842,17'd13466,17'd13843,17'd13844,17'd13845,17'd13846,17'd7410,17'd13847,17'd13848,17'd13849,17'd13850,17'd13851,17'd13477,17'd13852,17'd13728,17'd13853,17'd13854,17'd11484,17'd10433,17'd10700,17'd10569,17'd9015,17'd13612,17'd7266,17'd13614,17'd11365,17'd11366,17'd13855,17'd13856,17'd13857,17'd13858,17'd13859,17'd13860,17'd13861,17'd13862,17'd13863,17'd13619,17'd13864,17'd13113,17'd13343,17'd13114,17'd13865,17'd12080,17'd13866,17'd13745,17'd13867,17'd13868,17'd13869,17'd13237,17'd13238,17'd13870,17'd13871,17'd13872,17'd11500,17'd13873,17'd13874,17'd13875,17'd13633,17'd13633,17'd13500,17'd13635,17'd13502,17'd13752,17'd13876,17'd13877,17'd12710,17'd12402,17'd12851,17'd13878,17'd13879,17'd13880,17'd12717,17'd13881,17'd13519,17'd13517,17'd12997,17'd12860,17'd12418,17'd12257,17'd12110,17'd13882,17'd13883,17'd13135,17'd13762,17'd11129,17'd11129,17'd11964,17'd11807,17'd11961,17'd12580,17'd13517,17'd12418,17'd13884,17'd12859,17'd12856,17'd12575,17'd13763,17'd12718,17'd13885,17'd13886,17'd11671,17'd13887,17'd8568,17'd13888,17'd13889,17'd8426,17'd13890,17'd13891,17'd13892,17'd7790,17'd13893,17'd7458,17'd13894,17'd13771,17'd13772,17'd13895,17'd12870,17'd13896,17'd13774,17'd13897,17'd13898,17'd13775,17'd10036,17'd13533,17'd12874,17'd13899,17'd13900,17'd13901,17'd8132,17'd8132,17'd11413,17'd11413,17'd1197,17'd1197,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd133,17'd132,17'd132,17'd131,17'd13902,17'd13903,17'd13904,17'd13905,17'd13906,17'd13907,17'd13908,17'd13909,17'd13910,17'd13911,17'd13912,17'd13794,17'd9079,17'd13788,17'd13668,17'd13669,17'd13913,17'd13914,17'd10506,17'd13915,17'd13916,17'd13917,17'd8765,17'd8765,17'd12611,17'd11994,17'd12452,17'd12451,17'd13159,17'd13159,17'd8456,17'd12282,17'd12282,17'd12138,17'd8456,17'd7995,17'd7997,17'd8466,17'd8626,17'd8467,17'd8301,17'd9521,17'd9237,17'd9391,17'd9237,17'd9237,17'd9391,17'd13918,17'd9088,17'd7498,17'd9766,17'd9371,17'd10501,17'd7497,17'd8148,17'd13665,17'd13919,17'd13795,17'd9236,17'd9655,17'd9655,17'd9654,17'd10895,17'd9388,17'd9929,17'd9781,17'd9651,17'd9518,17'd9384,17'd10227,17'd12297,17'd12155,17'd12001,17'd12000,17'd12001,17'd11843,17'd12001,17'd12154,17'd12000,17'd12001,17'd11843,17'd11843,17'd12001,17'd12001,17'd11843,17'd11843,17'd12001,17'd12154,17'd12460,17'd12295,17'd13920,17'd13796,17'd13798,17'd13921,17'd13921,17'd13798,17'd13277,17'd13922,17'd13923,17'd13924,17'd13557,17'd13557,17'd13925,17'd12622,17'd12760,17'd12160,17'd13679,17'd12163,17'd13926,17'd13559,17'd13408,17'd12165,17'd8305,17'd8157,17'd7841,17'd7505,17'd13411,17'd13284,17'd13564,17'd13927,17'd13928,17'd13929,17'd13930,17'd13931,17'd13687,17'd13932,17'd13572,17'd13933,17'd4728,17'd2409,17'd1529,17'd13573,17'd1108,17'd1389,17'd1817,17'd3402,17'd5946,17'd6576,17'd6873,17'd7029,17'd7856,17'd8171,17'd8170,17'd8491,17'd13934,17'd13935,17'd13936,17'd11872,17'd12489,17'd13937,17'd13691,17'd13425,17'd12021,17'd12021,17'd11724,17'd11595,17'd9949,17'd9256,17'd9795,17'd9795,17'd11192,17'd11192,17'd9795,17'd11725,17'd11054,17'd9666,17'd13938,17'd12778,17'd9542,17'd9542,17'd13692,17'd8325,17'd8964,17'd9259,17'd8181,17'd7698,17'd8181,17'd9799,17'd10256,17'd12322,17'd12642,17'd12492,17'd13939,17'd12492,17'd8656,17'd10530,17'd9670,17'd5183,17'd5183,17'd4714,17'd3073,17'd5630,17'd11337,17'd1668,17'd952,17'd13940,17'd203,17'd4731
},
'{
17'd3250,17'd3250,17'd2422,17'd2935,17'd4246,17'd7545,17'd3250,17'd1689,17'd14,17'd12,17'd806,17'd2933,17'd4,17'd6,17'd5205,17'd5205,17'd8340,17'd8339,17'd8340,17'd8340,17'd8340,17'd8340,17'd8340,17'd8340,17'd8040,17'd10795,17'd10658,17'd12648,17'd9806,17'd8195,17'd7050,17'd13693,17'd13941,17'd13942,17'd6428,17'd8518,17'd9136,17'd6596,17'd6596,17'd8670,17'd7223,17'd6900,17'd7223,17'd5964,17'd12651,17'd9133,17'd9550,17'd10403,17'd9270,17'd10543,17'd1830,17'd2595,17'd466,17'd1831,17'd3427,17'd13943,17'd13944,17'd13945,17'd295,17'd13946,17'd13947,17'd13303,17'd13948,17'd13949,17'd13950,17'd13068,17'd13951,17'd13188,17'd13952,17'd3262,17'd1145,17'd13953,17'd13954,17'd13955,17'd13956,17'd5673,17'd13957,17'd13958,17'd13959,17'd13960,17'd13961,17'd13962,17'd13963,17'd13964,17'd12053,17'd11905,17'd13965,17'd13966,17'd12946,17'd13455,17'd13967,17'd12949,17'd12211,17'd12950,17'd13090,17'd13091,17'd13206,17'd13326,17'd13595,17'd13837,17'd13838,17'd13839,17'd13968,17'd13598,17'd13209,17'd13093,17'd13093,17'd13094,17'd12530,17'd11478,17'd11478,17'd11764,17'd13969,17'd12361,17'd12680,17'd11914,17'd12066,17'd13841,17'd13327,17'd8687,17'd9573,17'd8537,17'd9159,17'd9007,17'd9575,17'd13468,17'd13466,17'd13466,17'd13842,17'd13970,17'd13971,17'd13972,17'd13722,17'd6929,17'd13973,17'd13974,17'd13975,17'd13976,17'd13977,17'd13978,17'd13979,17'd13852,17'd13334,17'd13980,17'd10568,17'd10700,17'd10700,17'd9849,17'd9309,17'd13611,17'd12686,17'd9021,17'd11632,17'd11768,17'd13855,17'd11485,17'd13981,17'd13982,17'd13983,17'd13737,17'd13861,17'd13738,17'd13984,17'd13985,17'd13340,17'd13620,17'd13113,17'd13343,17'd12691,17'd13986,17'd13987,17'd13988,17'd13867,17'd13747,17'd13869,17'd13989,17'd13990,17'd13495,17'd13991,17'd13992,17'd13993,17'd13352,17'd12699,17'd13875,17'd13994,17'd13498,17'd13498,17'd13501,17'd13995,17'd13996,17'd13753,17'd12568,17'd12710,17'd13997,17'd13998,17'd13360,17'd13999,17'd14000,17'd14001,17'd12109,17'd12718,17'd14002,17'd13365,17'd12997,17'd12415,17'd14003,17'd12110,17'd12111,17'd13882,17'd13135,17'd11807,17'd11807,17'd11965,17'd11131,17'd10989,17'd11807,17'd11961,17'd12419,17'd12995,17'd12418,17'd13884,17'd12859,17'd12417,17'd12575,17'd13763,17'd12718,17'd13137,17'd10476,17'd11277,17'd9039,17'd14004,17'd14005,17'd14006,17'd14007,17'd14008,17'd14009,17'd8258,17'd14010,17'd14011,17'd14012,17'd12121,17'd14013,17'd14014,17'd8589,17'd12870,17'd13896,17'd13774,17'd13380,17'd14015,17'd13775,17'd10036,17'd13533,17'd11977,17'd13776,17'd14016,17'd14017,17'd11289,17'd11289,17'd11413,17'd11413,17'd1197,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd357,17'd14018,17'd14019,17'd10624,17'd14020,17'd14021,17'd14022,17'd14023,17'd14024,17'd14025,17'd14026,17'd14027,17'd14028,17'd14029,17'd14030,17'd13668,17'd14031,17'd13547,17'd14032,17'd13915,17'd14033,17'd14034,17'd10211,17'd8616,17'd8765,17'd12611,17'd11994,17'd12452,17'd12451,17'd13159,17'd13159,17'd14035,17'd12896,17'd8457,17'd12282,17'd8456,17'd7994,17'd7995,17'd7994,17'd14036,17'd7829,17'd7829,17'd8300,17'd14037,17'd14037,17'd13673,17'd13673,17'd13673,17'd7834,17'd7835,17'd9221,17'd9639,17'd14038,17'd14038,17'd14038,17'd9505,17'd7497,17'd14039,17'd13919,17'd14040,17'd14041,17'd13675,17'd14042,17'd10896,17'd10896,17'd14043,17'd9653,17'd9929,17'd14044,17'd9651,17'd9780,17'd12155,17'd11844,17'd11843,17'd12154,17'd12154,17'd12001,17'd11843,17'd12001,17'd12154,17'd12000,17'd12001,17'd12001,17'd12001,17'd12001,17'd12001,17'd11843,17'd12900,17'd12618,17'd12460,17'd12899,17'd12154,17'd11845,17'd13796,17'd13797,17'd13921,17'd13796,17'd13796,17'd13921,17'd13923,17'd13923,17'd13924,17'd13556,17'd14045,17'd14046,17'd14047,17'd14048,17'd14049,17'd14050,17'd14051,17'd13559,17'd13168,17'd13047,17'd6560,17'd14052,17'd7331,17'd7505,17'd13283,17'd13284,17'd14053,17'd14054,17'd14055,17'd14056,17'd14057,17'd14058,17'd14059,17'd13688,17'd13689,17'd14060,17'd4882,17'd2393,17'd1529,17'd195,17'd14061,17'd2751,17'd2913,17'd3403,17'd4720,17'd7193,17'd7030,17'd7029,17'd8169,17'd8171,17'd8170,17'd8491,17'd14062,17'd13690,17'd10077,17'd12487,17'd12178,17'd12178,17'd13691,17'd13425,17'd12021,17'd13425,17'd11873,17'd11874,17'd9949,17'd9256,17'd9795,17'd9795,17'd9795,17'd11192,17'd14063,17'd14064,17'd14065,17'd8807,17'd13938,17'd12920,17'd8324,17'd12921,17'd7691,17'd8026,17'd8964,17'd8027,17'd7867,17'd8327,17'd7698,17'd9955,17'd10256,17'd9120,17'd12642,17'd12642,17'd10256,17'd12182,17'd10910,17'd11880,17'd12494,17'd6581,17'd5183,17'd4714,17'd6889,17'd6415,17'd781,17'd1668,17'd1409,17'd14066,17'd1244,17'd1244
},
'{
17'd2422,17'd2422,17'd2935,17'd2935,17'd4246,17'd4887,17'd2781,17'd1127,17'd0,17'd12,17'd806,17'd4242,17'd5,17'd6,17'd5205,17'd5205,17'd8340,17'd8339,17'd8340,17'd8340,17'd8340,17'd8340,17'd8340,17'd8340,17'd8040,17'd10795,17'd10537,17'd7727,17'd9961,17'd14067,17'd14068,17'd7553,17'd7381,17'd13942,17'd6099,17'd9135,17'd6596,17'd6435,17'd8973,17'd8670,17'd8973,17'd7058,17'd6434,17'd6102,17'd9133,17'd9132,17'd10403,17'd6734,17'd6103,17'd14069,17'd4247,17'd4247,17'd4247,17'd14070,17'd3427,17'd14071,17'd14072,17'd14073,17'd659,17'd14074,17'd14075,17'd2262,17'd14076,17'd13949,17'd14077,17'd5805,17'd14078,17'd14079,17'd14080,17'd831,17'd14081,17'd2442,17'd14082,17'd14083,17'd4591,17'd14084,17'd14085,17'd14086,17'd14087,17'd14088,17'd14089,17'd14090,17'd14091,17'd14092,17'd12053,17'd13084,17'd13965,17'd14093,17'd12805,17'd14094,17'd14095,17'd14096,17'd13322,17'd13089,17'd13090,17'd14097,17'd12212,17'd13326,17'd13596,17'd13838,17'd14098,17'd13462,17'd13463,17'd13092,17'd13093,17'd11626,17'd13094,17'd12956,17'd11913,17'd11764,17'd11764,17'd11764,17'd12361,17'd12361,17'd11913,17'd12066,17'd13841,17'd10286,17'd8687,17'd9573,17'd8537,17'd10694,17'd9007,17'd9575,17'd13468,17'd14099,17'd14100,17'd14100,17'd13467,17'd13970,17'd13469,17'd6134,17'd14101,17'd14102,17'd14103,17'd14104,17'd14105,17'd13976,17'd14106,17'd14107,17'd13852,17'd13979,17'd14108,17'd13730,17'd10569,17'd9992,17'd9992,17'd14109,17'd9016,17'd8548,17'd13222,17'd7926,17'd11365,17'd12222,17'd13223,17'd10820,17'd13107,17'd14110,17'd13737,17'd14111,17'd13738,17'd14112,17'd14113,17'd14114,17'd13227,17'd13620,17'd13342,17'd13343,17'd12691,17'd14115,17'd14116,17'd14117,17'd14118,17'd13869,17'd12396,17'd12238,17'd13240,17'd13991,17'd13992,17'd14119,17'd13631,17'd14120,17'd13875,17'd14121,17'd13994,17'd14122,17'd14123,17'd14124,17'd12706,17'd14125,17'd12400,17'd12243,17'd11791,17'd14126,17'd14127,17'd14128,17'd14129,17'd12413,17'd14130,17'd11959,17'd13363,17'd12113,17'd13763,17'd12855,17'd12416,17'd14003,17'd12110,17'd12111,17'd14131,17'd13135,17'd11807,17'd11807,17'd11808,17'd14132,17'd11129,17'd11807,17'd11961,17'd13761,17'd12109,17'd12418,17'd13884,17'd12859,17'd12417,17'd12418,17'd12856,17'd13882,17'd14133,17'd14134,17'd11277,17'd9038,17'd14135,17'd14136,17'd7457,17'd14137,17'd14138,17'd14139,17'd13654,17'd14140,17'd8259,17'd14141,17'd12121,17'd14142,17'd14143,17'd8589,17'd14144,17'd13896,17'd13774,17'd14145,17'd13898,17'd13775,17'd10036,17'd13533,17'd11977,17'd13899,17'd13900,17'd14017,17'd11289,17'd11289,17'd11413,17'd11413,17'd1197,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd135,17'd131,17'd14146,17'd14147,17'd13904,17'd14148,17'd14021,17'd13265,17'd14149,17'd14150,17'd14151,17'd14152,17'd14153,17'd14040,17'd9079,17'd14030,17'd13668,17'd13669,17'd14154,17'd14032,17'd14155,17'd14156,17'd14157,17'd13792,17'd8616,17'd8616,17'd8457,17'd11994,17'd12452,17'd12451,17'd13159,17'd13159,17'd14035,17'd12611,17'd8295,17'd8615,17'd8614,17'd8614,17'd7994,17'd7994,17'd8613,17'd7834,17'd13673,17'd14037,17'd13673,17'd7830,17'd8300,17'd13673,17'd7828,17'd10501,17'd9221,17'd9370,17'd14038,17'd14158,17'd14159,17'd14160,17'd14161,17'd9640,17'd7497,17'd14039,17'd13919,17'd14040,17'd9236,17'd13675,17'd14162,17'd11033,17'd14162,17'd10896,17'd9388,17'd9929,17'd9781,17'd10063,17'd10377,17'd11846,17'd11844,17'd12001,17'd12154,17'd12460,17'd12154,17'd11843,17'd12295,17'd12000,17'd12001,17'd12001,17'd12001,17'd12001,17'd12001,17'd12001,17'd12617,17'd12618,17'd12154,17'd12460,17'd12460,17'd12000,17'd14163,17'd13797,17'd13921,17'd14164,17'd14164,17'd13921,17'd13923,17'd14165,17'd13799,17'd13557,17'd14045,17'd14046,17'd14045,17'd13045,17'd14166,17'd12760,17'd12622,17'd12162,17'd12162,17'd14167,17'd14168,17'd9395,17'd7331,17'd7503,17'd13680,17'd13681,17'd14169,17'd14170,17'd14055,17'd14171,17'd14172,17'd14173,17'd14174,17'd14175,17'd14176,17'd14177,17'd5958,17'd14178,17'd1529,17'd600,17'd14179,17'd5778,17'd2914,17'd3876,17'd3575,17'd7031,17'd8497,17'd6873,17'd8169,17'd8018,17'd7855,17'd7855,17'd14180,17'd13934,17'd13690,17'd12487,17'd11723,17'd12178,17'd13691,17'd13425,17'd13425,17'd13425,17'd12021,17'd11724,17'd9256,17'd9256,17'd9795,17'd9795,17'd9795,17'd9795,17'd14063,17'd14064,17'd14181,17'd8807,17'd13938,17'd13938,17'd12778,17'd8324,17'd7691,17'd8026,17'd8179,17'd8964,17'd8326,17'd8028,17'd7874,17'd8181,17'd10256,17'd9956,17'd12492,17'd12642,17'd9956,17'd9120,17'd8503,17'd12324,17'd9669,17'd6727,17'd5183,17'd4714,17'd6889,17'd8185,17'd14182,17'd1668,17'd1955,17'd1685,17'd1244,17'd1244
},
'{
17'd2784,17'd2935,17'd4246,17'd4887,17'd4887,17'd7711,17'd1689,17'd1127,17'd1,17'd806,17'd2933,17'd2421,17'd6,17'd5205,17'd5205,17'd8340,17'd8339,17'd8339,17'd8340,17'd10795,17'd8190,17'd8190,17'd8190,17'd8190,17'd5205,17'd8190,17'd14183,17'd14184,17'd7894,17'd9263,17'd807,17'd14185,17'd5798,17'd11730,17'd7713,17'd5796,17'd6266,17'd7223,17'd8670,17'd8670,17'd6900,17'd6900,17'd5965,17'd6104,17'd8342,17'd14186,17'd9680,17'd8983,17'd14187,17'd1830,17'd1688,17'd1688,17'd10535,17'd14188,17'd10924,17'd12653,17'd14189,17'd14190,17'd1279,17'd14191,17'd984,17'd470,17'd12198,17'd3259,17'd14192,17'd4253,17'd14193,17'd14194,17'd2788,17'd14195,17'd14196,17'd13954,17'd13955,17'd14197,17'd5673,17'd14198,17'd14199,17'd14200,17'd14201,17'd14202,17'd14090,17'd14203,17'd14204,17'd14205,17'd14206,17'd14207,17'd13831,17'd14208,17'd14209,17'd14210,17'd14096,17'd14211,17'd14212,17'd14213,17'd14214,17'd14215,17'd13459,17'd13326,17'd13460,17'd14216,17'd14217,17'd13462,17'd13598,17'd12954,17'd13093,17'd12065,17'd12218,17'd11627,17'd11764,17'd11629,17'd12532,17'd12532,17'd12362,17'd12361,17'd11913,17'd11764,17'd11629,17'd10427,17'd10286,17'd9158,17'd9159,17'd14218,17'd9301,17'd9575,17'd13466,17'd14100,17'd14219,17'd14219,17'd14220,17'd13470,17'd14221,17'd6301,17'd14222,17'd14223,17'd14224,17'd14225,17'd14105,17'd14226,17'd14227,17'd14107,17'd14228,17'd14228,17'd13980,17'd14229,17'd10700,17'd14230,17'd12822,17'd9016,17'd14231,17'd7590,17'd9169,17'd13614,17'd11768,17'd11769,17'd14232,17'd14233,17'd14234,17'd13983,17'd14111,17'd13861,17'd14235,17'd14236,17'd14237,17'd14238,17'd14239,17'd14240,17'd13342,17'd13343,17'd12833,17'd12693,17'd14241,17'd14242,17'd14243,17'd14244,17'd14245,17'd14246,17'd14247,17'd14248,17'd13630,17'd13241,17'd14249,17'd14250,17'd13875,17'd14121,17'd14251,17'd14252,17'd13635,17'd14253,17'd12706,17'd13130,17'd13129,17'd13507,17'd14254,17'd14255,17'd14256,17'd14257,17'd12111,17'd14258,17'd14259,17'd14260,17'd14261,17'd11960,17'd12109,17'd12575,17'd12575,17'd12575,17'd12109,17'd12580,17'd13882,17'd11806,17'd11807,17'd14262,17'd11131,17'd14263,17'd10989,17'd11667,17'd13363,17'd13882,17'd12109,17'd12253,17'd12997,17'd12859,17'd12417,17'd12418,17'd12579,17'd14130,17'd14264,17'd12584,17'd11277,17'd8873,17'd8100,17'd7787,17'd7622,17'd14265,17'd14266,17'd14267,17'd14268,17'd14140,17'd14269,17'd14270,17'd12121,17'd14271,17'd12122,17'd8589,17'd14272,17'd13896,17'd13774,17'd11819,17'd10616,17'd14273,17'd14274,17'd13533,17'd11977,17'd14275,17'd14276,17'd14017,17'd11289,17'd8132,17'd11413,17'd1045,17'd1197,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd135,17'd131,17'd14146,17'd4340,17'd14277,17'd14278,17'd14279,17'd14280,17'd14281,17'd14282,17'd14283,17'd14284,17'd14285,17'd14286,17'd14029,17'd14030,17'd13546,17'd14031,17'd13547,17'd14032,17'd14155,17'd14287,17'd14288,17'd14289,17'd14290,17'd14290,17'd8457,17'd11994,17'd12451,17'd13159,17'd13159,17'd12451,17'd12896,17'd12611,17'd8457,17'd8615,17'd12138,17'd12282,17'd8614,17'd13672,17'd8612,17'd8293,17'd8153,17'd8153,17'd8300,17'd7830,17'd7830,17'd7830,17'd14291,17'd10047,17'd9370,17'd14038,17'd14292,17'd14293,17'd14294,17'd14295,17'd14296,17'd14297,17'd9640,17'd11296,17'd14036,17'd13919,17'd13795,17'd14298,17'd14299,17'd13795,17'd14153,17'd14285,17'd10896,17'd14043,17'd9653,17'd9652,17'd10223,17'd14300,17'd11845,17'd11843,17'd12154,17'd12899,17'd12460,17'd12000,17'd12295,17'd12154,17'd12000,17'd12001,17'd12001,17'd12001,17'd12000,17'd12000,17'd12618,17'd12618,17'd12000,17'd12154,17'd12460,17'd12295,17'd13920,17'd13921,17'd13796,17'd14164,17'd14164,17'd13796,17'd13796,17'd14164,17'd13923,17'd13924,17'd13042,17'd13277,17'd13277,17'd13165,17'd11852,17'd14048,17'd14301,17'd12162,17'd12162,17'd12163,17'd14302,17'd14303,17'd6712,17'd7503,17'd14304,17'd13681,17'd14169,17'd14170,17'd14305,17'd14306,17'd14307,17'd14308,17'd14058,17'd14309,17'd14310,17'd14311,17'd14312,17'd14178,17'd1529,17'd416,17'd599,17'd1106,17'd2750,17'd1816,17'd4408,17'd5946,17'd6577,17'd7030,17'd7685,17'd8169,17'd8018,17'd7855,17'd14313,17'd14062,17'd13810,17'd11593,17'd11723,17'd12178,17'd13425,17'd13425,17'd13691,17'd13425,17'd12021,17'd11873,17'd10249,17'd9256,17'd9795,17'd9795,17'd9795,17'd9795,17'd14063,17'd14064,17'd14065,17'd8807,17'd13938,17'd13938,17'd13938,17'd12778,17'd7691,17'd8026,17'd8179,17'd8179,17'd8027,17'd8028,17'd7874,17'd8181,17'd10256,17'd10256,17'd12492,17'd12642,17'd9120,17'd9956,17'd8503,17'd14314,17'd13060,17'd9670,17'd5183,17'd5183,17'd6889,17'd5372,17'd1394,17'd1668,17'd1409,17'd971,17'd14315,17'd14316
},
'{
17'd2593,17'd2935,17'd4887,17'd4887,17'd4577,17'd6583,17'd1689,17'd1127,17'd3,17'd1275,17'd4242,17'd7215,17'd3753,17'd5205,17'd8190,17'd8340,17'd8339,17'd8339,17'd10795,17'd10795,17'd8190,17'd8190,17'd8190,17'd8190,17'd5205,17'd8190,17'd14183,17'd9672,17'd8196,17'd978,17'd977,17'd6587,17'd14317,17'd5796,17'd7893,17'd6098,17'd7713,17'd7223,17'd9136,17'd8815,17'd14318,17'd8973,17'd6102,17'd9551,17'd8822,17'd6740,17'd6430,17'd8823,17'd14319,17'd466,17'd1689,17'd3750,17'd3252,17'd3101,17'd2783,17'd14320,17'd14321,17'd14322,17'd14323,17'd2429,17'd2430,17'd12198,17'd14324,17'd14325,17'd2431,17'd14326,17'd14194,17'd480,17'd14327,17'd670,17'd2271,17'd14082,17'd14083,17'd4591,17'd14084,17'd14328,17'd14329,17'd14330,17'd14331,17'd14332,17'd14333,17'd14334,17'd14335,17'd12208,17'd13706,17'd14336,17'd14337,17'd14338,17'd12056,17'd14339,17'd14340,17'd14097,17'd14341,17'd14214,17'd14342,17'd14343,17'd13595,17'd12675,17'd13460,17'd14344,17'd13462,17'd13092,17'd12954,17'd12813,17'd12813,17'd13094,17'd11627,17'd11764,17'd11764,17'd12531,17'd12531,17'd12531,17'd12680,17'd11913,17'd11764,17'd11361,17'd10691,17'd13327,17'd9158,17'd9159,17'd10430,17'd9301,17'd12959,17'd13468,17'd14099,17'd14345,17'd14346,17'd14347,17'd13971,17'd13845,17'd6301,17'd6622,17'd14348,17'd14349,17'd14350,17'd14351,17'd13976,17'd14352,17'd14353,17'd14354,17'd14354,17'd14355,17'd14356,17'd14357,17'd14358,17'd14230,17'd9016,17'd14359,17'd12686,17'd7925,17'd9171,17'd14360,17'd11366,17'd13855,17'd9854,17'd13107,17'd13339,17'd13737,17'd14361,17'd14361,17'd14112,17'd14362,17'd13985,17'd14363,17'd14364,17'd13228,17'd13229,17'd12691,17'd12834,17'd14365,17'd14117,17'd14118,17'd13631,17'd12395,17'd14366,17'd14367,17'd14368,17'd14369,17'd14370,17'd14249,17'd14371,17'd14123,17'd14123,17'd14123,17'd14251,17'd14252,17'd14372,17'd14373,17'd14125,17'd14374,17'd13359,17'd14375,17'd13639,17'd14256,17'd14376,17'd14377,17'd13645,17'd14378,17'd14379,17'd14380,17'd13883,17'd12419,17'd12856,17'd12856,17'd12575,17'd12575,17'd12414,17'd12109,17'd13363,17'd11806,17'd11807,17'd11965,17'd14381,17'd11130,17'd11395,17'd13764,17'd13364,17'd12110,17'd12109,17'd12418,17'd12997,17'd12859,17'd12417,17'd12418,17'd12253,17'd14130,17'd14382,17'd12584,17'd14383,17'd9041,17'd14384,17'd14385,17'd8109,17'd14386,17'd14387,17'd14388,17'd14389,17'd14390,17'd14391,17'd14392,17'd12121,17'd14393,17'd14394,17'd14395,17'd14272,17'd14396,17'd14397,17'd11819,17'd14398,17'd14273,17'd14274,17'd14399,17'd14400,17'd14275,17'd14016,17'd14401,17'd8132,17'd8132,17'd11413,17'd1045,17'd1197,17'd1197,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd14146,17'd14402,17'd14403,17'd14404,17'd14279,17'd14405,17'd14406,17'd14407,17'd14408,17'd14409,17'd14410,17'd14411,17'd14412,17'd14030,17'd13546,17'd13789,17'd13547,17'd14413,17'd14155,17'd14287,17'd14414,17'd14034,17'd8458,17'd14290,17'd12611,17'd12450,17'd12451,17'd13159,17'd13159,17'd8294,17'd12611,17'd12611,17'd12896,17'd14035,17'd12282,17'd12282,17'd12138,17'd12137,17'd13672,17'd7994,17'd7994,17'd7994,17'd13673,17'd14037,17'd14036,17'd8613,17'd10047,17'd9640,17'd14038,17'd14415,17'd14159,17'd14294,17'd14416,17'd14417,17'd14418,17'd14419,17'd9370,17'd8761,17'd8148,17'd13665,17'd13786,17'd14028,17'd14420,17'd14299,17'd13795,17'd14298,17'd14298,17'd14162,17'd11177,17'd9929,17'd9517,17'd10224,17'd10225,17'd12155,17'd12154,17'd12154,17'd12295,17'd12899,17'd12295,17'd12295,17'd12000,17'd12001,17'd12001,17'd12001,17'd12000,17'd12154,17'd12617,17'd12617,17'd12001,17'd12001,17'd12295,17'd12899,17'd14421,17'd14422,17'd14164,17'd14164,17'd14164,17'd14164,17'd14164,17'd13796,17'd13923,17'd13799,17'd13042,17'd13043,17'd13277,17'd13042,17'd12306,17'd12904,17'd12467,17'd14423,17'd14424,17'd12163,17'd14425,17'd14426,17'd6712,17'd7331,17'd14427,17'd13411,17'd14428,17'd14170,17'd14429,17'd14430,17'd14431,17'd14432,17'd14058,17'd14433,17'd14434,17'd14311,17'd14312,17'd6889,17'd2589,17'd419,17'd418,17'd14435,17'd1386,17'd2913,17'd3403,17'd4720,17'd6243,17'd8497,17'd7346,17'd7685,17'd8018,17'd7854,17'd14436,17'd14180,17'd13810,17'd10077,17'd12488,17'd12489,17'd12178,17'd13691,17'd13691,17'd13425,17'd12021,17'd12021,17'd11724,17'd9256,17'd9795,17'd9795,17'd9795,17'd9795,17'd14063,17'd14064,17'd14065,17'd8807,17'd13938,17'd14437,17'd13938,17'd12920,17'd7691,17'd7691,17'd8179,17'd8179,17'd8964,17'd8809,17'd14438,17'd7698,17'd10256,17'd10256,17'd12182,17'd12490,17'd8181,17'd10256,17'd8810,17'd14439,17'd13180,17'd11334,17'd8187,17'd5183,17'd3570,17'd5940,17'd10911,17'd1668,17'd1098,17'd205,17'd972,17'd1098
},
'{
17'd4733,17'd4733,17'd4733,17'd4246,17'd3252,17'd1688,17'd1127,17'd2,17'd10,17'd25,17'd4,17'd6,17'd5205,17'd8040,17'd8340,17'd8340,17'd8339,17'd8339,17'd13295,17'd8339,17'd8040,17'd8040,17'd5205,17'd5205,17'd6,17'd7,17'd7374,17'd5206,17'd8,17'd4,17'd8,17'd5647,17'd5794,17'd5794,17'd5513,17'd12649,17'd7724,17'd8825,17'd8511,17'd7057,17'd11067,17'd14440,17'd9681,17'd8982,17'd7217,17'd7051,17'd7217,17'd14441,17'd14442,17'd17,17'd466,17'd4247,17'd7545,17'd4245,17'd4736,17'd14443,17'd14444,17'd14445,17'd37,17'd14446,17'd3596,17'd3106,17'd2945,17'd14447,17'd14448,17'd14449,17'd826,17'd14450,17'd14451,17'd2270,17'd14452,17'd14453,17'd3767,17'd14454,17'd13823,17'd14455,17'd14456,17'd14331,17'd14457,17'd14458,17'd13590,17'd13706,17'd14459,17'd13706,17'd14460,17'd14208,17'd14461,17'd12210,17'd14462,17'd14463,17'd14464,17'd14097,17'd14097,17'd14097,17'd14465,17'd14343,17'd12212,17'd13460,17'd14466,17'd14467,17'd14468,17'd14469,17'd13092,17'd13093,17'd13211,17'd14470,17'd12361,17'd13969,17'd14471,17'd13840,17'd12218,17'd11360,17'd12957,17'd14472,17'd11361,17'd13841,17'd8687,17'd12220,17'd12219,17'd10430,17'd9704,17'd13842,17'd14099,17'd14100,17'd14473,17'd14474,17'd14475,17'd13467,17'd9703,17'd9300,17'd14476,17'd14477,17'd14478,17'd14479,17'd14480,17'd14481,17'd14482,17'd14483,17'd14484,17'd14485,17'd14486,17'd14357,17'd14487,17'd14488,17'd14489,17'd14109,17'd13611,17'd7265,17'd9021,17'd14490,17'd14491,17'd14492,17'd9592,17'd10437,17'd14493,17'd14494,17'd13737,17'd14495,17'd14496,17'd14497,17'd14498,17'd14499,17'd14114,17'd14500,17'd14240,17'd14501,17'd13114,17'd14502,17'd11928,17'd14503,17'd14504,17'd14505,17'd12396,17'd14506,17'd14507,17'd14508,17'd14509,17'd14510,17'd14511,17'd14371,17'd13355,17'd13246,17'd13501,17'd13127,17'd14512,17'd14512,17'd12393,17'd14513,17'd13504,17'd12094,17'd14514,17'd14515,17'd13132,17'd14516,17'd14517,17'd14518,17'd14519,17'd12584,17'd14520,17'd11960,17'd13519,17'd14521,17'd12856,17'd12575,17'd12414,17'd12109,17'd12110,17'd12718,17'd13135,17'd11962,17'd14262,17'd11129,17'd14522,17'd13645,17'd11962,17'd13363,17'd12110,17'd12414,17'd12418,17'd14523,17'd14524,17'd14525,17'd14526,17'd12256,17'd12577,17'd11961,17'd11274,17'd14134,17'd11809,17'd12118,17'd14527,17'd9351,17'd14528,17'd14529,17'd14530,17'd14010,17'd10180,17'd14531,17'd14392,17'd14532,17'd14533,17'd14393,17'd14534,17'd14535,17'd14144,17'd14536,17'd14537,17'd14538,17'd14539,17'd14540,17'd14541,17'd13533,17'd8597,17'd8444,17'd14016,17'd11152,17'd14017,17'd3025,17'd1197,17'd1197,17'd1197,17'd1197,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd131,17'd7484,17'd14542,17'd10624,17'd14543,17'd14544,17'd14545,17'd14546,17'd14547,17'd14548,17'd14549,17'd14550,17'd14551,17'd14029,17'd14552,17'd14553,17'd13548,17'd13670,17'd14033,17'd14287,17'd14554,17'd14555,17'd14556,17'd14557,17'd14558,17'd8151,17'd14559,17'd12289,17'd13159,17'd12282,17'd12282,17'd8456,17'd12451,17'd13159,17'd8456,17'd12282,17'd9767,17'd14560,17'd9506,17'd13665,17'd8300,17'd8300,17'd13673,17'd7995,17'd7833,17'd10047,17'd14038,17'd14158,17'd14158,17'd14561,17'd14562,17'd14159,17'd14160,17'd14563,17'd14564,17'd14297,17'd11423,17'd11551,17'd9639,17'd8610,17'd7497,17'd14039,17'd13393,17'd14565,17'd14039,17'd14039,17'd13786,17'd14286,17'd13795,17'd14566,17'd14567,17'd9929,17'd9652,17'd9651,17'd10226,17'd12297,17'd12295,17'd13035,17'd14568,17'd14568,17'd14569,17'd13162,17'd12900,17'd12618,17'd13162,17'd12617,17'd13162,17'd12618,17'd12618,17'd12618,17'd12900,17'd12618,17'd12899,17'd14570,17'd14571,17'd14572,17'd14573,17'd14163,17'd14164,17'd13923,17'd14165,17'd14165,17'd14165,17'd13799,17'd13677,17'd13677,17'd13923,17'd13558,17'd14166,17'd11853,17'd12467,17'd12162,17'd12163,17'd13408,17'd14574,17'd14575,17'd7331,17'd7505,17'd14576,17'd14577,17'd14170,17'd14578,17'd14305,17'd14579,17'd14580,17'd14581,17'd14582,17'd14583,17'd14584,17'd14585,17'd14312,17'd14586,17'd941,17'd14587,17'd14588,17'd2748,17'd14589,17'd3080,17'd5032,17'd7521,17'd7520,17'd6873,17'd7685,17'd14590,17'd14591,17'd14592,17'd14180,17'd8795,17'd10076,17'd12319,17'd12487,17'd11723,17'd12178,17'd13425,17'd13691,17'd14593,17'd14594,17'd14595,17'd11873,17'd14063,17'd14063,17'd12777,17'd9795,17'd9795,17'd12777,17'd11725,17'd11054,17'd11054,17'd9666,17'd13938,17'd13938,17'd8026,17'd7691,17'd13692,17'd14596,17'd8325,17'd12641,17'd7698,17'd14438,17'd9956,17'd10256,17'd9120,17'd9120,17'd7524,17'd9668,17'd10654,17'd11196,17'd10793,17'd10083,17'd9544,17'd4714,17'd4714,17'd2098,17'd1525,17'd424,17'd1685,17'd1124,17'd1687,17'd14597
},
'{
17'd3904,17'd3904,17'd6584,17'd4887,17'd2422,17'd4247,17'd2,17'd12,17'd10,17'd23,17'd6,17'd5205,17'd8040,17'd8040,17'd8340,17'd8340,17'd8339,17'd8339,17'd8339,17'd8339,17'd8040,17'd8040,17'd5205,17'd5205,17'd7,17'd7,17'd5378,17'd8,17'd4,17'd23,17'd4,17'd8,17'd5513,17'd5513,17'd7375,17'd12649,17'd13431,17'd8670,17'd8511,17'd9137,17'd10919,17'd11342,17'd9132,17'd6741,17'd7722,17'd7546,17'd6270,17'd10923,17'd9422,17'd17,17'd2595,17'd1688,17'd4246,17'd4428,17'd5202,17'd14598,17'd14322,17'd14599,17'd1553,17'd14446,17'd14600,17'd14600,17'd2606,17'd2433,17'd14601,17'd14602,17'd482,17'd14603,17'd14604,17'd2127,17'd14605,17'd2449,17'd14606,17'd14607,17'd14608,17'd14200,17'd14609,17'd14610,17'd14611,17'd14612,17'd14613,17'd14206,17'd13830,17'd14614,17'd14615,17'd14616,17'd14617,17'd12807,17'd14618,17'd14619,17'd13715,17'd13206,17'd13206,17'd13715,17'd14465,17'd13595,17'd14620,17'd14216,17'd14466,17'd14217,17'd14469,17'd13092,17'd12813,17'd13093,17'd14621,17'd14622,17'd12361,17'd13969,17'd13840,17'd12530,17'd12814,17'd12956,17'd11914,17'd10815,17'd13841,17'd10286,17'd12535,17'd12219,17'd10430,17'd9007,17'd13842,17'd14623,17'd14624,17'd14625,17'd14474,17'd14626,17'd14345,17'd13468,17'd9703,17'd9440,17'd14627,17'd14628,17'd14629,17'd14630,17'd14631,17'd14632,17'd14633,17'd14634,17'd14485,17'd14635,17'd14636,17'd14637,17'd14638,17'd14639,17'd14230,17'd9016,17'd14640,17'd12823,17'd9171,17'd14641,17'd12825,17'd9452,17'd10437,17'd14642,17'd14643,17'd14644,17'd14495,17'd14645,17'd14646,17'd14647,17'd14648,17'd14649,17'd14238,17'd14239,17'd13228,17'd14650,17'd14651,17'd14652,17'd14653,17'd14654,17'd14655,17'd12562,17'd11501,17'd14656,17'd14657,17'd14658,17'd14659,17'd14660,17'd14661,17'd14252,17'd13355,17'd13355,17'd14123,17'd14512,17'd14251,17'd12558,17'd13127,17'd14662,17'd12093,17'd12099,17'd14663,17'd12853,17'd14664,17'd14665,17'd14666,17'd14667,17'd10169,17'd14668,17'd14669,17'd11960,17'd14670,17'd14521,17'd12856,17'd12414,17'd12579,17'd12580,17'd12419,17'd12718,17'd12861,17'd11963,17'd14262,17'd11965,17'd14671,17'd13516,17'd13135,17'd13882,17'd12109,17'd12575,17'd13643,17'd14523,17'd14672,17'd14525,17'd14526,17'd12256,17'd12577,17'd11962,17'd14673,17'd11670,17'd14674,17'd14675,17'd14676,17'd13141,17'd14677,17'd14678,17'd14679,17'd14680,17'd14681,17'd14682,17'd14683,17'd14684,17'd13529,17'd7627,17'd14534,17'd14685,17'd14686,17'd14687,17'd14688,17'd14689,17'd14690,17'd14691,17'd14541,17'd14692,17'd14693,17'd14694,17'd14016,17'd10874,17'd11413,17'd3025,17'd1197,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd131,17'd4815,17'd14695,17'd14696,17'd14697,17'd14698,17'd14699,17'd14700,17'd14547,17'd14701,17'd14409,17'd14702,17'd14551,17'd14029,17'd14703,17'd14553,17'd13548,17'd13670,17'd14704,17'd14705,17'd14554,17'd14555,17'd14706,17'd12745,17'd12282,17'd12289,17'd14559,17'd12289,17'd13159,17'd12282,17'd12282,17'd8456,17'd12451,17'd13159,17'd13159,17'd12138,17'd9767,17'd11017,17'd14707,17'd13665,17'd9088,17'd8300,17'd14036,17'd7832,17'd11016,17'd14708,17'd14709,17'd14710,17'd14711,17'd14711,17'd14712,17'd14159,17'd14713,17'd14714,17'd14714,17'd14715,17'd11423,17'd11551,17'd11551,17'd11551,17'd8610,17'd14716,17'd13153,17'd14565,17'd14039,17'd14039,17'd14565,17'd13919,17'd14717,17'd14551,17'd14718,17'd14719,17'd14720,17'd9387,17'd10773,17'd12155,17'd12000,17'd12154,17'd14721,17'd14568,17'd14568,17'd14721,17'd12618,17'd12617,17'd12618,17'd14721,17'd13162,17'd13162,17'd13162,17'd12618,17'd12617,17'd12618,17'd14721,17'd14570,17'd14722,17'd14723,17'd14573,17'd14164,17'd14163,17'd14724,17'd14165,17'd13923,17'd14724,17'd13799,17'd13677,17'd13677,17'd13799,17'd13925,17'd13407,17'd14049,17'd12760,17'd12468,17'd12163,17'd13408,17'd14725,17'd14726,17'd6856,17'd7841,17'd14576,17'd14428,17'd14727,17'd14728,17'd14729,17'd14730,17'd14731,17'd14732,17'd14733,17'd14734,17'd14735,17'd14584,17'd14736,17'd4714,17'd12644,17'd1811,17'd11883,17'd14737,17'd14738,17'd2911,17'd3399,17'd5032,17'd7520,17'd7030,17'd7346,17'd14590,17'd14591,17'd14592,17'd14180,17'd8491,17'd9253,17'd14739,17'd14740,17'd12320,17'd11723,17'd13059,17'd13691,17'd14593,17'd14594,17'd14741,17'd14595,17'd11330,17'd14063,17'd9795,17'd9795,17'd9795,17'd12777,17'd11725,17'd11054,17'd9666,17'd9666,17'd13938,17'd13938,17'd8026,17'd7691,17'd13692,17'd14596,17'd8325,17'd11193,17'd8181,17'd14438,17'd9120,17'd10256,17'd9956,17'd9120,17'd7524,17'd9800,17'd11597,17'd11196,17'd12324,17'd10530,17'd9670,17'd6416,17'd9123,17'd14178,17'd10911,17'd204,17'd972,17'd206,17'd272,17'd273
},
'{
17'd4733,17'd6584,17'd4887,17'd7711,17'd1688,17'd1127,17'd0,17'd806,17'd21,17'd23,17'd6,17'd5205,17'd8340,17'd8340,17'd8340,17'd8340,17'd8339,17'd8339,17'd8339,17'd8339,17'd8040,17'd8040,17'd5205,17'd5205,17'd6,17'd7,17'd8,17'd4,17'd22,17'd22,17'd23,17'd4,17'd7216,17'd5514,17'd7375,17'd8519,17'd7223,17'd8815,17'd6900,17'd8973,17'd5965,17'd9137,17'd9966,17'd6432,17'd10261,17'd7546,17'd6267,17'd14742,17'd1,17'd2,17'd4247,17'd1831,17'd14743,17'd4244,17'd14744,17'd14745,17'd14746,17'd986,17'd14747,17'd14748,17'd14600,17'd1975,17'd1974,17'd1701,17'd14602,17'd14749,17'd14750,17'd14451,17'd14751,17'd14752,17'd14753,17'd14754,17'd14755,17'd14756,17'd14757,17'd14456,17'd14758,17'd14759,17'd14458,17'd14760,17'd13829,17'd14206,17'd13706,17'd14615,17'd14761,17'd11907,17'd14762,17'd14462,17'd14096,17'd14211,17'd14465,17'd13715,17'd13715,17'd13715,17'd13595,17'd13595,17'd13460,17'd13461,17'd14763,17'd14468,17'd14469,17'd14469,17'd12679,17'd12955,17'd14764,17'd14764,17'd13969,17'd12361,17'd12218,17'd12218,17'd12814,17'd12218,17'd11913,17'd10815,17'd10691,17'd10286,17'd12535,17'd9006,17'd12534,17'd9301,17'd13468,17'd14099,17'd14765,17'd14766,17'd14767,17'd14768,17'd14100,17'd14769,17'd14221,17'd6622,17'd14770,17'd14771,17'd14772,17'd14773,17'd14774,17'd14775,17'd14352,17'd14776,17'd14777,17'd14778,17'd14779,17'd14780,17'd14781,17'd14782,17'd12822,17'd14231,17'd12686,17'd7764,17'd12221,17'd12072,17'd11366,17'd9995,17'd14783,17'd14784,17'd14785,17'd14111,17'd14786,17'd14496,17'd14497,17'd14787,17'd14788,17'd14789,17'd14790,17'd13341,17'd14791,17'd14650,17'd13743,17'd14792,17'd14793,17'd14794,17'd12845,17'd13628,17'd14795,17'd14796,17'd14797,17'd14509,17'd14244,17'd12086,17'd13127,17'd14251,17'd14798,17'd14799,17'd14250,17'd14512,17'd14251,17'd12558,17'd13635,17'd13504,17'd11791,17'd11951,17'd14800,17'd14801,17'd14802,17'd14803,17'd14804,17'd14805,17'd9741,17'd14806,17'd11667,17'd11960,17'd14670,17'd13136,17'd13763,17'd12109,17'd14807,17'd14130,17'd12419,17'd12111,17'd12861,17'd11395,17'd10989,17'd11965,17'd13516,17'd11964,17'd11806,17'd14808,17'd12577,17'd12575,17'd13643,17'd14672,17'd14672,17'd14525,17'd14809,17'd13512,17'd12576,17'd11963,17'd14810,17'd9884,17'd14811,17'd14812,17'd10179,17'd14813,17'd14814,17'd14815,17'd7457,17'd14680,17'd14681,17'd8258,17'd14816,17'd14817,17'd14142,17'd14818,17'd14534,17'd14819,17'd12870,17'd14820,17'd14821,17'd14822,17'd14823,17'd14824,17'd14541,17'd9755,17'd14825,17'd14694,17'd11152,17'd7980,17'd1045,17'd1197,17'd1197,17'd1197,17'd133,17'd133,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd132,17'd132,17'd133,17'd131,17'd2865,17'd14826,17'd14827,17'd14828,17'd14829,17'd14405,17'd14830,17'd14150,17'd14831,17'd14409,17'd14832,17'd14833,17'd13787,17'd13667,17'd14834,17'd14835,17'd14836,17'd14704,17'd14837,17'd14704,17'd14838,17'd14706,17'd14839,17'd8615,17'd12145,17'd14840,17'd12451,17'd8456,17'd12282,17'd12282,17'd8294,17'd13159,17'd13159,17'd8456,17'd9767,17'd11017,17'd8916,17'd14841,17'd14842,17'd9238,17'd13673,17'd7832,17'd9641,17'd14843,17'd14844,17'd14845,17'd14845,17'd14293,17'd14293,17'd14846,17'd14415,17'd14161,17'd14038,17'd9370,17'd11295,17'd11295,17'd14161,17'd14161,17'd14297,17'd14161,17'd14038,17'd10630,17'd14707,17'd9506,17'd13153,17'd14847,17'd13393,17'd13393,17'd14848,17'd14286,17'd14718,17'd14719,17'd9929,17'd9518,17'd10226,17'd12155,17'd12001,17'd12000,17'd12899,17'd12460,17'd12899,17'd12460,17'd12001,17'd12000,17'd13035,17'd14721,17'd14568,17'd13035,17'd13162,17'd12618,17'd12617,17'd13162,17'd14722,17'd14570,17'd14421,17'd14849,17'd13796,17'd14422,17'd14850,17'd14165,17'd13923,17'd14724,17'd14165,17'd13799,17'd13677,17'd13924,17'd13925,17'd13558,17'd13407,17'd14049,17'd12307,17'd12163,17'd14851,17'd14852,17'd14853,17'd14854,17'd7841,17'd14304,17'd13412,17'd13803,17'd14855,17'd14578,17'd14856,17'd14056,17'd14432,17'd14857,17'd14583,17'd14735,17'd14584,17'd14858,17'd4714,17'd12644,17'd197,17'd1813,17'd14859,17'd14859,17'd14860,17'd14861,17'd14862,17'd14863,17'd14864,17'd6872,17'd7684,17'd8018,17'd14592,17'd14180,17'd8491,17'd8795,17'd14865,17'd12319,17'd12320,17'd11723,17'd12489,17'd13937,17'd14594,17'd14594,17'd14741,17'd14741,17'd11330,17'd11330,17'd9795,17'd9795,17'd9795,17'd9795,17'd11725,17'd11054,17'd9541,17'd9541,17'd14437,17'd14437,17'd8026,17'd7691,17'd13692,17'd8325,17'd8325,17'd13692,17'd9955,17'd14438,17'd12490,17'd10256,17'd10256,17'd9956,17'd14866,17'd7034,17'd8655,17'd12493,17'd14439,17'd10655,17'd9958,17'd6727,17'd6889,17'd14178,17'd10911,17'd775,17'd425,17'd269,17'd1407,17'd267
},
'{
17'd4733,17'd4887,17'd4887,17'd7711,17'd1127,17'd2,17'd3,17'd1275,17'd25,17'd5,17'd5205,17'd8190,17'd8340,17'd8340,17'd8340,17'd8340,17'd8339,17'd8339,17'd8339,17'd8040,17'd8040,17'd5205,17'd3753,17'd6,17'd5,17'd5,17'd4,17'd22,17'd22,17'd22,17'd4,17'd5206,17'd5206,17'd5514,17'd5649,17'd8671,17'd8518,17'd8815,17'd13299,17'd9135,17'd8042,17'd9966,17'd8045,17'd6432,17'd10261,17'd7376,17'd14867,17'd15,17'd2,17'd466,17'd1688,17'd2935,17'd4428,17'd4426,17'd7049,17'd14868,17'd986,17'd985,17'd14869,17'd14870,17'd14748,17'd1702,17'd1557,17'd1421,17'd58,17'd14871,17'd14872,17'd14873,17'd14874,17'd14875,17'd14876,17'd5672,17'd14877,17'd14878,17'd14879,17'd14880,17'd14881,17'd14882,17'd14883,17'd14884,17'd11754,17'd13706,17'd14885,17'd11906,17'd14886,17'd14887,17'd14888,17'd14889,17'd14463,17'd14619,17'd14465,17'd13715,17'd13715,17'd13595,17'd13595,17'd13460,17'd14344,17'd14344,17'd14763,17'd14469,17'd14469,17'd13092,17'd12955,17'd14890,17'd14764,17'd14891,17'd12361,17'd12361,17'd13094,17'd13094,17'd12814,17'd11627,17'd11361,17'd10691,17'd13327,17'd9573,17'd9006,17'd10694,17'd9301,17'd12959,17'd14099,17'd14625,17'd14892,17'd14893,17'd14768,17'd14346,17'd14623,17'd14894,17'd14895,17'd14896,17'd14897,17'd14898,17'd14899,17'd14631,17'd14900,17'd14775,17'd14106,17'd13978,17'd14901,17'd14902,17'd14780,17'd14781,17'd14903,17'd14904,17'd13106,17'd12371,17'd12823,17'd9318,17'd10703,17'd14905,17'd10819,17'd10437,17'd14906,17'd14907,17'd14908,17'd14909,17'd14496,17'd14496,17'd14647,17'd14910,17'd14911,17'd14912,17'd13741,17'd14913,17'd13113,17'd13114,17'd13987,17'd11106,17'd14914,17'd12984,17'd11501,17'd14915,17'd14916,17'd14917,17'd14918,17'd14919,17'd12705,17'd12565,17'd14920,17'd14122,17'd14921,17'd14922,17'd12699,17'd14512,17'd14512,17'd13355,17'd14125,17'd14923,17'd13998,17'd14924,17'd14925,17'd14664,17'd14926,17'd11136,17'd14927,17'd9191,17'd14928,17'd14929,17'd11667,17'd13883,17'd12719,17'd12420,17'd12110,17'd13882,17'd14130,17'd14130,17'd12580,17'd13363,17'd13253,17'd14262,17'd11965,17'd10989,17'd11964,17'd13762,17'd11806,17'd14131,17'd12414,17'd12418,17'd14930,17'd14672,17'd14672,17'd14525,17'd13643,17'd12256,17'd12577,17'd11963,17'd14931,17'd9741,17'd8886,17'd8419,17'd14932,17'd14933,17'd14934,17'd14935,17'd14936,17'd14937,17'd12266,17'd14938,17'd14816,17'd12430,17'd14142,17'd14939,17'd12268,17'd14940,17'd14941,17'd14942,17'd14943,17'd14822,17'd14944,17'd14945,17'd10619,17'd12274,17'd14693,17'd9059,17'd11152,17'd7980,17'd1045,17'd3025,17'd3025,17'd1197,17'd133,17'd133,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd132,17'd132,17'd132,17'd131,17'd6369,17'd14946,17'd14947,17'd14948,17'd14949,17'd14950,17'd14406,17'd13909,17'd14951,17'd14284,17'd14952,17'd14718,17'd14953,17'd13395,17'd14834,17'd13668,17'd14954,17'd14704,17'd14955,17'd14413,17'd14704,17'd14956,17'd14957,17'd8457,17'd12145,17'd12895,17'd8294,17'd12282,17'd12282,17'd12282,17'd8294,17'd14958,17'd8456,17'd12138,17'd14560,17'd10884,17'd14558,17'd8293,17'd9088,17'd9238,17'd13665,17'd9505,17'd14959,17'd14960,17'd14961,17'd14962,17'd14963,17'd14964,17'd14293,17'd14846,17'd14038,17'd8610,17'd8611,17'd8611,17'd11831,17'd11831,17'd14038,17'd14161,17'd14297,17'd14297,17'd14161,17'd14161,17'd9640,17'd8761,17'd13153,17'd14965,17'd13270,17'd14848,17'd13393,17'd14565,17'd14966,17'd14967,17'd14720,17'd9387,17'd9518,17'd10226,17'd12155,17'd12000,17'd12154,17'd12460,17'd13036,17'd12899,17'd12154,17'd12000,17'd14721,17'd14721,17'd14569,17'd14568,17'd13035,17'd14721,17'd12618,17'd12617,17'd14421,17'd14570,17'd14570,17'd14723,17'd14164,17'd14422,17'd14968,17'd14969,17'd14724,17'd14724,17'd14724,17'd13923,17'd13924,17'd13677,17'd14970,17'd14971,17'd13406,17'd11575,17'd11854,17'd12468,17'd12163,17'd13408,17'd14972,17'd14726,17'd7330,17'd7505,17'd13681,17'd13285,17'd13564,17'd14728,17'd14973,17'd14974,17'd14580,17'd14975,17'd14976,17'd14735,17'd14584,17'd14858,17'd4714,17'd12644,17'd197,17'd14977,17'd14978,17'd14979,17'd2567,17'd14980,17'd14981,17'd14982,17'd6575,17'd6871,17'd7684,17'd14983,17'd14591,17'd14592,17'd8491,17'd8795,17'd14984,17'd12319,17'd12487,17'd11723,17'd12178,17'd12489,17'd13425,17'd14594,17'd14594,17'd14741,17'd12640,17'd11330,17'd9795,17'd9795,17'd9795,17'd9795,17'd12777,17'd11725,17'd9541,17'd9541,17'd14437,17'd14437,17'd8498,17'd7691,17'd13692,17'd8325,17'd8325,17'd8325,17'd10653,17'd14438,17'd12491,17'd9956,17'd10080,17'd9956,17'd8330,17'd7034,17'd8655,17'd12493,17'd14985,17'd14986,17'd12184,17'd6727,17'd4559,17'd3073,17'd11062,17'd425,17'd206,17'd258,17'd264,17'd457
},
'{
17'd5508,17'd7545,17'd7711,17'd4886,17'd1127,17'd0,17'd283,17'd2591,17'd4,17'd6,17'd5205,17'd8190,17'd8340,17'd8340,17'd8339,17'd8339,17'd8339,17'd8339,17'd8040,17'd8040,17'd8040,17'd3753,17'd3753,17'd6,17'd5,17'd4,17'd23,17'd22,17'd5518,17'd22,17'd4,17'd5206,17'd8,17'd5513,17'd8519,17'd12185,17'd8518,17'd8670,17'd14987,17'd9673,17'd9136,17'd10542,17'd10263,17'd6432,17'd10663,17'd6103,17'd14988,17'd12,17'd13,17'd466,17'd3250,17'd2593,17'd6730,17'd7049,17'd14868,17'd14989,17'd659,17'd35,17'd14869,17'd14869,17'd14990,17'd1971,17'd1700,17'd822,17'd14991,17'd305,17'd1291,17'd2270,17'd14992,17'd14993,17'd13192,17'd14994,17'd14995,17'd14996,17'd14997,17'd14998,17'd14999,17'd15000,17'd15001,17'd15002,17'd13706,17'd12208,17'd12349,17'd14761,17'd15003,17'd14888,17'd15004,17'd15005,17'd13714,17'd14619,17'd14465,17'd14465,17'd12212,17'd13595,17'd13460,17'd12355,17'd14344,17'd14468,17'd14469,17'd14469,17'd14469,17'd13209,17'd12955,17'd14890,17'd14764,17'd14764,17'd12530,17'd12218,17'd11360,17'd12956,17'd11627,17'd11478,17'd11361,17'd10691,17'd12533,17'd9158,17'd9006,17'd15006,17'd12959,17'd13466,17'd15007,17'd14768,17'd15008,17'd14893,17'd14346,17'd15009,17'd15010,17'd15011,17'd15012,17'd15013,17'd15014,17'd15015,17'd15016,17'd15017,17'd15018,17'd14482,17'd14633,17'd14483,17'd15019,17'd15020,17'd15021,17'd15022,17'd15023,17'd8700,17'd14640,17'd7924,17'd10702,17'd9319,17'd15024,17'd10819,17'd13734,17'd15025,17'd15026,17'd15027,17'd15028,17'd15029,17'd15030,17'd15031,17'd15032,17'd14362,17'd14114,17'd13227,17'd13620,17'd15033,17'd15034,17'd13743,17'd15035,17'd11107,17'd11500,17'd13495,17'd15036,17'd15037,17'd15038,17'd15039,17'd13630,17'd13748,17'd13995,17'd12708,17'd13634,17'd15040,17'd15041,17'd15042,17'd14120,17'd14250,17'd14372,17'd13503,17'd11788,17'd15043,17'd15044,17'd15045,17'd15046,17'd15047,17'd15048,17'd15049,17'd15050,17'd12117,17'd15051,17'd15052,17'd13764,17'd15053,17'd11958,17'd12419,17'd14131,17'd15054,17'd15055,17'd14130,17'd12580,17'd12419,17'd12861,17'd14262,17'd11965,17'd10989,17'd11964,17'd13762,17'd11806,17'd12577,17'd12575,17'd12418,17'd14930,17'd14672,17'd14672,17'd14930,17'd12859,17'd12256,17'd12110,17'd11963,17'd10475,17'd9619,17'd9886,17'd15056,17'd14682,17'd15057,17'd15058,17'd15059,17'd14680,17'd15060,17'd14531,17'd7621,17'd13528,17'd15061,17'd14013,17'd15062,17'd15063,17'd15064,17'd15065,17'd10614,17'd15066,17'd15067,17'd14273,17'd15068,17'd15069,17'd7978,17'd9360,17'd9059,17'd14016,17'd8132,17'd3025,17'd3025,17'd3025,17'd1197,17'd133,17'd133,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd133,17'd132,17'd12127,17'd4655,17'd15070,17'd15071,17'd15072,17'd15073,17'd15074,17'd15075,17'd15076,17'd15077,17'd15078,17'd14967,17'd14953,17'd13271,17'd15079,17'd14835,17'd14555,17'd14704,17'd14955,17'd14837,17'd14704,17'd15080,17'd15081,17'd11994,17'd11994,17'd12896,17'd8294,17'd12282,17'd12282,17'd12282,17'd8456,17'd14958,17'd8614,17'd11987,17'd14038,17'd10630,17'd14707,17'd8293,17'd9088,17'd14420,17'd13672,17'd14708,17'd15082,17'd15083,17'd15084,17'd15084,17'd15085,17'd14961,17'd14844,17'd14709,17'd10630,17'd8611,17'd8759,17'd9372,17'd11831,17'd14038,17'd14158,17'd14415,17'd15086,17'd14296,17'd15086,17'd15086,17'd14161,17'd10630,17'd9222,17'd15087,17'd12743,17'd13154,17'd13270,17'd14965,17'd15088,17'd14966,17'd15089,17'd15090,17'd14044,17'd9385,17'd10227,17'd12155,17'd12155,17'd15091,17'd15092,17'd13163,17'd12899,17'd12295,17'd12618,17'd13162,17'd14569,17'd14569,17'd14569,17'd14568,17'd14721,17'd12618,17'd14571,17'd14722,17'd15093,17'd14571,17'd14723,17'd14849,17'd14850,17'd14968,17'd14850,17'd14724,17'd14969,17'd14724,17'd14970,17'd13925,17'd14970,17'd15094,17'd13925,17'd14166,17'd14049,17'd12161,17'd14167,17'd13408,17'd15095,17'd15096,17'd7671,17'd7841,17'd13411,17'd13412,17'd15097,17'd13803,17'd15098,17'd15099,17'd15100,17'd15101,17'd15102,17'd15103,17'd15104,17'd6890,17'd5183,17'd12644,17'd776,17'd417,17'd2102,17'd2398,17'd2567,17'd15105,17'd14861,17'd15106,17'd5635,17'd7028,17'd7516,17'd7684,17'd7854,17'd7855,17'd8170,17'd8491,17'd14984,17'd11722,17'd12487,17'd15107,17'd12178,17'd12489,17'd13425,17'd13425,17'd14594,17'd14594,17'd12918,17'd12640,17'd11330,17'd14063,17'd9795,17'd9795,17'd14064,17'd14064,17'd9666,17'd9666,17'd8651,17'd15108,17'd8651,17'd8026,17'd13692,17'd8325,17'd8325,17'd14596,17'd12641,17'd7698,17'd7531,17'd9120,17'd10080,17'd10256,17'd7034,17'd8330,17'd12182,17'd15109,17'd15110,17'd15111,17'd15112,17'd10258,17'd4559,17'd2097,17'd6407,17'd1666,17'd261,17'd262,17'd1274,17'd15113
},
'{
17'd5508,17'd7545,17'd4886,17'd6419,17'd2,17'd3,17'd1275,17'd2591,17'd8,17'd6,17'd5205,17'd8190,17'd8340,17'd8340,17'd8339,17'd8339,17'd8339,17'd8040,17'd8040,17'd5793,17'd3753,17'd3753,17'd6,17'd5,17'd8,17'd4,17'd23,17'd22,17'd5518,17'd22,17'd4,17'd8,17'd5206,17'd13062,17'd15114,17'd15115,17'd8973,17'd13182,17'd15116,17'd8347,17'd7892,17'd10542,17'd6271,17'd6271,17'd6595,17'd14187,17'd3,17'd806,17'd12,17'd14,17'd2592,17'd4738,17'd15117,17'd14745,17'd14868,17'd15118,17'd36,17'd35,17'd15119,17'd15120,17'd15121,17'd1836,17'd1699,17'd665,17'd15122,17'd68,17'd2269,17'd2128,17'd14875,17'd14876,17'd5395,17'd15123,17'd15124,17'd15125,17'd15126,17'd15127,17'd14882,17'd15128,17'd15129,17'd15130,17'd13706,17'd15131,17'd12209,17'd15132,17'd15133,17'd15134,17'd15135,17'd15136,17'd14619,17'd14619,17'd14465,17'd14619,17'd12212,17'd13596,17'd13461,17'd13461,17'd14468,17'd14469,17'd14469,17'd13092,17'd13209,17'd13210,17'd14890,17'd15137,17'd14764,17'd12218,17'd12218,17'd12218,17'd12956,17'd12956,17'd11627,17'd11361,17'd10691,17'd10286,17'd9158,17'd9574,17'd10694,17'd15138,17'd13466,17'd14100,17'd14765,17'd14767,17'd15008,17'd14892,17'd15009,17'd15139,17'd15011,17'd15140,17'd15141,17'd15142,17'd15143,17'd15144,17'd15017,17'd15145,17'd13976,17'd15146,17'd14633,17'd14483,17'd15147,17'd15148,17'd15149,17'd15150,17'd9016,17'd15151,17'd15152,17'd9021,17'd9591,17'd14360,17'd15024,17'd13734,17'd13857,17'd15153,17'd14785,17'd15154,17'd15155,17'd15156,17'd15157,17'd15031,17'd15158,17'd15159,17'd13111,17'd15160,17'd14913,17'd15161,17'd15162,17'd12385,17'd15163,17'd15164,17'd12982,17'd11111,17'd15165,17'd15166,17'd15167,17'd13872,17'd15168,17'd15169,17'd14662,17'd13246,17'd14122,17'd15170,17'd15171,17'd13874,17'd12699,17'd14371,17'd14124,17'd15172,17'd11948,17'd15173,17'd12250,17'd15174,17'd15175,17'd15176,17'd15177,17'd15178,17'd15179,17'd15180,17'd15181,17'd15182,17'd11806,17'd12719,17'd12420,17'd13882,17'd15183,17'd15054,17'd15055,17'd15184,17'd12109,17'd12420,17'd11962,17'd14262,17'd11965,17'd10989,17'd11964,17'd15185,17'd11960,17'd12414,17'd12418,17'd12418,17'd14672,17'd14524,17'd14930,17'd14930,17'd12859,17'd12575,17'd12111,17'd15186,17'd10473,17'd15187,17'd10178,17'd15188,17'd15189,17'd15190,17'd15191,17'd14680,17'd15192,17'd15193,17'd10747,17'd15194,17'd13528,17'd15061,17'd14013,17'd15195,17'd15196,17'd15197,17'd15198,17'd11146,17'd15199,17'd15200,17'd13382,17'd15201,17'd12435,17'd9756,17'd8131,17'd9059,17'd14016,17'd11289,17'd3025,17'd3025,17'd3025,17'd1197,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd15202,17'd5470,17'd15203,17'd15204,17'd15205,17'd15206,17'd15207,17'd15208,17'd13910,17'd14026,17'd14952,17'd14719,17'd14411,17'd15209,17'd13272,17'd13668,17'd14954,17'd14704,17'd14837,17'd14837,17'd14287,17'd15080,17'd14033,17'd9649,17'd11994,17'd12896,17'd12283,17'd12282,17'd12282,17'd8456,17'd13159,17'd8614,17'd12138,17'd9767,17'd10630,17'd15210,17'd13672,17'd7994,17'd14036,17'd8148,17'd11693,17'd14844,17'd15211,17'd15212,17'd15213,17'd15213,17'd15085,17'd14961,17'd15214,17'd14708,17'd9640,17'd8611,17'd7993,17'd8759,17'd11295,17'd14161,17'd14415,17'd15086,17'd14296,17'd14296,17'd14296,17'd14296,17'd14161,17'd10630,17'd15215,17'd9222,17'd12886,17'd15216,17'd15217,17'd15217,17'd14965,17'd15088,17'd15218,17'd15090,17'd15219,17'd15220,17'd10773,17'd10227,17'd11309,17'd12757,17'd13163,17'd13163,17'd15221,17'd12899,17'd12618,17'd13162,17'd14721,17'd14568,17'd15222,17'd15222,17'd14568,17'd14721,17'd14421,17'd14421,17'd14570,17'd14570,17'd14571,17'd15223,17'd14850,17'd15224,17'd15225,17'd14969,17'd14850,17'd14969,17'd15094,17'd14970,17'd14970,17'd15094,17'd14970,17'd13278,17'd11854,17'd12760,17'd12161,17'd14167,17'd15226,17'd15227,17'd15228,17'd7330,17'd13680,17'd13284,17'd13412,17'd13564,17'd14054,17'd14055,17'd15229,17'd15230,17'd15231,17'd15232,17'd15104,17'd6890,17'd5183,17'd15233,17'd776,17'd943,17'd15234,17'd2397,17'd2566,17'd15235,17'd14980,17'd15236,17'd4065,17'd5365,17'd7343,17'd7684,17'd7514,17'd7855,17'd8170,17'd8491,17'd15237,17'd10076,17'd10077,17'd12487,17'd11723,17'd12489,17'd13425,17'd13425,17'd14594,17'd14594,17'd15238,17'd12918,17'd12640,17'd11330,17'd9795,17'd9795,17'd14063,17'd14064,17'd11054,17'd9666,17'd8651,17'd15108,17'd8651,17'd8498,17'd8325,17'd8325,17'd8325,17'd14596,17'd13692,17'd9955,17'd7531,17'd12490,17'd10256,17'd10256,17'd9800,17'd8330,17'd12182,17'd11332,17'd12493,17'd14314,17'd10530,17'd9670,17'd4559,17'd1946,17'd6407,17'd1956,17'd15239,17'd2115,17'd15240,17'd15240
},
'{
17'd7214,17'd7214,17'd1127,17'd14,17'd0,17'd3,17'd25,17'd4,17'd7,17'd7,17'd5205,17'd8040,17'd8040,17'd8040,17'd8340,17'd8340,17'd8340,17'd8040,17'd5793,17'd3753,17'd3753,17'd3753,17'd5,17'd5,17'd8,17'd4,17'd23,17'd22,17'd5518,17'd22,17'd23,17'd4,17'd7216,17'd12925,17'd9135,17'd6732,17'd8825,17'd6427,17'd9673,17'd7724,17'd8824,17'd9420,17'd6271,17'd9272,17'd6596,17'd15241,17'd8814,17'd8814,17'd15242,17'd6419,17'd2934,17'd6730,17'd14746,17'd15243,17'd14599,17'd15244,17'd35,17'd35,17'd2261,17'd1694,17'd15245,17'd15246,17'd15247,17'd53,17'd15248,17'd1291,17'd2270,17'd14752,17'd13442,17'd15249,17'd15250,17'd15251,17'd15252,17'd15253,17'd15254,17'd15255,17'd15000,17'd13705,17'd15130,17'd13591,17'd14614,17'd15256,17'd12521,17'd15257,17'd15258,17'd15259,17'd13596,17'd13595,17'd12212,17'd13715,17'd14619,17'd14619,17'd13596,17'd13716,17'd13461,17'd12357,17'd14469,17'd14469,17'd14469,17'd13092,17'd13209,17'd13210,17'd15137,17'd14764,17'd12530,17'd12218,17'd13094,17'd12956,17'd11627,17'd11627,17'd12066,17'd12066,17'd10691,17'd10286,17'd11232,17'd10428,17'd10113,17'd13601,17'd14345,17'd14473,17'd14767,17'd14893,17'd14892,17'd15260,17'd15261,17'd15262,17'd15140,17'd15263,17'd15264,17'd15265,17'd15266,17'd15267,17'd15268,17'd15269,17'd13977,17'd14633,17'd14106,17'd15270,17'd15271,17'd15272,17'd14903,17'd9017,17'd15273,17'd15274,17'd7764,17'd9591,17'd14360,17'd11096,17'd15275,17'd10437,17'd15153,17'd15276,17'd15277,17'd15278,17'd15279,17'd15280,17'd15281,17'd14497,17'd15158,17'd15159,17'd14363,17'd13112,17'd13228,17'd11491,17'd15282,17'd15283,17'd15284,17'd15285,17'd15286,17'd15165,17'd15287,17'd15288,17'd15289,17'd15290,17'd12564,17'd14124,17'd15291,17'd13634,17'd14251,17'd14250,17'd15292,17'd15292,17'd13127,17'd14253,17'd13753,17'd11789,17'd15293,17'd14925,17'd15294,17'd14669,17'd14134,17'd15295,17'd15296,17'd12264,17'd15297,17'd15298,17'd10477,17'd15175,17'd12581,17'd12106,17'd12580,17'd13882,17'd15054,17'd15299,17'd13761,17'd14131,17'd12580,17'd11958,17'd11963,17'd11395,17'd14262,17'd14262,17'd13762,17'd13520,17'd13761,17'd12414,17'd12418,17'd12416,17'd14672,17'd14524,17'd14930,17'd14930,17'd12997,17'd12575,17'd12113,17'd10737,17'd15300,17'd8720,17'd15301,17'd15302,17'd8891,17'd11141,17'd15303,17'd14932,17'd10995,17'd10180,17'd10747,17'd15304,17'd15305,17'd15306,17'd15307,17'd15308,17'd15309,17'd12731,17'd15310,17'd12872,17'd15311,17'd15312,17'd15313,17'd10619,17'd10621,17'd7812,17'd8131,17'd9059,17'd14276,17'd8132,17'd3025,17'd1197,17'd1197,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd133,17'd132,17'd357,17'd3028,17'd15314,17'd15315,17'd15316,17'd14698,17'd15317,17'd14700,17'd15076,17'd14701,17'd14409,17'd15089,17'd14953,17'd13154,17'd13155,17'd14553,17'd13789,17'd15318,17'd15319,17'd15319,17'd15320,17'd15321,17'd14837,17'd9776,17'd11994,17'd8615,17'd15322,17'd12282,17'd12282,17'd8294,17'd14958,17'd8456,17'd9506,17'd15215,17'd15210,17'd9506,17'd7832,17'd7994,17'd8149,17'd8762,17'd15323,17'd14961,17'd15212,17'd15324,17'd15325,17'd15213,17'd15085,17'd15326,17'd14843,17'd9640,17'd8611,17'd10501,17'd8454,17'd8454,17'd11295,17'd14161,17'd14161,17'd14297,17'd14713,17'd15327,17'd15327,17'd14564,17'd14713,17'd15328,17'd14158,17'd15329,17'd15330,17'd12605,17'd12743,17'd15331,17'd13023,17'd13270,17'd14966,17'd15089,17'd15332,17'd15333,17'd10773,17'd15334,17'd10894,17'd15335,17'd12757,17'd13163,17'd15221,17'd15221,17'd14568,17'd14721,17'd12618,17'd13035,17'd15222,17'd15222,17'd14569,17'd14568,17'd15336,17'd15337,17'd14722,17'd15093,17'd14722,17'd15338,17'd15223,17'd15339,17'd15339,17'd14723,17'd14850,17'd14850,17'd15340,17'd14971,17'd14970,17'd14971,17'd14971,17'd13925,17'd13407,17'd14049,17'd12307,17'd15341,17'd14425,17'd15342,17'd15343,17'd15344,17'd13680,17'd13411,17'd13681,17'd15097,17'd13803,17'd15098,17'd15345,17'd15346,17'd15347,17'd15348,17'd14858,17'd8187,17'd5631,17'd12644,17'd776,17'd196,17'd14977,17'd2397,17'd2400,17'd2566,17'd15105,17'd15349,17'd3717,17'd15350,17'd6870,17'd7345,17'd7514,17'd7854,17'd8170,17'd8491,17'd11191,17'd14984,17'd11722,17'd11593,17'd15107,17'd15351,17'd13937,17'd13937,17'd14594,17'd14741,17'd15352,17'd15238,17'd12640,17'd11330,17'd11330,17'd14063,17'd14063,17'd14064,17'd12777,17'd11054,17'd8651,17'd15108,17'd15108,17'd8651,17'd8325,17'd13692,17'd8325,17'd8325,17'd8325,17'd10653,17'd12491,17'd12491,17'd9120,17'd9956,17'd9956,17'd12322,17'd12492,17'd12182,17'd11879,17'd14439,17'd10655,17'd12494,17'd4401,17'd6415,17'd6407,17'd260,17'd15353,17'd1123,17'd15354,17'd15355
},
'{
17'd7214,17'd13436,17'd1127,17'd0,17'd3,17'd1275,17'd4,17'd4,17'd7,17'd5205,17'd8040,17'd8040,17'd8040,17'd8040,17'd8340,17'd8340,17'd8340,17'd8040,17'd3753,17'd3753,17'd3753,17'd6,17'd5,17'd5,17'd23,17'd22,17'd22,17'd5518,17'd5518,17'd22,17'd4,17'd8,17'd7375,17'd12782,17'd8661,17'd6435,17'd13299,17'd15116,17'd6588,17'd7058,17'd8824,17'd9272,17'd6271,17'd9137,17'd13941,17'd2591,17'd2933,17'd8814,17'd15356,17'd15357,17'd15358,17'd15359,17'd15360,17'd15361,17'd15362,17'd473,17'd35,17'd471,17'd2428,17'd15363,17'd15246,17'd15364,17'd988,17'd15365,17'd15366,17'd487,17'd15367,17'd15368,17'd15369,17'd15370,17'd5071,17'd15371,17'd15372,17'd15373,17'd15374,17'd15375,17'd15376,17'd13450,17'd13591,17'd14336,17'd14615,17'd15377,17'd15378,17'd15379,17'd15380,17'd13716,17'd13326,17'd15381,17'd13459,17'd13595,17'd14619,17'd15382,17'd13838,17'd12356,17'd12357,17'd14469,17'd14469,17'd13092,17'd13092,17'd13599,17'd13210,17'd15383,17'd14764,17'd14764,17'd12530,17'd12218,17'd11360,17'd12956,17'd11627,17'd11361,17'd12066,17'd10562,17'd13327,17'd11232,17'd10693,17'd15138,17'd13470,17'd13843,17'd14473,17'd15384,17'd15385,17'd14893,17'd15386,17'd15387,17'd15139,17'd15262,17'd15140,17'd15388,17'd15389,17'd15390,17'd15266,17'd15391,17'd15392,17'd15393,17'd15394,17'd15395,17'd15396,17'd15397,17'd15398,17'd15399,17'd15400,17'd13733,17'd15401,17'd15402,17'd9318,17'd14360,17'd15403,17'd10436,17'd15404,17'd15405,17'd15406,17'd15407,17'd15408,17'd15409,17'd15410,17'd15280,17'd15281,17'd15411,17'd15158,17'd15159,17'd13340,17'd12832,17'd13113,17'd11492,17'd15412,17'd15413,17'd15414,17'd15415,17'd15416,17'd15417,17'd15418,17'd15419,17'd12983,17'd15420,17'd13503,17'd13356,17'd15421,17'd15040,17'd14250,17'd12558,17'd15422,17'd15422,17'd14253,17'd15423,17'd11940,17'd15424,17'd15425,17'd12112,17'd15426,17'd15427,17'd9620,17'd15428,17'd9744,17'd15429,17'd15430,17'd15431,17'd15432,17'd13135,17'd13252,17'd15433,17'd12579,17'd15184,17'd15054,17'd13366,17'd13761,17'd12577,17'd12995,17'd12719,17'd13362,17'd11395,17'd11395,17'd11964,17'd13762,17'd11806,17'd12110,17'd15434,17'd12416,17'd12416,17'd14672,17'd14524,17'd14930,17'd14930,17'd12997,17'd12577,17'd12861,17'd10739,17'd9473,17'd11530,17'd15435,17'd15436,17'd15437,17'd15438,17'd15439,17'd15440,17'd15441,17'd9890,17'd15442,17'd14266,17'd15443,17'd13259,17'd15444,17'd15445,17'd15446,17'd15447,17'd12124,17'd12125,17'd14689,17'd15448,17'd12434,17'd13533,17'd11977,17'd13776,17'd8131,17'd14276,17'd14276,17'd11413,17'd1197,17'd133,17'd133,17'd133,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd357,17'd4816,17'd15449,17'd15450,17'd15451,17'd15452,17'd15453,17'd14700,17'd15454,17'd15455,17'd15456,17'd15457,17'd15458,17'd15459,17'd15460,17'd14553,17'd13789,17'd15318,17'd14032,17'd14032,17'd15320,17'd15319,17'd15461,17'd15462,17'd11994,17'd8615,17'd15322,17'd12282,17'd8456,17'd8294,17'd14958,17'd8294,17'd9506,17'd15215,17'd15463,17'd14841,17'd7832,17'd13159,17'd8457,17'd11162,17'd14961,17'd15212,17'd15464,17'd15465,17'd15466,17'd15212,17'd14961,17'd15214,17'd14708,17'd9640,17'd10629,17'd8610,17'd8610,17'd11831,17'd14038,17'd14038,17'd14038,17'd14161,17'd15328,17'd14713,17'd14713,17'd15327,17'd14564,17'd14713,17'd14415,17'd14158,17'd15330,17'd15467,17'd15216,17'd15216,17'd15331,17'd15468,17'd15469,17'd14833,17'd14719,17'd15470,17'd15471,17'd15472,17'd11175,17'd10894,17'd12296,17'd13163,17'd13036,17'd15473,17'd15474,17'd14721,17'd12900,17'd13035,17'd14569,17'd14569,17'd14569,17'd15222,17'd15475,17'd15336,17'd14722,17'd15093,17'd14570,17'd15339,17'd14723,17'd15338,17'd14571,17'd15339,17'd14850,17'd14968,17'd15476,17'd15094,17'd14970,17'd14970,17'd14971,17'd15094,17'd13406,17'd14166,17'd12760,17'd14050,17'd15477,17'd15478,17'd15479,17'd14575,17'd7505,17'd13411,17'd13680,17'd13681,17'd13564,17'd14578,17'd15480,17'd15481,17'd15482,17'd15483,17'd15484,17'd4714,17'd14586,17'd12644,17'd941,17'd1671,17'd943,17'd2241,17'd2246,17'd2400,17'd14860,17'd15485,17'd15486,17'd15487,17'd6869,17'd7345,17'd7514,17'd7854,17'd8170,17'd8491,17'd11191,17'd11050,17'd10076,17'd10077,17'd12487,17'd15488,17'd13424,17'd13937,17'd13425,17'd14741,17'd15352,17'd15238,17'd12776,17'd11330,17'd11330,17'd11330,17'd14063,17'd14063,17'd9795,17'd11054,17'd8651,17'd8651,17'd15489,17'd15108,17'd14596,17'd13692,17'd8325,17'd8325,17'd8325,17'd11195,17'd12491,17'd7531,17'd12322,17'd9956,17'd9956,17'd12322,17'd12492,17'd12182,17'd15490,17'd15490,17'd10793,17'd9413,17'd15491,17'd1946,17'd7210,17'd427,17'd15353,17'd405,17'd15492,17'd770
},
'{
17'd2594,17'd1127,17'd0,17'd12,17'd2423,17'd2933,17'd4,17'd7374,17'd8190,17'd5205,17'd8040,17'd8040,17'd8340,17'd8340,17'd8340,17'd8040,17'd3594,17'd3594,17'd3753,17'd3753,17'd6,17'd5,17'd24,17'd23,17'd23,17'd5518,17'd5518,17'd5518,17'd22,17'd22,17'd8,17'd5514,17'd5649,17'd13297,17'd8661,17'd13431,17'd15493,17'd9673,17'd8825,17'd7892,17'd6105,17'd10542,17'd9682,17'd6428,17'd807,17'd15494,17'd8814,17'd465,17'd15495,17'd7372,17'd15496,17'd14744,17'd15360,17'd15497,17'd986,17'd295,17'd294,17'd471,17'd2428,17'd660,17'd1698,17'd15498,17'd301,17'd15248,17'd1291,17'd2270,17'd15499,17'd14753,17'd15500,17'd15501,17'd15502,17'd15503,17'd15504,17'd15505,17'd15506,17'd15507,17'd15508,17'd15509,17'd15510,17'd15131,17'd15511,17'd15512,17'd15513,17'd15514,17'd15515,17'd13460,17'd13326,17'd13325,17'd13595,17'd13595,17'd14619,17'd15136,17'd13716,17'd13597,17'd14469,17'd12527,17'd12527,17'd12527,17'd15516,17'd13093,17'd14890,17'd14764,17'd14764,17'd14622,17'd12218,17'd13094,17'd12956,17'd11627,17'd12066,17'd11914,17'd11914,17'd10427,17'd10692,17'd9574,17'd15517,17'd13470,17'd15518,17'd14345,17'd14474,17'd15519,17'd14892,17'd15520,17'd15521,17'd15522,17'd15523,17'd15524,17'd15011,17'd15525,17'd15526,17'd15527,17'd15528,17'd15529,17'd15269,17'd15530,17'd15531,17'd15532,17'd15533,17'd15534,17'd15535,17'd15536,17'd13106,17'd12685,17'd15537,17'd15538,17'd9853,17'd10703,17'd10436,17'd15539,17'd15540,17'd15541,17'd15542,17'd15543,17'd15279,17'd15410,17'd15280,17'd15544,17'd15545,17'd15546,17'd15158,17'd14237,17'd13340,17'd15547,17'd11637,17'd15548,17'd15549,17'd15550,17'd13991,17'd15286,17'd15551,17'd15552,17'd14797,17'd15553,17'd15554,17'd13130,17'd15555,17'd15556,17'd15557,17'd15558,17'd12558,17'd15559,17'd15560,17'd13130,17'd14125,17'd14923,17'd15561,17'd15562,17'd15563,17'd15564,17'd15565,17'd15566,17'd15567,17'd15568,17'd15429,17'd8569,17'd15569,17'd14666,17'd11666,17'd11958,17'd15570,17'd12417,17'd12579,17'd12109,17'd13761,17'd13761,17'd12718,17'd12252,17'd13365,17'd14002,17'd11963,17'd11395,17'd13516,17'd11964,17'd11963,17'd11961,17'd12110,17'd12109,17'd12859,17'd14930,17'd15571,17'd15571,17'd14672,17'd14672,17'd12859,17'd12419,17'd14262,17'd10477,17'd9342,17'd15568,17'd12726,17'd15572,17'd15573,17'd12429,17'd14681,17'd10995,17'd10746,17'd10029,17'd15194,17'd15574,17'd15575,17'd13259,17'd14939,17'd15576,17'd15577,17'd15578,17'd10867,17'd12433,17'd15067,17'd13657,17'd15069,17'd9495,17'd8597,17'd14275,17'd14275,17'd14016,17'd11289,17'd11413,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd135,17'd131,17'd15579,17'd4500,17'd6058,17'd15580,17'd15581,17'd15582,17'd15583,17'd15584,17'd14408,17'd14549,17'd15585,17'd14966,17'd14965,17'd15586,17'd14835,17'd13548,17'd14838,17'd14704,17'd15587,17'd15588,17'd14032,17'd15589,17'd15590,17'd12611,17'd8295,17'd12282,17'd12283,17'd8456,17'd13159,17'd8456,17'd8456,17'd8761,17'd15215,17'd14707,17'd13672,17'd7998,17'd12451,17'd11988,17'd15591,17'd15212,17'd15324,17'd15465,17'd15466,17'd15592,17'd15593,17'd14159,17'd15594,17'd9370,17'd10047,17'd9640,17'd9370,17'd14415,17'd14415,17'd14038,17'd14161,17'd15594,17'd15594,17'd15594,17'd15594,17'd14713,17'd15327,17'd15327,17'd14713,17'd15328,17'd14709,17'd10884,17'd11017,17'd15595,17'd12605,17'd15596,17'd15331,17'd15217,17'd15597,17'd14718,17'd15598,17'd15599,17'd15600,17'd15601,17'd10894,17'd12155,17'd12756,17'd13036,17'd15222,17'd15474,17'd15602,17'd13035,17'd13162,17'd14721,17'd15222,17'd15473,17'd15474,17'd15603,17'd15604,17'd14722,17'd14570,17'd15605,17'd15093,17'd14421,17'd15338,17'd15339,17'd14722,17'd15606,17'd15606,17'd15607,17'd15608,17'd15609,17'd15610,17'd13923,17'd13923,17'd14970,17'd14166,17'd11853,17'd12307,17'd15611,17'd15612,17'd15479,17'd15096,17'd14427,17'd15613,17'd13680,17'd15614,17'd13564,17'd14578,17'd15615,17'd15616,17'd15617,17'd15618,17'd14858,17'd4714,17'd15233,17'd941,17'd415,17'd196,17'd15619,17'd1948,17'd2104,17'd2400,17'd15620,17'd15621,17'd15622,17'd6408,17'd5502,17'd6870,17'd7684,17'd14983,17'd8018,17'd8491,17'd11191,17'd11191,17'd10076,17'd11722,17'd12320,17'd15488,17'd12489,17'd13937,17'd13425,17'd13691,17'd15623,17'd15352,17'd15238,17'd12640,17'd11330,17'd11330,17'd11330,17'd14064,17'd14063,17'd14181,17'd8651,17'd8651,17'd15108,17'd15489,17'd15624,17'd8325,17'd8325,17'd8325,17'd8325,17'd11193,17'd9956,17'd7531,17'd12922,17'd12182,17'd11332,17'd11332,17'd12182,17'd12642,17'd15490,17'd11879,17'd10793,17'd8332,17'd3875,17'd7041,17'd3742,17'd7512,17'd15625,17'd15626,17'd1542,17'd15627
},
'{
17'd4247,17'd466,17'd12,17'd3,17'd806,17'd2933,17'd8,17'd7374,17'd5205,17'd5205,17'd8040,17'd8040,17'd8040,17'd8040,17'd8040,17'd5205,17'd3753,17'd3753,17'd3753,17'd5,17'd5,17'd24,17'd4,17'd4,17'd23,17'd5518,17'd5518,17'd22,17'd22,17'd4,17'd5378,17'd5513,17'd12649,17'd13181,17'd13431,17'd14987,17'd15628,17'd15116,17'd8973,17'd7380,17'd9272,17'd9420,17'd6434,17'd5797,17'd7725,17'd7215,17'd8814,17'd13,17'd15357,17'd13428,17'd15496,17'd15629,17'd14599,17'd15362,17'd814,17'd36,17'd471,17'd811,17'd1553,17'd474,17'd15364,17'd15630,17'd15365,17'd15366,17'd15631,17'd13954,17'd14875,17'd2959,17'd4106,17'd4594,17'd15632,17'd15633,17'd15634,17'd15127,17'd15635,17'd15636,17'd15508,17'd13316,17'd15510,17'd14885,17'd15637,17'd15638,17'd15379,17'd15639,17'd13716,17'd13326,17'd12952,17'd13325,17'd13595,17'd13596,17'd15136,17'd13838,17'd12356,17'd12357,17'd12527,17'd12527,17'd12527,17'd12527,17'd12813,17'd13211,17'd14764,17'd14891,17'd14622,17'd14470,17'd12218,17'd12218,17'd12956,17'd15640,17'd12066,17'd12066,17'd10691,17'd10817,17'd9574,17'd10429,17'd13469,17'd13843,17'd14345,17'd14473,17'd15641,17'd15384,17'd15520,17'd15642,17'd15643,17'd15644,17'd15645,17'd15645,17'd15646,17'd15647,17'd15527,17'd15648,17'd15528,17'd15649,17'd15650,17'd15651,17'd15652,17'd15653,17'd15654,17'd15398,17'd15655,17'd15656,17'd14640,17'd7265,17'd15402,17'd15657,17'd9451,17'd15275,17'd15539,17'd15658,17'd15541,17'd15659,17'd15660,17'd15278,17'd15410,17'd15661,17'd15280,17'd15281,17'd15411,17'd15662,17'd15663,17'd13985,17'd15160,17'd15664,17'd12382,17'd15665,17'd15666,17'd15667,17'd10714,17'd15668,17'd15552,17'd15669,17'd13992,17'd15670,17'd15560,17'd15671,17'd13637,17'd15672,17'd15673,17'd14371,17'd12705,17'd15674,17'd15675,17'd15676,17'd12710,17'd11949,17'd15677,17'd15678,17'd15679,17'd15680,17'd15681,17'd15682,17'd15683,17'd14675,17'd8725,17'd15684,17'd14928,17'd14810,17'd13135,17'd15685,17'd15570,17'd13515,17'd12579,17'd12579,17'd14130,17'd13761,17'd12718,17'd15686,17'd13365,17'd14002,17'd11963,17'd11395,17'd11964,17'd13762,17'd13135,17'd13761,17'd12414,17'd12418,17'd14930,17'd14930,17'd15687,17'd15571,17'd14930,17'd12859,17'd12575,17'd12857,17'd12720,17'd15688,17'd8873,17'd12867,17'd15689,17'd15690,17'd12591,17'd15691,17'd15692,17'd15693,17'd15694,17'd12727,17'd14392,17'd15575,17'd12267,17'd15695,17'd15696,17'd15697,17'd15698,17'd15699,17'd11818,17'd10615,17'd15700,17'd15313,17'd15701,17'd15702,17'd14693,17'd14016,17'd14016,17'd11152,17'd11413,17'd1045,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd131,17'd6691,17'd15703,17'd13384,17'd15704,17'd15705,17'd15706,17'd15707,17'd15708,17'd15455,17'd15456,17'd15332,17'd15709,17'd15710,17'd12888,17'd14553,17'd13548,17'd14838,17'd14033,17'd15711,17'd15320,17'd14032,17'd15589,17'd15712,17'd8296,17'd8615,17'd12282,17'd8456,17'd13159,17'd13159,17'd8614,17'd12138,17'd8761,17'd8761,17'd13672,17'd7994,17'd7998,17'd12611,17'd11298,17'd15713,17'd15714,17'd15715,17'd15466,17'd15716,17'd15717,17'd15718,17'd15086,17'd14161,17'd9370,17'd10363,17'd9370,17'd15594,17'd15328,17'd15328,17'd14161,17'd14161,17'd15594,17'd15594,17'd15594,17'd15594,17'd14713,17'd15327,17'd15327,17'd15327,17'd15328,17'd15328,17'd14709,17'd10884,17'd10631,17'd15595,17'd15719,17'd15468,17'd15217,17'd14953,17'd15709,17'd15090,17'd15720,17'd15600,17'd15721,17'd15721,17'd15335,17'd12756,17'd12899,17'd15222,17'd15722,17'd15602,17'd14569,17'd13035,17'd13035,17'd14569,17'd15474,17'd15474,17'd15723,17'd15723,17'd15724,17'd15605,17'd15605,17'd15093,17'd14722,17'd15339,17'd15339,17'd14571,17'd15725,17'd15607,17'd15607,17'd15726,17'd15727,17'd15610,17'd13923,17'd13923,17'd14971,17'd13278,17'd11854,17'd11854,17'd15728,17'd15611,17'd15612,17'd15729,17'd15730,17'd13680,17'd13680,17'd15614,17'd13564,17'd14578,17'd15731,17'd15732,17'd15733,17'd15734,17'd15735,17'd4714,17'd15233,17'd776,17'd415,17'd415,17'd196,17'd1947,17'd2103,17'd2246,17'd15736,17'd15737,17'd15738,17'd6241,17'd5366,17'd6870,17'd7684,17'd14983,17'd8018,17'd8491,17'd11191,17'd11444,17'd9405,17'd12018,17'd12019,17'd12320,17'd13423,17'd12489,17'd13425,17'd13425,17'd15623,17'd15623,17'd15238,17'd12776,17'd12640,17'd11330,17'd11330,17'd14063,17'd14064,17'd14181,17'd15108,17'd15108,17'd15108,17'd15108,17'd15624,17'd14596,17'd14596,17'd8325,17'd13692,17'd11193,17'd9956,17'd12491,17'd12922,17'd12182,17'd12182,17'd11332,17'd12492,17'd12642,17'd15490,17'd12493,17'd15739,17'd8331,17'd8952,17'd3875,17'd4422,17'd208,17'd15740,17'd15741,17'd399,17'd15742
},
'{
17'd2595,17'd466,17'd12,17'd806,17'd21,17'd23,17'd6,17'd7,17'd5205,17'd3753,17'd3753,17'd5205,17'd5205,17'd5205,17'd3753,17'd3753,17'd3753,17'd6,17'd6,17'd5,17'd24,17'd23,17'd4,17'd8,17'd22,17'd5518,17'd20,17'd21,17'd25,17'd5647,17'd8510,17'd13574,17'd6427,17'd8347,17'd15743,17'd15744,17'd10659,17'd6427,17'd13183,17'd8815,17'd9966,17'd8511,17'd5796,17'd6425,17'd978,17'd2421,17'd1128,17'd15745,17'd7214,17'd15746,17'd15496,17'd15118,17'd1279,17'd814,17'd985,17'd36,17'd811,17'd811,17'd37,17'd1836,17'd1133,17'd15747,17'd65,17'd1291,17'd15748,17'd14082,17'd15749,17'd2627,17'd15750,17'd15751,17'd15752,17'd15753,17'd15754,17'd15755,17'd15756,17'd15508,17'd13450,17'd13450,17'd13591,17'd15757,17'd15758,17'd15759,17'd15258,17'd15760,17'd15761,17'd13326,17'd13325,17'd13325,17'd13595,17'd13596,17'd13838,17'd14098,17'd13597,17'd15762,17'd14469,17'd15763,17'd12527,17'd12527,17'd13093,17'd14621,17'd14764,17'd15764,17'd12361,17'd12362,17'd12530,17'd12530,17'd11627,17'd15640,17'd12066,17'd13841,17'd10563,17'd11087,17'd15765,17'd15766,17'd13843,17'd14219,17'd14473,17'd15641,17'd15641,17'd15767,17'd15386,17'd15387,17'd15768,17'd15769,17'd15770,17'd15771,17'd15772,17'd15773,17'd15527,17'd15774,17'd15775,17'd15776,17'd15777,17'd15778,17'd15779,17'd15780,17'd15781,17'd15782,17'd15783,17'd13106,17'd8702,17'd8856,17'd9589,17'd15784,17'd15785,17'd15786,17'd15787,17'd15788,17'd15789,17'd15790,17'd15791,17'd15409,17'd15661,17'd15280,17'd15544,17'd15792,17'd15032,17'd14236,17'd15793,17'd13226,17'd15794,17'd15795,17'd15796,17'd15797,17'd15550,17'd14658,17'd15287,17'd15798,17'd15799,17'd15800,17'd15553,17'd15559,17'd15801,17'd15802,17'd13504,17'd13996,17'd14513,17'd14253,17'd12706,17'd12236,17'd12240,17'd11788,17'd11949,17'd12714,17'd15803,17'd15804,17'd15805,17'd15806,17'd8873,17'd15178,17'd9482,17'd8726,17'd8886,17'd15807,17'd14134,17'd11667,17'd11958,17'd15433,17'd15570,17'd13517,17'd12579,17'd12579,17'd12580,17'd12419,17'd12258,17'd15808,17'd15809,17'd14002,17'd13362,17'd15810,17'd12262,17'd11963,17'd11806,17'd13882,17'd12414,17'd12859,17'd14672,17'd15811,17'd15687,17'd15687,17'd12415,17'd12859,17'd12575,17'd12861,17'd15052,17'd15569,17'd8724,17'd15812,17'd15813,17'd8259,17'd15442,17'd14390,17'd15814,17'd15188,17'd10180,17'd14938,17'd14270,17'd15575,17'd15306,17'd14393,17'd15815,17'd15816,17'd8117,17'd15817,17'd15818,17'd15819,17'd15820,17'd15201,17'd15821,17'd15822,17'd14275,17'd11289,17'd10874,17'd15823,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd135,17'd132,17'd132,17'd3512,17'd15824,17'd15825,17'd15826,17'd15827,17'd15828,17'd15829,17'd15830,17'd15831,17'd14284,17'd15585,17'd15832,17'd13270,17'd15216,17'd15833,17'd15834,17'd15835,17'd14838,17'd15836,17'd14706,17'd14287,17'd15837,17'd15838,17'd10054,17'd8764,17'd12611,17'd14035,17'd13159,17'd13159,17'd8614,17'd12138,17'd8762,17'd8762,17'd8614,17'd13159,17'd14958,17'd15839,17'd15840,17'd15841,17'd15842,17'd15715,17'd15843,17'd15716,17'd15844,17'd15718,17'd15086,17'd11295,17'd11551,17'd9504,17'd14161,17'd15594,17'd15328,17'd14846,17'd14415,17'd14161,17'd15594,17'd15594,17'd15594,17'd15594,17'd14713,17'd15327,17'd14417,17'd14160,17'd14159,17'd14159,17'd14159,17'd14846,17'd15845,17'd15846,17'd15467,17'd15719,17'd15847,17'd13787,17'd15709,17'd9381,17'd15598,17'd15848,17'd15849,17'd15601,17'd15850,17'd12756,17'd12460,17'd14569,17'd15722,17'd15851,17'd15473,17'd15222,17'd14569,17'd14569,17'd15603,17'd15604,17'd15604,17'd15723,17'd15852,17'd15723,17'd15475,17'd15475,17'd15093,17'd14421,17'd15339,17'd15339,17'd14722,17'd14571,17'd15725,17'd15607,17'd15853,17'd15854,17'd13923,17'd13923,17'd14971,17'd14970,17'd12760,17'd12160,17'd15855,17'd15856,17'd15857,17'd15858,17'd15859,17'd14427,17'd15613,17'd13681,17'd14053,17'd13927,17'd14055,17'd15860,17'd15861,17'd15231,17'd15862,17'd8507,17'd14586,17'd15233,17'd415,17'd415,17'd196,17'd418,17'd2102,17'd2246,17'd15863,17'd15864,17'd15865,17'd15622,17'd5366,17'd6869,17'd7516,17'd7684,17'd8018,17'd8170,17'd11444,17'd11444,17'd11191,17'd14984,17'd12319,17'd12487,17'd11723,17'd12489,17'd13425,17'd13425,17'd15866,17'd15866,17'd15238,17'd15238,17'd12776,17'd11330,17'd15867,17'd15867,17'd14064,17'd14181,17'd15489,17'd15108,17'd15108,17'd15108,17'd15868,17'd15624,17'd14596,17'd8325,17'd15869,17'd15870,17'd10080,17'd12322,17'd12922,17'd12492,17'd12182,17'd12182,17'd12492,17'd12642,17'd8810,17'd12493,17'd13294,17'd13427,17'd15871,17'd4060,17'd5788,17'd209,17'd406,17'd15872,17'd15873,17'd15874
},
'{
17'd466,17'd466,17'd12,17'd806,17'd25,17'd4,17'd6,17'd7,17'd3753,17'd3753,17'd5205,17'd5205,17'd5205,17'd5205,17'd3753,17'd3753,17'd7,17'd6,17'd5,17'd24,17'd23,17'd23,17'd23,17'd23,17'd5518,17'd5518,17'd20,17'd21,17'd9,17'd5512,17'd11063,17'd12925,17'd13431,17'd8347,17'd15875,17'd15628,17'd6588,17'd8825,17'd8670,17'd8815,17'd9272,17'd6106,17'd6426,17'd2421,17'd10260,17'd8814,17'd4089,17'd2594,17'd13428,17'd15876,17'd15877,17'd15878,17'd659,17'd985,17'd36,17'd36,17'd811,17'd295,17'd1553,17'd1836,17'd15879,17'd14871,17'd15366,17'd2269,17'd15880,17'd15881,17'd15882,17'd15883,17'd15884,17'd15885,17'd15886,17'd15887,17'd15888,17'd15889,17'd15890,17'd13199,17'd15891,17'd15892,17'd15893,17'd15894,17'd15895,17'd15896,17'd15639,17'd15259,17'd15761,17'd13326,17'd13325,17'd13326,17'd13596,17'd13838,17'd14098,17'd13597,17'd15762,17'd13092,17'd14469,17'd15763,17'd12527,17'd13093,17'd13211,17'd14764,17'd15764,17'd15764,17'd12362,17'd12815,17'd12218,17'd11478,17'd15897,17'd11229,17'd10111,17'd10427,17'd11915,17'd10943,17'd15898,17'd15899,17'd14219,17'd14346,17'd15641,17'd15384,17'd15767,17'd15900,17'd15901,17'd15261,17'd15769,17'd15902,17'd15010,17'd15903,17'd15904,17'd15905,17'd15906,17'd15907,17'd15908,17'd15909,17'd15777,17'd15910,17'd15911,17'd15912,17'd15913,17'd15914,17'd8700,17'd13612,17'd7590,17'd9851,17'd15784,17'd15915,17'd15916,17'd15917,17'd15918,17'd15919,17'd15920,17'd15921,17'd15922,17'd15923,17'd15924,17'd15280,17'd15281,17'd15411,17'd15662,17'd14237,17'd15925,17'd12548,17'd15664,17'd15926,17'd15927,17'd15928,17'd15929,17'd15930,17'd15798,17'd15931,17'd15932,17'd14369,17'd12704,17'd12565,17'd15933,17'd15802,17'd13995,17'd14513,17'd15674,17'd12236,17'd15934,17'd12088,17'd15935,17'd15936,17'd15937,17'd15938,17'd15939,17'd13137,17'd15940,17'd9345,17'd15941,17'd14675,17'd8569,17'd8886,17'd10175,17'd15566,17'd13138,17'd11806,17'd13252,17'd15942,17'd12995,17'd12109,17'd12579,17'd12579,17'd12580,17'd12580,17'd15809,17'd15808,17'd12998,17'd12858,17'd12262,17'd12262,17'd13362,17'd13135,17'd11960,17'd12414,17'd12859,17'd12415,17'd15687,17'd15687,17'd15687,17'd15687,17'd12415,17'd15434,17'd12414,17'd11667,17'd15943,17'd15944,17'd15945,17'd7951,17'd8425,17'd8259,17'd7620,17'd15946,17'd15947,17'd15948,17'd15949,17'd14269,17'd14816,17'd15950,17'd13529,17'd15951,17'd15952,17'd15953,17'd15954,17'd12124,17'd15955,17'd15956,17'd15957,17'd15958,17'd15959,17'd15960,17'd15961,17'd8132,17'd15823,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd135,17'd132,17'd135,17'd12127,17'd13903,17'd15962,17'd15963,17'd15964,17'd15965,17'd15966,17'd15967,17'd15968,17'd15969,17'd15332,17'd15970,17'd13394,17'd15971,17'd15972,17'd15834,17'd15973,17'd14555,17'd14706,17'd14956,17'd15080,17'd14156,17'd14413,17'd10505,17'd8764,17'd11994,17'd14035,17'd14958,17'd8614,17'd11987,17'd11987,17'd8762,17'd12137,17'd13159,17'd13159,17'd8614,17'd9223,17'd15714,17'd15974,17'd15975,17'd15715,17'd15976,17'd15977,17'd15593,17'd14159,17'd14415,17'd11295,17'd11295,17'd14161,17'd14161,17'd15594,17'd15214,17'd15328,17'd14161,17'd14161,17'd15594,17'd15594,17'd15594,17'd15594,17'd14713,17'd15327,17'd15978,17'd14417,17'd14160,17'd14160,17'd14160,17'd14159,17'd14710,17'd15845,17'd15979,17'd15980,17'd15216,17'd13271,17'd15981,17'd15982,17'd15090,17'd15470,17'd15471,17'd15983,17'd15984,17'd15985,17'd12757,17'd12899,17'd15474,17'd15473,17'd15986,17'd15987,17'd15474,17'd14569,17'd15603,17'd15852,17'd15852,17'd15604,17'd15852,17'd15604,17'd15603,17'd15603,17'd15605,17'd14570,17'd14421,17'd14571,17'd14722,17'd14421,17'd15988,17'd15988,17'd15607,17'd15989,17'd13799,17'd13799,17'd14971,17'd15094,17'd14301,17'd11853,17'd15990,17'd15855,17'd15991,17'd15227,17'd15992,17'd15730,17'd15993,17'd13681,17'd15994,17'd15995,17'd14055,17'd15996,17'd15997,17'd15998,17'd15999,17'd6418,17'd9123,17'd15233,17'd415,17'd1529,17'd197,17'd417,17'd1948,17'd2104,17'd12497,17'd15864,17'd16000,17'd15738,17'd3877,17'd6869,17'd7516,17'd7684,17'd14983,17'd8170,17'd11444,17'd11444,17'd11191,17'd11050,17'd12018,17'd12019,17'd11723,17'd12489,17'd13425,17'd13425,17'd15866,17'd15866,17'd15623,17'd15623,17'd12918,17'd11330,17'd15867,17'd16001,17'd14064,17'd14064,17'd15489,17'd15489,17'd15108,17'd15108,17'd15868,17'd15868,17'd15624,17'd8325,17'd15869,17'd15870,17'd11059,17'd9120,17'd12642,17'd12922,17'd12182,17'd12182,17'd12492,17'd12642,17'd8810,17'd11196,17'd13294,17'd16002,17'd9669,17'd16003,17'd6885,17'd233,17'd16004,17'd1398,17'd16005,17'd16006
},
'{
17'd3430,17'd13,17'd2423,17'd1275,17'd25,17'd4,17'd6,17'd6,17'd5205,17'd5205,17'd5205,17'd5205,17'd7,17'd6,17'd6,17'd6,17'd6,17'd5,17'd22,17'd23,17'd4,17'd8,17'd23,17'd5518,17'd2598,17'd20,17'd20,17'd21,17'd1413,17'd5513,17'd12781,17'd16007,17'd14987,17'd16008,17'd15744,17'd13813,17'd8661,17'd6900,17'd9136,17'd7892,17'd6105,17'd6428,17'd14068,17'd16009,17'd20,17'd3905,17'd1416,17'd2258,17'd3251,17'd3428,17'd16010,17'd16011,17'd471,17'd294,17'd294,17'd471,17'd295,17'd295,17'd1553,17'd1836,17'd58,17'd64,17'd487,17'd2127,17'd16012,17'd3116,17'd16013,17'd16014,17'd16015,17'd16016,17'd16017,17'd16018,17'd16019,17'd16020,17'd15890,17'd16021,17'd14091,17'd16022,17'd16023,17'd16024,17'd15896,17'd16025,17'd16026,17'd13716,17'd13596,17'd13595,17'd13595,17'd13595,17'd13596,17'd13716,17'd13597,17'd15762,17'd13598,17'd13092,17'd14469,17'd14469,17'd12527,17'd12528,17'd15137,17'd14891,17'd15764,17'd16027,17'd12362,17'd12362,17'd12956,17'd11478,17'd15640,17'd11229,17'd10111,17'd10563,17'd10944,17'd11231,17'd16028,17'd15524,17'd14347,17'd14768,17'd15641,17'd16029,17'd16030,17'd16031,17'd15261,17'd16032,17'd16033,17'd16034,17'd14895,17'd14897,17'd15773,17'd15906,17'd16035,17'd15529,17'd16036,17'd16037,17'd16038,17'd16039,17'd16040,17'd16041,17'd15022,17'd12822,17'd16042,17'd16043,17'd16044,17'd9589,17'd16045,17'd15916,17'd16046,17'd16047,17'd16048,17'd15659,17'd16049,17'd16050,17'd15922,17'd15923,17'd15924,17'd15280,17'd15545,17'd15411,17'd14362,17'd14114,17'd14363,17'd16051,17'd16052,17'd10710,17'd16053,17'd16054,17'd16055,17'd15288,17'd16056,17'd16057,17'd16058,17'd16059,17'd14373,17'd12709,17'd16060,17'd13129,17'd14372,17'd12705,17'd15675,17'd15934,17'd12089,17'd12710,17'd16061,17'd11656,17'd16062,17'd16063,17'd16064,17'd14806,17'd16065,17'd16066,17'd15941,17'd8878,17'd9046,17'd16067,17'd9339,17'd11134,17'd16068,17'd11960,17'd13252,17'd13518,17'd13763,17'd12577,17'd12109,17'd12579,17'd12579,17'd12995,17'd15809,17'd15809,17'd12857,17'd12996,17'd12115,17'd12262,17'd13362,17'd11806,17'd12419,17'd12414,17'd12859,17'd12415,17'd15687,17'd15687,17'd15571,17'd14672,17'd12859,17'd13514,17'd12577,17'd16069,17'd16070,17'd16071,17'd16072,17'd16073,17'd16074,17'd16075,17'd9890,17'd16076,17'd15947,17'd16077,17'd16078,17'd15194,17'd13528,17'd16079,17'd15695,17'd15444,17'd16080,17'd16081,17'd16082,17'd16083,17'd16084,17'd16085,17'd16086,17'd16087,17'd16088,17'd16089,17'd6530,17'd1045,17'd16090,17'd133,17'd132,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd542,17'd542,17'd132,17'd132,17'd135,17'd132,17'd134,17'd3811,17'd16091,17'd16092,17'd16093,17'd16094,17'd16095,17'd16096,17'd16097,17'd15831,17'd14152,17'd16098,17'd16099,17'd13271,17'd14558,17'd16100,17'd16101,17'd16102,17'd16103,17'd16104,17'd16105,17'd16106,17'd14704,17'd15080,17'd14555,17'd8457,17'd12611,17'd16107,17'd14035,17'd14035,17'd8916,17'd9767,17'd8762,17'd11987,17'd8614,17'd8456,17'd8916,17'd16108,17'd16109,17'd16110,17'd16111,17'd15325,17'd15324,17'd15212,17'd15211,17'd16112,17'd14710,17'd14415,17'd14415,17'd14161,17'd14161,17'd14038,17'd14708,17'd14708,17'd14161,17'd14161,17'd14415,17'd14415,17'd14709,17'd15328,17'd14159,17'd14160,17'd14295,17'd14295,17'd14416,17'd14416,17'd14294,17'd15718,17'd14293,17'd16113,17'd16114,17'd12604,17'd15463,17'd16115,17'd15981,17'd16116,17'd15457,17'd15332,17'd15848,17'd16117,17'd15984,17'd15985,17'd12756,17'd12460,17'd15221,17'd15474,17'd16118,17'd16118,17'd15604,17'd15603,17'd15603,17'd15852,17'd16118,17'd15852,17'd15852,17'd15852,17'd15852,17'd15604,17'd15603,17'd16119,17'd15336,17'd16120,17'd14421,17'd14421,17'd14421,17'd14722,17'd16121,17'd15726,17'd15854,17'd16122,17'd13925,17'd15094,17'd16123,17'd13678,17'd16124,17'd16125,17'd16126,17'd15343,17'd16127,17'd16128,17'd7505,17'd13411,17'd14727,17'd15995,17'd14973,17'd16129,17'd16130,17'd16131,17'd15618,17'd16132,17'd9123,17'd12644,17'd1529,17'd1529,17'd416,17'd196,17'd1947,17'd2103,17'd2398,17'd2565,17'd2745,17'd15738,17'd3877,17'd5502,17'd7516,17'd7685,17'd8169,17'd8019,17'd8795,17'd8795,17'd16133,17'd11050,17'd12018,17'd12319,17'd12488,17'd12489,17'd13425,17'd13691,17'd16134,17'd15866,17'd16134,17'd16134,17'd16135,17'd16001,17'd15867,17'd16001,17'd14064,17'd14064,17'd16136,17'd15489,17'd15108,17'd15108,17'd15868,17'd16137,17'd15868,17'd14596,17'd15869,17'd15870,17'd16138,17'd10256,17'd12492,17'd12922,17'd12492,17'd12492,17'd12492,17'd12492,17'd8810,17'd8810,17'd9121,17'd13294,17'd8644,17'd7209,17'd5192,17'd782,17'd16139,17'd614,17'd177,17'd16140
},
'{
17'd3430,17'd12,17'd1275,17'd465,17'd25,17'd4,17'd5,17'd6,17'd5205,17'd5205,17'd5205,17'd5205,17'd6,17'd6,17'd6,17'd6,17'd6,17'd24,17'd22,17'd23,17'd8,17'd8,17'd22,17'd16141,17'd2598,17'd20,17'd21,17'd9,17'd5647,17'd13062,17'd16142,17'd16143,17'd16008,17'd16008,17'd16144,17'd10659,17'd8973,17'd7380,17'd6105,17'd7892,17'd6732,17'd5797,17'd2421,17'd10260,17'd11,17'd17,17'd2257,17'd3252,17'd6420,17'd4428,17'd3427,17'd10925,17'd656,17'd656,17'd294,17'd471,17'd36,17'd985,17'd15363,17'd1836,17'd482,17'd668,17'd16145,17'd16146,17'd16147,17'd16013,17'd16148,17'd16149,17'd16150,17'd16151,17'd16152,17'd16153,17'd16154,17'd16155,17'd16156,17'd16157,17'd16158,17'd16159,17'd16160,17'd16161,17'd16162,17'd15762,17'd14098,17'd13716,17'd13596,17'd13595,17'd13595,17'd13596,17'd13716,17'd12356,17'd15762,17'd13092,17'd13092,17'd13092,17'd14469,17'd14469,17'd12528,17'd14890,17'd14764,17'd15764,17'd16163,17'd16027,17'd12362,17'd12362,17'd12956,17'd11627,17'd15640,17'd12066,17'd10691,17'd11087,17'd10944,17'd16164,17'd15899,17'd16165,17'd14346,17'd14892,17'd15767,17'd16166,17'd16167,17'd16031,17'd14765,17'd16168,17'd16169,17'd16170,17'd16171,17'd16172,17'd16173,17'd16174,17'd16175,17'd16176,17'd15909,17'd16037,17'd16177,17'd16178,17'd16041,17'd16179,17'd12822,17'd13611,17'd12685,17'd7428,17'd9588,17'd16180,17'd15915,17'd15916,17'd16181,17'd16182,17'd16183,17'd16184,17'd15790,17'd15921,17'd15922,17'd16185,17'd15924,17'd16186,17'd15545,17'd16187,17'd14237,17'd13226,17'd15160,17'd16188,17'd16189,17'd16190,17'd16191,17'd16192,17'd16193,17'd16194,17'd14917,17'd14368,17'd16195,17'd13237,17'd13753,17'd15555,17'd12400,17'd14253,17'd12558,17'd12558,17'd12087,17'd12088,17'd11788,17'd11790,17'd12247,17'd16196,17'd16197,17'd16198,17'd16199,17'd16200,17'd16201,17'd16202,17'd8884,17'd8886,17'd8567,17'd9038,17'd9341,17'd11133,17'd11667,17'd12420,17'd13252,17'd13365,17'd12252,17'd14808,17'd15184,17'd16203,17'd12579,17'd13517,17'd13365,17'd12111,17'd11806,17'd16204,17'd12115,17'd12262,17'd12996,17'd11960,17'd12109,17'd15434,17'd12415,17'd12860,17'd15687,17'd15687,17'd15571,17'd12860,17'd15434,17'd13514,17'd13882,17'd14673,17'd15566,17'd16205,17'd8254,17'd16206,17'd14813,17'd13141,17'd10746,17'd16207,17'd16208,17'd16209,17'd16210,17'd14270,17'd12267,17'd7958,17'd11676,17'd16211,17'd16212,17'd16213,17'd16214,17'd16215,17'd16216,17'd14539,17'd16217,17'd16218,17'd16219,17'd16220,17'd3025,17'd133,17'd133,17'd133,17'd132,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd132,17'd542,17'd542,17'd132,17'd132,17'd132,17'd132,17'd132,17'd2861,17'd16221,17'd16222,17'd16223,17'd16224,17'd16225,17'd16226,17'd14700,17'd16227,17'd14026,17'd15332,17'd16228,17'd13156,17'd15839,17'd16229,17'd16230,17'd16231,17'd16103,17'd16103,17'd16105,17'd16232,17'd16233,17'd14706,17'd16233,17'd9921,17'd12611,17'd16107,17'd16234,17'd8764,17'd10631,17'd10631,17'd8916,17'd11987,17'd8614,17'd12282,17'd10631,17'd15593,17'd16235,17'd16236,17'd15325,17'd16237,17'd15084,17'd15212,17'd15083,17'd14961,17'd16238,17'd14846,17'd14846,17'd14415,17'd14038,17'd14038,17'd14708,17'd14708,17'd14161,17'd14161,17'd14415,17'd14415,17'd15328,17'd15328,17'd14159,17'd14160,17'd14416,17'd14416,17'd14416,17'd14416,17'd14416,17'd14294,17'd14293,17'd16113,17'd14292,17'd16239,17'd15330,17'd15216,17'd16240,17'd16241,17'd16242,17'd15090,17'd16243,17'd16244,17'd16245,17'd15984,17'd15985,17'd15091,17'd15092,17'd15221,17'd15852,17'd16118,17'd16118,17'd15604,17'd15723,17'd15852,17'd16118,17'd16118,17'd16118,17'd16246,17'd16246,17'd15852,17'd15723,17'd15475,17'd15336,17'd15337,17'd14571,17'd14421,17'd14421,17'd14722,17'd16247,17'd15725,17'd15989,17'd16122,17'd13925,17'd14971,17'd16123,17'd12307,17'd15855,17'd16248,17'd16249,17'd16126,17'd16250,17'd16251,17'd7504,17'd13411,17'd14727,17'd15995,17'd16252,17'd16253,17'd16254,17'd15230,17'd16255,17'd15862,17'd8186,17'd16256,17'd413,17'd1529,17'd416,17'd197,17'd14977,17'd2102,17'd2397,17'd2399,17'd2564,17'd16257,17'd5036,17'd5502,17'd7343,17'd7346,17'd8169,17'd8171,17'd8795,17'd8795,17'd16133,17'd16133,17'd9253,17'd12319,17'd12487,17'd13423,17'd13059,17'd13691,17'd16258,17'd16134,17'd16134,17'd16134,17'd15866,17'd16259,17'd16001,17'd15867,17'd14063,17'd14063,17'd16136,17'd15489,17'd15489,17'd15108,17'd16137,17'd16137,17'd15868,17'd15624,17'd16260,17'd15870,17'd16138,17'd10256,17'd12492,17'd12922,17'd12642,17'd12492,17'd12182,17'd12492,17'd8810,17'd8810,17'd9121,17'd16261,17'd16262,17'd8184,17'd6885,17'd794,17'd1547,17'd613,17'd16263,17'd16264
},
'{
17'd3430,17'd12,17'd808,17'd9,17'd23,17'd23,17'd5,17'd5,17'd5205,17'd5205,17'd5205,17'd3753,17'd5,17'd5,17'd4,17'd8,17'd23,17'd23,17'd23,17'd23,17'd23,17'd23,17'd20,17'd2598,17'd2598,17'd21,17'd9,17'd1413,17'd5514,17'd13574,17'd16007,17'd16265,17'd15493,17'd15628,17'd8195,17'd6427,17'd6900,17'd8511,17'd6595,17'd8815,17'd6588,17'd807,17'd15494,17'd8814,17'd18,17'd17,17'd2257,17'd10547,17'd3901,17'd4738,17'd11071,17'd10669,17'd32,17'd1130,17'd656,17'd294,17'd12504,17'd985,17'd15363,17'd989,17'd14450,17'd2613,17'd16266,17'd16267,17'd3116,17'd16268,17'd16269,17'd16270,17'd16271,17'd16272,17'd16273,17'd16274,17'd13314,17'd16275,17'd16276,17'd16277,17'd16278,17'd16279,17'd16280,17'd16281,17'd16282,17'd12677,17'd12356,17'd13596,17'd13595,17'd16283,17'd16283,17'd15761,17'd13716,17'd13597,17'd13598,17'd12954,17'd13092,17'd12527,17'd16284,17'd16284,17'd12529,17'd16285,17'd16286,17'd14891,17'd14622,17'd16287,17'd12361,17'd12361,17'd11627,17'd11627,17'd15640,17'd15897,17'd16288,17'd11087,17'd10945,17'd16289,17'd15902,17'd16290,17'd14346,17'd14892,17'd15767,17'd15900,17'd15260,17'd15260,17'd14768,17'd16168,17'd16028,17'd16291,17'd16292,17'd14898,17'd15648,17'd15144,17'd15268,17'd15269,17'd15650,17'd15650,17'd16177,17'd16177,17'd16293,17'd14782,17'd9016,17'd9165,17'd12071,17'd16294,17'd9589,17'd16295,17'd16296,17'd15916,17'd16182,17'd16297,17'd16298,17'd16298,17'd15790,17'd15543,17'd15279,17'd15279,17'd16186,17'd15156,17'd15545,17'd16187,17'd13985,17'd13340,17'd12832,17'd16299,17'd16300,17'd16301,17'd10582,17'd16302,17'd16303,17'd16304,17'd16305,17'd11377,17'd13237,17'd16306,17'd13754,17'd16307,17'd15169,17'd16308,17'd13353,17'd13632,17'd16309,17'd11936,17'd12712,17'd16310,17'd16311,17'd16312,17'd16313,17'd12862,17'd16314,17'd10172,17'd16315,17'd16316,17'd16317,17'd9195,17'd8567,17'd16318,17'd16319,17'd16320,17'd11806,17'd16321,17'd13136,17'd13763,17'd16322,17'd16323,17'd15054,17'd16324,17'd12253,17'd12417,17'd13365,17'd12420,17'd16325,17'd16326,17'd12115,17'd13362,17'd12113,17'd12111,17'd12413,17'd13514,17'd12997,17'd14672,17'd15571,17'd16327,17'd15571,17'd14672,17'd12859,17'd12578,17'd11960,17'd11399,17'd16328,17'd11531,17'd16329,17'd8425,17'd16330,17'd16331,17'd16332,17'd16333,17'd16334,17'd16335,17'd15690,17'd14266,17'd13894,17'd16336,17'd11676,17'd7466,17'd16337,17'd16338,17'd16339,17'd16340,17'd16341,17'd14823,17'd16342,17'd14399,17'd14276,17'd4163,17'd356,17'd132,17'd131,17'd11541,17'd132,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd542,17'd542,17'd132,17'd132,17'd131,17'd132,17'd132,17'd3168,17'd6057,17'd12598,17'd9497,17'd16343,17'd16344,17'd16345,17'd13020,17'd13910,17'd13911,17'd16346,17'd16099,17'd13667,17'd16347,17'd16348,17'd16349,17'd16350,17'd16351,17'd16352,17'd16105,17'd16232,17'd16353,17'd14556,17'd14556,17'd14957,17'd14035,17'd12895,17'd16234,17'd16354,17'd11297,17'd11297,17'd8917,17'd8763,17'd14035,17'd8764,17'd10885,17'd16355,17'd16356,17'd15843,17'd15465,17'd16357,17'd16358,17'd15212,17'd15212,17'd14962,17'd14963,17'd14964,17'd14293,17'd14846,17'd14158,17'd14038,17'd9370,17'd9370,17'd14161,17'd15086,17'd15086,17'd15086,17'd14159,17'd14159,17'd15718,17'd14294,17'd16359,17'd16360,17'd16361,17'd16361,17'd16361,17'd16360,17'd16362,17'd16363,17'd14293,17'd14710,17'd12604,17'd9222,17'd14965,17'd14029,17'd16364,17'd16346,17'd16365,17'd15848,17'd16366,17'd16367,17'd16368,17'd16369,17'd15091,17'd13036,17'd15723,17'd15852,17'd16246,17'd16118,17'd15604,17'd15604,17'd15852,17'd16246,17'd16118,17'd16246,17'd16370,17'd16118,17'd15604,17'd15723,17'd15475,17'd15336,17'd12000,17'd12295,17'd14421,17'd14421,17'd16371,17'd16247,17'd15608,17'd15854,17'd14970,17'd13925,17'd14423,17'd12468,17'd15855,17'd16248,17'd16249,17'd16249,17'd16372,17'd16373,17'd16374,17'd13411,17'd16375,17'd15995,17'd16376,17'd16377,17'd16378,17'd16379,17'd16380,17'd16381,17'd6258,17'd16382,17'd413,17'd1529,17'd416,17'd419,17'd1811,17'd1948,17'd2241,17'd2398,17'd14737,17'd15865,17'd3574,17'd5635,17'd6576,17'd7346,17'd8169,17'd8171,17'd8491,17'd8491,17'd16133,17'd11050,17'd10076,17'd11722,17'd11593,17'd12178,17'd13425,17'd13425,17'd16134,17'd16134,17'd16383,17'd16384,17'd15866,17'd16135,17'd16259,17'd15867,17'd11330,17'd14063,17'd16136,17'd15489,17'd15489,17'd15489,17'd16137,17'd16137,17'd16137,17'd15624,17'd16260,17'd15869,17'd16138,17'd10256,17'd12182,17'd12642,17'd16385,17'd12492,17'd8655,17'd7034,17'd8330,17'd8503,17'd6089,17'd16261,17'd16262,17'd16386,17'd5788,17'd794,17'd247,17'd433,17'd16387,17'd16388
},
'{
17'd3430,17'd806,17'd808,17'd16389,17'd25,17'd22,17'd23,17'd5,17'd7,17'd5205,17'd3753,17'd5,17'd24,17'd23,17'd4,17'd8,17'd22,17'd23,17'd4,17'd23,17'd22,17'd20,17'd20,17'd20,17'd20,17'd25,17'd1413,17'd5647,17'd5513,17'd10916,17'd12782,17'd16390,17'd16391,17'd16144,17'd7893,17'd7724,17'd6900,17'd6105,17'd9272,17'd8518,17'd6426,17'd4242,17'd15494,17'd806,17'd3905,17'd2257,17'd2258,17'd2935,17'd4245,17'd3904,17'd2592,17'd10546,17'd292,17'd32,17'd656,17'd34,17'd16392,17'd659,17'd1837,17'd825,17'd831,17'd2615,17'd2128,17'd1990,17'd16393,17'd16394,17'd16395,17'd16396,17'd16397,17'd16398,17'd16399,17'd16400,17'd12942,17'd16275,17'd16401,17'd16402,17'd16403,17'd16404,17'd16161,17'd16405,17'd16406,17'd16407,17'd12215,17'd13838,17'd15136,17'd15136,17'd16408,17'd15761,17'd14344,17'd13597,17'd13092,17'd12954,17'd12527,17'd12527,17'd16284,17'd12679,17'd14890,17'd15137,17'd14891,17'd15764,17'd14470,17'd14470,17'd12361,17'd13840,17'd11627,17'd12956,17'd15640,17'd16288,17'd16409,17'd10944,17'd16410,17'd15899,17'd16411,17'd14346,17'd14766,17'd14892,17'd15767,17'd15900,17'd15260,17'd15386,17'd14768,17'd14219,17'd16412,17'd16413,17'd16414,17'd16415,17'd16174,17'd15267,17'd15776,17'd16416,17'd15650,17'd15650,17'd16177,17'd16417,17'd15399,17'd13105,17'd9165,17'd11920,17'd7428,17'd15402,17'd9993,17'd16418,17'd16418,17'd16419,17'd16183,17'd15790,17'd15790,17'd15790,17'd15921,17'd15543,17'd16420,17'd16186,17'd16186,17'd15157,17'd16421,17'd16422,17'd13226,17'd12077,17'd15664,17'd10709,17'd16423,17'd16424,17'd16425,17'd16302,17'd16426,17'd16427,17'd16428,17'd16429,17'd13996,17'd13753,17'd13752,17'd16430,17'd16431,17'd16432,17'd13632,17'd16433,17'd11786,17'd12850,17'd11799,17'd13878,17'd16312,17'd16434,17'd16435,17'd16436,17'd9479,17'd16437,17'd16438,17'd16439,17'd16440,17'd16067,17'd16441,17'd13887,17'd10741,17'd14810,17'd11961,17'd16321,17'd12420,17'd12110,17'd13364,17'd13363,17'd14130,17'd16324,17'd12253,17'd12417,17'd12995,17'd12420,17'd16442,17'd16326,17'd12115,17'd13362,17'd12420,17'd12109,17'd15434,17'd12860,17'd12860,17'd14672,17'd15571,17'd15571,17'd15571,17'd14672,17'd12859,17'd16443,17'd13520,17'd11400,17'd16440,17'd12426,17'd8583,17'd16444,17'd14936,17'd16445,17'd16446,17'd9622,17'd16447,17'd16448,17'd15437,17'd13528,17'd12121,17'd16449,17'd14142,17'd16450,17'd16451,17'd16452,17'd16453,17'd16454,17'd16455,17'd16456,17'd16457,17'd16458,17'd11289,17'd356,17'd130,17'd132,17'd11541,17'd11541,17'd132,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd135,17'd132,17'd3168,17'd6831,17'd16459,17'd16460,17'd16461,17'd16462,17'd16463,17'd16464,17'd16465,17'd15455,17'd16346,17'd16466,17'd13396,17'd16467,17'd12284,17'd16468,17'd16350,17'd16469,17'd16470,17'd16471,17'd16232,17'd16104,17'd16353,17'd14556,17'd13548,17'd16234,17'd12896,17'd10202,17'd16354,17'd16472,17'd16472,17'd8917,17'd8763,17'd8763,17'd16354,17'd16473,17'd16474,17'd15976,17'd15464,17'd16357,17'd16475,17'd16476,17'd16477,17'd15213,17'd16358,17'd14963,17'd16112,17'd14846,17'd14561,17'd14158,17'd14038,17'd9370,17'd9370,17'd14161,17'd15086,17'd15327,17'd14160,17'd16478,17'd16478,17'd16478,17'd14294,17'd15718,17'd14294,17'd14295,17'd16479,17'd16361,17'd16360,17'd16480,17'd16362,17'd14293,17'd15845,17'd12604,17'd12604,17'd9222,17'd15217,17'd16481,17'd16482,17'd16483,17'd16243,17'd16484,17'd16485,17'd16486,17'd16369,17'd12757,17'd13036,17'd15724,17'd15852,17'd16246,17'd16246,17'd15852,17'd15723,17'd15852,17'd16246,17'd15852,17'd16118,17'd16246,17'd16118,17'd15852,17'd15852,17'd15723,17'd15475,17'd13162,17'd12460,17'd14421,17'd14571,17'd16371,17'd16371,17'd15607,17'd16487,17'd14971,17'd13925,17'd14423,17'd12162,17'd16488,17'd16248,17'd16125,17'd16249,17'd16126,17'd16489,17'd15730,17'd13283,17'd13285,17'd14054,17'd16376,17'd16377,17'd16490,17'd15346,17'd16491,17'd15232,17'd16492,17'd5776,17'd14178,17'd413,17'd415,17'd419,17'd197,17'd1948,17'd2241,17'd2241,17'd2399,17'd2745,17'd6087,17'd3877,17'd4872,17'd6724,17'd7685,17'd7856,17'd8491,17'd8491,17'd9253,17'd11191,17'd9405,17'd11592,17'd11593,17'd12488,17'd12178,17'd13425,17'd13691,17'd16134,17'd15866,17'd16493,17'd15866,17'd16134,17'd16135,17'd16001,17'd11330,17'd14063,17'd16136,17'd15489,17'd15489,17'd15489,17'd16137,17'd15868,17'd16137,17'd15868,17'd14596,17'd15869,17'd11059,17'd10256,17'd12182,17'd12642,17'd16494,17'd12492,17'd7034,17'd7034,17'd8330,17'd8503,17'd10910,17'd16261,17'd9803,17'd16495,17'd4422,17'd794,17'd16139,17'd614,17'd16496,17'd16497
},
'{
17'd16498,17'd806,17'd651,17'd465,17'd1275,17'd2933,17'd977,17'd978,17'd7373,17'd7215,17'd16009,17'd16009,17'd16009,17'd2421,17'd2591,17'd2933,17'd10260,17'd4242,17'd23,17'd25,17'd21,17'd20,17'd20,17'd20,17'd22,17'd24,17'd5,17'd7216,17'd12925,17'd13063,17'd8347,17'd15743,17'd16265,17'd13574,17'd8347,17'd13183,17'd8815,17'd9137,17'd7380,17'd6435,17'd465,17'd10260,17'd16499,17'd16500,17'd13,17'd1127,17'd2422,17'd2935,17'd7545,17'd2422,17'd3429,17'd3593,17'd292,17'd33,17'd11071,17'd12196,17'd16501,17'd295,17'd1700,17'd667,17'd2613,17'd13581,17'd14605,17'd16502,17'd16503,17'd16504,17'd16505,17'd16506,17'd16507,17'd15125,17'd16508,17'd13197,17'd13198,17'd16509,17'd15128,17'd16510,17'd16511,17'd16512,17'd16513,17'd16514,17'd16025,17'd16515,17'd11224,17'd16516,17'd16516,17'd11909,17'd13838,17'd13716,17'd13597,17'd13462,17'd13092,17'd13092,17'd12813,17'd12813,17'd13093,17'd12955,17'd16517,17'd13969,17'd12361,17'd12218,17'd12530,17'd12530,17'd12530,17'd12530,17'd12956,17'd11627,17'd11361,17'd10691,17'd16518,17'd16164,17'd16519,17'd15524,17'd14346,17'd16030,17'd15641,17'd15641,17'd16520,17'd16521,17'd14766,17'd14892,17'd16165,17'd16522,17'd16523,17'd16524,17'd16525,17'd16526,17'd16527,17'd16528,17'd16037,17'd16529,17'd16177,17'd16530,17'd16040,17'd15272,17'd14358,17'd12822,17'd12370,17'd7428,17'd9589,17'd16180,17'd16419,17'd16531,17'd16532,17'd16533,17'd16534,17'd16535,17'd16536,17'd15543,17'd15791,17'd16537,17'd16186,17'd16186,17'd15544,17'd15030,17'd16538,17'd14113,17'd12831,17'd12549,17'd16052,17'd16539,17'd16540,17'd16541,17'd16542,17'd16543,17'd16544,17'd16545,17'd12702,17'd12397,17'd15672,17'd14662,17'd14252,17'd16546,17'd16546,17'd12842,17'd12847,17'd12560,17'd12850,17'd16547,17'd15293,17'd15803,17'd16548,17'd13000,17'd16436,17'd16549,17'd16550,17'd16551,17'd16201,17'd16552,17'd10175,17'd8873,17'd16553,17'd16554,17'd16555,17'd13362,17'd11960,17'd12420,17'd12420,17'd12419,17'd12414,17'd12414,17'd12109,17'd12579,17'd12579,17'd12579,17'd12580,17'd15053,17'd16204,17'd12262,17'd13362,17'd16204,17'd16321,17'd12415,17'd16556,17'd16557,17'd16558,17'd12860,17'd16559,17'd14524,17'd16560,17'd13642,17'd12859,17'd13882,17'd13254,17'd16561,17'd16562,17'd16563,17'd16564,17'd16565,17'd10746,17'd16332,17'd7947,17'd16566,17'd16567,17'd15438,17'd16568,17'd7957,17'd7793,17'd16569,17'd16570,17'd16571,17'd16572,17'd16573,17'd16574,17'd16575,17'd16576,17'd16577,17'd16578,17'd14016,17'd1197,17'd1197,17'd1197,17'd1045,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd130,17'd130,17'd130,17'd132,17'd132,17'd134,17'd3168,17'd16579,17'd16580,17'd16581,17'd16582,17'd14949,17'd16583,17'd16584,17'd15830,17'd16585,17'd16364,17'd16586,17'd14552,17'd12889,17'd8458,17'd8617,17'd16587,17'd16588,17'd16589,17'd16590,17'd16591,17'd16592,17'd16353,17'd14706,17'd13669,17'd8770,17'd8614,17'd8763,17'd11694,17'd10048,17'd8917,17'd10202,17'd11987,17'd16354,17'd10048,17'd15085,17'd16593,17'd16594,17'd15213,17'd15464,17'd16595,17'd16596,17'd16597,17'd16598,17'd16477,17'd16599,17'd14297,17'd11295,17'd11831,17'd10884,17'd15328,17'd9504,17'd9504,17'd14297,17'd14713,17'd16478,17'd15844,17'd15977,17'd15977,17'd15211,17'd16478,17'd14417,17'd14160,17'd16600,17'd16601,17'd16602,17'd16479,17'd16360,17'd15593,17'd16113,17'd14846,17'd14846,17'd15329,17'd12604,17'd9222,17'd15847,17'd16603,17'd16604,17'd16605,17'd16606,17'd16607,17'd16608,17'd16609,17'd15092,17'd13036,17'd16610,17'd16611,17'd15986,17'd16612,17'd16613,17'd15987,17'd15473,17'd15986,17'd16370,17'd16246,17'd16246,17'd16370,17'd16246,17'd15604,17'd16614,17'd15723,17'd14569,17'd13035,17'd14722,17'd14421,17'd15988,17'd16371,17'd16121,17'd15608,17'd15727,17'd15610,17'd16615,17'd14051,17'd16616,17'd16617,17'd16618,17'd16249,17'd14426,17'd16619,17'd15730,17'd14304,17'd13284,17'd13050,17'd16620,17'd16621,17'd14171,17'd16622,17'd15347,17'd15348,17'd16623,17'd7365,17'd12496,17'd193,17'd422,17'd416,17'd197,17'd196,17'd1248,17'd1248,17'd2397,17'd15235,17'd15349,17'd16624,17'd7028,17'd7028,17'd7346,17'd7856,17'd8796,17'd8019,17'd9405,17'd9405,17'd10076,17'd12018,17'd10077,17'd12487,17'd12488,17'd12489,17'd13424,17'd13425,17'd15623,17'd15623,17'd16134,17'd16134,17'd16625,17'd16626,17'd11330,17'd11330,17'd16627,17'd16136,17'd15489,17'd15108,17'd15108,17'd15108,17'd16628,17'd16629,17'd16630,17'd13692,17'd9542,17'd7692,17'd7034,17'd8503,17'd10910,17'd8810,17'd9120,17'd12322,17'd12492,17'd12493,17'd11196,17'd10910,17'd10793,17'd16631,17'd16632,17'd623,17'd1826,17'd16633,17'd16634,17'd16635
},
'{
17'd16636,17'd1275,17'd465,17'd465,17'd1275,17'd1275,17'd977,17'd807,17'd978,17'd7215,17'd16009,17'd2421,17'd2421,17'd2591,17'd1275,17'd8814,17'd4242,17'd4242,17'd25,17'd25,17'd10,17'd11,17'd20,17'd20,17'd22,17'd5,17'd7,17'd12648,17'd12781,17'd13063,17'd6427,17'd7724,17'd12925,17'd10916,17'd13431,17'd8670,17'd8815,17'd7892,17'd8973,17'd7381,17'd465,17'd2933,17'd16499,17'd16500,17'd3430,17'd1127,17'd2422,17'd2935,17'd4886,17'd4247,17'd2597,17'd3752,17'd292,17'd33,17'd33,17'd11071,17'd11888,17'd1694,17'd990,17'd16637,17'd2792,17'd16638,17'd16639,17'd16640,17'd16641,17'd16642,17'd16643,17'd16644,17'd16645,17'd16646,17'd16647,17'd16648,17'd13198,17'd16649,17'd14760,17'd16650,17'd16651,17'd16652,17'd16653,17'd16654,17'd16655,17'd16656,17'd16515,17'd16515,17'd16516,17'd16516,17'd16657,17'd13597,17'd13462,17'd14469,17'd13092,17'd13092,17'd12813,17'd13093,17'd13211,17'd14470,17'd16658,17'd12532,17'd12361,17'd12362,17'd12530,17'd12360,17'd12360,17'd12360,17'd12956,17'd11361,17'd10427,17'd10816,17'd15765,17'd16659,17'd15524,17'd14765,17'd15641,17'd16030,17'd16030,17'd16030,17'd15260,17'd15386,17'd14766,17'd14346,17'd15644,17'd16660,17'd16661,17'd16662,17'd15017,17'd16527,17'd15145,17'd16036,17'd16663,17'd16663,17'd16178,17'd16177,17'd16664,17'd16665,17'd13104,17'd9165,17'd16666,17'd15402,17'd9993,17'd16045,17'd16419,17'd16667,17'd16668,17'd16669,17'd16534,17'd16535,17'd16670,17'd15791,17'd15922,17'd16671,17'd16186,17'd15156,17'd15281,17'd15031,17'd15662,17'd16672,17'd16673,17'd10824,17'd10826,17'd16190,17'd16674,17'd16675,17'd16676,17'd16677,17'd16055,17'd11109,17'd12843,17'd13996,17'd14662,17'd14124,17'd14799,17'd14249,17'd14661,17'd12397,17'd11935,17'd12089,17'd16678,17'd16679,17'd12249,17'd11956,17'd11666,17'd15427,17'd16680,17'd15682,17'd16681,17'd9041,17'd10336,17'd16682,17'd8874,17'd15944,17'd15180,17'd16683,17'd11965,17'd12996,17'd13761,17'd11960,17'd12420,17'd12580,17'd12417,17'd12417,17'd12417,17'd12417,17'd12579,17'd12109,17'd13761,17'd13135,17'd13362,17'd12262,17'd15186,17'd12996,17'd14807,17'd16557,17'd16684,17'd16684,17'd16558,17'd16685,17'd13361,17'd14524,17'd16560,17'd16686,17'd12859,17'd15299,17'd16687,17'd10334,17'd12587,17'd16688,17'd16689,17'd10609,17'd15693,17'd16690,17'd16691,17'd13140,17'd15442,17'd16692,17'd16693,17'd12729,17'd16694,17'd14142,17'd16695,17'd16696,17'd16697,17'd16698,17'd16454,17'd16085,17'd16699,17'd11977,17'd10874,17'd11289,17'd1197,17'd1197,17'd1045,17'd133,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd130,17'd130,17'd130,17'd130,17'd134,17'd132,17'd132,17'd357,17'd3027,17'd16700,17'd7816,17'd16701,17'd16702,17'd16703,17'd14699,17'd16704,17'd16705,17'd16706,17'd16707,17'd14703,17'd8923,17'd8295,17'd16708,17'd16709,17'd16710,17'd16711,17'd16712,17'd16713,17'd16714,17'd14288,17'd14033,17'd13669,17'd16715,17'd8456,17'd10202,17'd11694,17'd16716,17'd16717,17'd10202,17'd11987,17'd16354,17'd16718,17'd15085,17'd16594,17'd16719,17'd16476,17'd16595,17'd16720,17'd16721,17'd16722,17'd16723,17'd16724,17'd16599,17'd14715,17'd11551,17'd11831,17'd10884,17'd15328,17'd14161,17'd9504,17'd14419,17'd15327,17'd16725,17'd16726,17'd16727,17'd16727,17'd16728,17'd16729,17'd16730,17'd14160,17'd16600,17'd16601,17'd16602,17'd16361,17'd15844,17'd15593,17'd15718,17'd14159,17'd14710,17'd15846,17'd12604,17'd15330,17'd12886,17'd12887,17'd16603,17'd16466,17'd16731,17'd16732,17'd16117,17'd16733,17'd15091,17'd12295,17'd13036,17'd16610,17'd15987,17'd15986,17'd16613,17'd15986,17'd15987,17'd15473,17'd16118,17'd16246,17'd16370,17'd16370,17'd16246,17'd16118,17'd16734,17'd16614,17'd14569,17'd13035,17'd14722,17'd14421,17'd15988,17'd16371,17'd16371,17'd15607,17'd16735,17'd15609,17'd12906,17'd12761,17'd12468,17'd16488,17'd16618,17'd16736,17'd16737,17'd16738,17'd15730,17'd14576,17'd16739,17'd13050,17'd16620,17'd16621,17'd14171,17'd16622,17'd15347,17'd15483,17'd16132,17'd7365,17'd5630,17'd412,17'd598,17'd2763,17'd419,17'd197,17'd1384,17'd1384,17'd2241,17'd14737,17'd15865,17'd16740,17'd6869,17'd5365,17'd7516,17'd7856,17'd8796,17'd8796,17'd9405,17'd9405,17'd10076,17'd12018,17'd10391,17'd10077,17'd12320,17'd15488,17'd13424,17'd12489,17'd13425,17'd15352,17'd16134,17'd15866,17'd16741,17'd16742,17'd11330,17'd11330,17'd16627,17'd16136,17'd15489,17'd15489,17'd15108,17'd15108,17'd16629,17'd16629,17'd16743,17'd8179,17'd9411,17'd7523,17'd9800,17'd8810,17'd10910,17'd8810,17'd9120,17'd9120,17'd12182,17'd11879,17'd11196,17'd10910,17'd12324,17'd16631,17'd16744,17'd623,17'd1826,17'd16745,17'd16633,17'd16746
},
'{
17'd806,17'd283,17'd283,17'd3,17'd806,17'd1275,17'd977,17'd977,17'd2421,17'd4242,17'd4242,17'd978,17'd2421,17'd2933,17'd2423,17'd16747,17'd4242,17'd16009,17'd4242,17'd2933,17'd11,17'd11,17'd20,17'd5518,17'd24,17'd6,17'd10658,17'd10796,17'd12781,17'd13063,17'd13297,17'd13181,17'd13062,17'd13063,17'd12926,17'd16748,17'd6900,17'd7058,17'd6596,17'd4732,17'd1275,17'd8814,17'd16500,17'd16749,17'd3430,17'd4247,17'd3250,17'd2422,17'd1689,17'd1127,17'd2596,17'd469,17'd2940,17'd2943,17'd3253,17'd3103,17'd2939,17'd1971,17'd824,17'd832,17'd2271,17'd2130,17'd16750,17'd16751,17'd16752,17'd16753,17'd16754,17'd16755,17'd16756,17'd16757,17'd13314,17'd16275,17'd16758,17'd16157,17'd16759,17'd16760,17'd16761,17'd16653,17'd16762,17'd15896,17'd16763,17'd16656,17'd16515,17'd16764,17'd16516,17'd16516,17'd14098,17'd13462,17'd13462,17'd14469,17'd13092,17'd12527,17'd13093,17'd12955,17'd14621,17'd14891,17'd13969,17'd16765,17'd12361,17'd12361,17'd12530,17'd12530,17'd12360,17'd12360,17'd11627,17'd11764,17'd11362,17'd16766,17'd16410,17'd16767,17'd16169,17'd14347,17'd14474,17'd16030,17'd15386,17'd15260,17'd15260,17'd14768,17'd16768,17'd16769,17'd16770,17'd16771,17'd16772,17'd16525,17'd16773,17'd16774,17'd16176,17'd15909,17'd16775,17'd16776,17'd16178,17'd16777,17'd16778,17'd16779,17'd9016,17'd12370,17'd7428,17'd16044,17'd9589,17'd16780,17'd16781,17'd16782,17'd16533,17'd16669,17'd16534,17'd16670,17'd15543,17'd15791,17'd16185,17'd16185,17'd15544,17'd15281,17'd15031,17'd15032,17'd14362,17'd13111,17'd11490,17'd16783,17'd16784,17'd16785,17'd16786,17'd16787,17'd16676,17'd16788,17'd13872,17'd12561,17'd12236,17'd12849,17'd16789,17'd14371,17'd16432,17'd16546,17'd12235,17'd16790,17'd15934,17'd12711,17'd11655,17'd16196,17'd11955,17'd16791,17'd16792,17'd10478,17'd16793,17'd16794,17'd8883,17'd16795,17'd10173,17'd9481,17'd9345,17'd15569,17'd10743,17'd16796,17'd13762,17'd13883,17'd12419,17'd12420,17'd16321,17'd12109,17'd12417,17'd13517,17'd12579,17'd14807,17'd12580,17'd12580,17'd11960,17'd12996,17'd12262,17'd12262,17'd16797,17'd12113,17'd12418,17'd16557,17'd16684,17'd16327,17'd16558,17'd12860,17'd16798,17'd16799,17'd16686,17'd14524,17'd12578,17'd11667,17'd10330,17'd10175,17'd9745,17'd16800,17'd16801,17'd16802,17'd13765,17'd16803,17'd11968,17'd16804,17'd14391,17'd10482,17'd14532,17'd15695,17'd16805,17'd16806,17'd16807,17'd14940,17'd16808,17'd16809,17'd16341,17'd11004,17'd16810,17'd16811,17'd889,17'd1197,17'd1481,17'd1481,17'd133,17'd133,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd542,17'd133,17'd132,17'd130,17'd130,17'd134,17'd132,17'd132,17'd131,17'd2866,17'd14826,17'd16812,17'd16813,17'd4009,17'd16814,17'd16815,17'd16816,17'd16817,17'd16818,17'd16481,17'd16819,17'd15460,17'd8458,17'd16820,17'd16821,17'd16822,17'd16823,17'd16824,17'd16825,17'd16714,17'd16104,17'd14555,17'd13669,17'd14030,17'd12447,17'd9642,17'd11694,17'd16716,17'd9642,17'd8762,17'd8916,17'd9223,17'd16718,17'd15085,17'd16594,17'd16826,17'd15841,17'd16827,17'd16828,17'd16829,17'd16830,17'd16831,17'd16477,17'd15326,17'd14161,17'd11295,17'd11831,17'd14709,17'd15328,17'd14161,17'd14161,17'd14714,17'd15327,17'd15844,17'd16726,17'd16832,17'd16236,17'd16833,17'd16834,17'd16478,17'd14416,17'd14416,17'd16360,17'd16361,17'd16835,17'd15844,17'd15844,17'd14416,17'd14294,17'd14293,17'd16836,17'd16114,17'd16114,17'd15979,17'd12605,17'd16837,17'd16604,17'd16838,17'd16839,17'd16244,17'd16733,17'd16840,17'd15091,17'd15091,17'd16841,17'd16611,17'd16842,17'd15986,17'd16612,17'd16246,17'd15604,17'd16843,17'd16844,17'd16845,17'd16844,17'd16246,17'd16246,17'd16846,17'd16614,17'd15222,17'd13035,17'd14722,17'd14722,17'd16121,17'd16247,17'd16371,17'd16247,17'd16847,17'd15727,17'd12906,17'd12469,17'd12163,17'd15611,17'd16848,17'd16849,17'd16850,17'd14854,17'd16851,17'd15614,17'd12907,17'd16852,17'd13414,17'd16377,17'd16853,17'd16622,17'd16491,17'd16854,17'd16855,17'd4882,17'd6415,17'd412,17'd952,17'd422,17'd421,17'd941,17'd945,17'd1105,17'd2099,17'd2399,17'd16856,17'd15486,17'd5366,17'd5365,17'd7343,17'd14983,17'd8171,17'd8019,17'd9405,17'd10076,17'd10076,17'd12018,17'd10391,17'd10077,17'd12487,17'd12488,17'd12489,17'd12489,17'd13691,17'd13691,17'd15866,17'd15866,17'd16741,17'd16741,17'd16001,17'd11330,17'd16627,17'd16136,17'd15489,17'd15489,17'd15489,17'd15489,17'd16629,17'd16629,17'd16629,17'd16857,17'd13692,17'd11195,17'd9668,17'd8655,17'd10910,17'd8810,17'd9120,17'd9120,17'd12182,17'd11879,17'd8810,17'd8503,17'd8656,17'd7533,17'd9105,17'd16858,17'd1683,17'd16859,17'd16860,17'd16861
},
'{
17'd1,17'd1,17'd12,17'd12,17'd806,17'd2933,17'd2591,17'd977,17'd4242,17'd4242,17'd2421,17'd807,17'd2591,17'd16747,17'd16636,17'd8814,17'd2421,17'd4242,17'd2933,17'd8814,17'd1128,17'd11,17'd20,17'd22,17'd5,17'd6,17'd10658,17'd16862,17'd13296,17'd16143,17'd16390,17'd12649,17'd5649,17'd16390,17'd16863,17'd16748,17'd16864,17'd8825,17'd16865,17'd3,17'd1275,17'd16747,17'd16500,17'd16749,17'd8971,17'd1127,17'd1688,17'd1688,17'd14,17'd1414,17'd31,17'd31,17'd3254,17'd2940,17'd16866,17'd2262,17'd2600,17'd1281,17'd480,17'd2439,17'd16867,17'd16868,17'd16869,17'd16870,17'd16871,17'd16753,17'd16872,17'd16873,17'd16874,17'd13446,17'd13447,17'd16155,17'd16156,17'd16875,17'd16876,17'd16877,17'd16761,17'd16878,17'd15895,17'd16654,17'd16879,17'd16656,17'd16764,17'd16764,17'd15259,17'd14098,17'd13597,17'd13968,17'd14469,17'd13092,17'd12527,17'd12813,17'd13093,17'd14621,17'd14764,17'd15764,17'd12361,17'd16765,17'd12361,17'd12361,17'd12530,17'd12530,17'd12360,17'd11627,17'd11913,17'd11362,17'd11915,17'd10945,17'd16880,17'd16034,17'd14347,17'd14346,17'd15641,17'd16030,17'd15386,17'd15260,17'd14346,17'd16881,17'd15902,17'd16882,17'd16883,17'd16884,17'd15016,17'd16773,17'd15145,17'd15268,17'd16885,17'd16886,17'd16887,17'd16888,17'd16038,17'd16889,17'd16890,17'd13105,17'd12370,17'd8703,17'd16044,17'd15402,17'd9588,17'd16891,17'd16782,17'd16892,17'd16893,17'd16894,17'd16534,17'd16670,17'd15791,17'd16537,17'd16185,17'd15279,17'd15544,17'd16895,17'd15411,17'd16896,17'd14114,17'd12077,17'd10824,17'd16897,17'd16190,17'd16898,17'd16899,17'd16787,17'd16900,17'd15414,17'd13124,17'd15420,17'd15423,17'd12567,17'd14252,17'd12842,17'd16546,17'd11934,17'd16790,17'd16901,17'd16902,17'd16903,17'd16904,17'd16905,17'd16906,17'd16907,17'd16908,17'd9341,17'd16909,17'd16910,17'd10336,17'd16911,17'd10173,17'd9344,17'd16065,17'd10742,17'd16912,17'd10476,17'd13253,17'd11960,17'd12419,17'd12420,17'd12580,17'd12109,17'd12417,17'd13517,17'd12579,17'd14807,17'd12580,17'd12420,17'd11806,17'd12996,17'd12262,17'd13362,17'd11962,17'd12857,17'd12418,17'd16913,17'd16327,17'd16327,17'd14524,17'd14524,17'd16798,17'd14672,17'd16914,17'd16915,17'd12577,17'd14810,17'd9885,17'd8881,17'd16916,17'd16917,17'd16918,17'd16919,17'd16333,17'd13765,17'd16802,17'd14531,17'd11141,17'd16920,17'd16921,17'd7626,17'd8738,17'd16922,17'd16923,17'd16924,17'd16925,17'd12433,17'd14015,17'd11976,17'd9756,17'd10873,17'd11413,17'd133,17'd1481,17'd1481,17'd133,17'd133,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd130,17'd130,17'd134,17'd132,17'd132,17'd131,17'd12127,17'd13535,17'd16926,17'd16927,17'd13016,17'd16928,17'd16929,17'd16930,17'd16931,17'd16932,17'd16706,17'd16586,17'd14703,17'd9077,17'd16820,17'd16933,17'd16934,17'd16935,17'd16936,17'd16937,17'd16938,17'd16471,17'd14555,17'd13547,17'd13547,17'd8459,17'd8764,17'd16717,17'd16716,17'd9642,17'd8762,17'd9767,17'd9223,17'd16718,17'd15085,17'd16358,17'd16826,17'd16939,17'd16828,17'd16940,17'd16941,17'd16942,17'd16943,17'd16476,17'd15326,17'd15594,17'd14038,17'd14158,17'd14292,17'd14561,17'd14415,17'd14297,17'd14714,17'd16730,17'd16729,17'd16944,17'd16945,17'd15975,17'd16477,17'd16946,17'd15211,17'd15844,17'd16947,17'd16355,17'd16355,17'd15717,17'd16729,17'd16729,17'd15844,17'd14416,17'd14294,17'd14293,17'd14292,17'd16239,17'd15330,17'd12605,17'd15331,17'd16948,17'd16605,17'd16949,17'd16244,17'd16950,17'd16951,17'd16952,17'd16840,17'd15092,17'd15221,17'd16611,17'd15986,17'd16612,17'd16246,17'd15852,17'd16843,17'd16844,17'd16845,17'd16845,17'd16370,17'd16370,17'd16953,17'd16954,17'd15473,17'd14569,17'd14570,17'd14722,17'd16121,17'd15988,17'd16247,17'd16371,17'd16955,17'd16956,17'd15610,17'd13046,17'd12162,17'd14167,17'd16617,17'd16736,17'd16957,17'd14854,17'd16851,17'd15614,17'd12907,17'd12764,17'd13804,17'd16377,17'd16958,17'd16622,17'd16491,17'd16959,17'd15735,17'd6095,17'd4729,17'd5372,17'd1272,17'd1245,17'd1382,17'd421,17'd417,17'd945,17'd15234,17'd2397,17'd2567,17'd16960,17'd5036,17'd5502,17'd7513,17'd7684,17'd8018,17'd8171,17'd9405,17'd9405,17'd10076,17'd10076,17'd10391,17'd10077,17'd12487,17'd12320,17'd13423,17'd12489,17'd13691,17'd13691,17'd15866,17'd15866,17'd16961,17'd16384,17'd16259,17'd12640,17'd16962,17'd16136,17'd15489,17'd15489,17'd15489,17'd15489,17'd16743,17'd16629,17'd16629,17'd16630,17'd13692,17'd16138,17'd10654,17'd8655,17'd10910,17'd8810,17'd9120,17'd9120,17'd12182,17'd15109,17'd8655,17'd8503,17'd10910,17'd16963,17'd16964,17'd2578,17'd639,17'd16745,17'd649,17'd16861
},
'{
17'd15,17'd14,17'd466,17'd16636,17'd8814,17'd10260,17'd4242,17'd2421,17'd2933,17'd2591,17'd977,17'd465,17'd2423,17'd16749,17'd16747,17'd2591,17'd4242,17'd4242,17'd2933,17'd8814,17'd1128,17'd11,17'd21,17'd23,17'd7,17'd5205,17'd10658,17'd16862,17'd12781,17'd16007,17'd13063,17'd5649,17'd13430,17'd16390,17'd12926,17'd16863,17'd16965,17'd15114,17'd15241,17'd283,17'd806,17'd2423,17'd16636,17'd3430,17'd466,17'd466,17'd1127,17'd1127,17'd1415,17'd1415,17'd30,17'd30,17'd3595,17'd4249,17'd2944,17'd2602,17'd16966,17'd16967,17'd994,17'd16266,17'd16968,17'd16969,17'd16970,17'd16971,17'd16972,17'd16973,17'd16974,17'd14996,17'd16975,17'd16976,17'd16977,17'd16155,17'd16978,17'd16979,17'd16980,17'd16760,17'd16651,17'd16981,17'd16982,17'd15133,17'd16983,17'd16984,17'd16985,17'd16985,17'd15259,17'd16026,17'd13839,17'd13968,17'd13092,17'd13092,17'd12527,17'd13093,17'd12065,17'd12218,17'd12530,17'd13969,17'd12361,17'd12361,17'd12530,17'd12530,17'd12530,17'd12530,17'd11627,17'd11627,17'd11764,17'd11362,17'd16766,17'd16986,17'd16519,17'd16033,17'd16168,17'd14346,17'd14892,17'd15386,17'd16290,17'd16987,17'd16411,17'd16411,17'd16028,17'd16988,17'd16989,17'd16990,17'd16991,17'd16773,17'd15145,17'd14481,17'd15909,17'd16992,17'd16993,17'd16994,17'd16995,17'd16665,17'd13104,17'd9165,17'd8703,17'd16294,17'd9588,17'd9588,17'd16996,17'd16997,17'd16533,17'd16533,17'd16183,17'd15407,17'd16535,17'd16998,17'd15923,17'd16185,17'd15279,17'd15156,17'd15281,17'd16895,17'd15032,17'd16999,17'd17000,17'd11490,17'd10709,17'd17001,17'd10446,17'd17002,17'd17003,17'd16676,17'd17004,17'd17005,17'd17006,17'd14373,17'd13995,17'd13501,17'd14799,17'd13126,17'd11934,17'd12087,17'd12088,17'd11939,17'd11652,17'd17007,17'd17008,17'd15939,17'd11664,17'd17009,17'd9477,17'd17010,17'd15567,17'd15684,17'd15807,17'd15807,17'd9345,17'd15569,17'd17011,17'd17012,17'd10329,17'd16069,17'd13363,17'd12419,17'd16321,17'd16321,17'd12580,17'd12109,17'd12109,17'd12580,17'd12580,17'd16321,17'd12420,17'd12420,17'd13135,17'd16204,17'd13362,17'd13362,17'd12114,17'd12419,17'd12859,17'd15687,17'd16560,17'd17013,17'd17014,17'd17015,17'd17014,17'd13642,17'd15571,17'd13884,17'd13363,17'd14518,17'd9346,17'd14675,17'd8104,17'd13140,17'd13649,17'd17016,17'd17017,17'd16332,17'd13377,17'd17018,17'd16568,17'd17019,17'd14013,17'd10182,17'd17020,17'd17021,17'd17022,17'd13010,17'd17023,17'd15067,17'd17024,17'd17025,17'd7812,17'd7980,17'd3025,17'd130,17'd130,17'd130,17'd133,17'd133,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd542,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd357,17'd10759,17'd5470,17'd9362,17'd17026,17'd17027,17'd17028,17'd17029,17'd17030,17'd17031,17'd17032,17'd17033,17'd17034,17'd17035,17'd17036,17'd17037,17'd17038,17'd17039,17'd17040,17'd17041,17'd16936,17'd17042,17'd16471,17'd14838,17'd13668,17'd13547,17'd13396,17'd8458,17'd9912,17'd9912,17'd8917,17'd11987,17'd9767,17'd9223,17'd11018,17'd15084,17'd16237,17'd17043,17'd17044,17'd17045,17'd17046,17'd17047,17'd17048,17'd17049,17'd16358,17'd14844,17'd14709,17'd14158,17'd14292,17'd14561,17'd14561,17'd14415,17'd14713,17'd17050,17'd17051,17'd16593,17'd16111,17'd15975,17'd15975,17'd15842,17'd17052,17'd15714,17'd16728,17'd17053,17'd17054,17'd17054,17'd15977,17'd17055,17'd16947,17'd16360,17'd16360,17'd16360,17'd16359,17'd14712,17'd14711,17'd16239,17'd17056,17'd17057,17'd17058,17'd16603,17'd16099,17'd16606,17'd16244,17'd16950,17'd17059,17'd16952,17'd17060,17'd17061,17'd17062,17'd17063,17'd16844,17'd16246,17'd16370,17'd17063,17'd17063,17'd17063,17'd16845,17'd17064,17'd16845,17'd16246,17'd16246,17'd15852,17'd15603,17'd14570,17'd14722,17'd16121,17'd15988,17'd16121,17'd17065,17'd16247,17'd17066,17'd15609,17'd12905,17'd12468,17'd14167,17'd15856,17'd14168,17'd16957,17'd15344,17'd17067,17'd17068,17'd17069,17'd17070,17'd13286,17'd17071,17'd17072,17'd14172,17'd15347,17'd16854,17'd15104,17'd4730,17'd4085,17'd5371,17'd1272,17'd952,17'd202,17'd1526,17'd198,17'd417,17'd945,17'd1384,17'd2399,17'd16000,17'd6241,17'd15350,17'd6869,17'd17073,17'd14983,17'd8018,17'd8795,17'd8795,17'd10076,17'd10076,17'd10391,17'd10391,17'd12487,17'd12487,17'd11723,17'd12489,17'd13691,17'd13691,17'd15866,17'd15866,17'd16384,17'd16383,17'd16259,17'd16001,17'd16962,17'd16627,17'd16136,17'd15489,17'd16629,17'd16629,17'd16630,17'd16629,17'd16629,17'd16630,17'd8325,17'd15870,17'd17074,17'd8655,17'd10910,17'd8810,17'd9956,17'd9956,17'd11332,17'd15109,17'd12182,17'd12492,17'd10910,17'd8657,17'd16964,17'd2578,17'd186,17'd17075,17'd16633,17'd17076
},
'{
17'd1688,17'd4247,17'd466,17'd2423,17'd2933,17'd4242,17'd4242,17'd4242,17'd2933,17'd465,17'd465,17'd2423,17'd16749,17'd16749,17'd8814,17'd977,17'd4242,17'd10260,17'd8814,17'd16747,17'd1128,17'd20,17'd23,17'd4,17'd7374,17'd8190,17'd10658,17'd17077,17'd17078,17'd16142,17'd10916,17'd5648,17'd12782,17'd12782,17'd13297,17'd12926,17'd13297,17'd7224,17'd283,17'd1275,17'd806,17'd12,17'd13,17'd3430,17'd466,17'd466,17'd2,17'd14,17'd1415,17'd1415,17'd30,17'd809,17'd3755,17'd5208,17'd2944,17'd2265,17'd1703,17'd17079,17'd1843,17'd17080,17'd17081,17'd17082,17'd17083,17'd17084,17'd16753,17'd17085,17'd17086,17'd17087,17'd17088,17'd17089,17'd17090,17'd16276,17'd17091,17'd17092,17'd17093,17'd16404,17'd17094,17'd15895,17'd17095,17'd15133,17'd16983,17'd16984,17'd16985,17'd16985,17'd15259,17'd13839,17'd13968,17'd13463,17'd13092,17'd12813,17'd12813,17'd17096,17'd12218,17'd12361,17'd12361,17'd13969,17'd12361,17'd12361,17'd12530,17'd12530,17'd12530,17'd12530,17'd11627,17'd12066,17'd11629,17'd11915,17'd16986,17'd16289,17'd15524,17'd16987,17'd14768,17'd14346,17'd14766,17'd15386,17'd16987,17'd16768,17'd16033,17'd15899,17'd17097,17'd17098,17'd17099,17'd17100,17'd16773,17'd15017,17'd17101,17'd17102,17'd16886,17'd16887,17'd17103,17'd17104,17'd16778,17'd17105,17'd9017,17'd12370,17'd7428,17'd7429,17'd9588,17'd16891,17'd16997,17'd17106,17'd17107,17'd17107,17'd16183,17'd15407,17'd16536,17'd15278,17'd17108,17'd17109,17'd16420,17'd15157,17'd15281,17'd15031,17'd16896,17'd12967,17'd17110,17'd17111,17'd17112,17'd17113,17'd17114,17'd17115,17'd17116,17'd17117,17'd17118,17'd17119,17'd12564,17'd14124,17'd14123,17'd14251,17'd12699,17'd13632,17'd12235,17'd15934,17'd11937,17'd11789,17'd11951,17'd17120,17'd11804,17'd11666,17'd17121,17'd9739,17'd17122,17'd15179,17'd16067,17'd17123,17'd15807,17'd9480,17'd11809,17'd17011,17'd17012,17'd17124,17'd11524,17'd17125,17'd13761,17'd12420,17'd16321,17'd16321,17'd12580,17'd12109,17'd12580,17'd12580,17'd12580,17'd16321,17'd12420,17'd11958,17'd12996,17'd16204,17'd13362,17'd11963,17'd12858,17'd12856,17'd16799,17'd14672,17'd16560,17'd17013,17'd16686,17'd17014,17'd17014,17'd16686,17'd15571,17'd15434,17'd11666,17'd10479,17'd8873,17'd17126,17'd7951,17'd13140,17'd15435,17'd17127,17'd17128,17'd17129,17'd13654,17'd17130,17'd17131,17'd15061,17'd17132,17'd8429,17'd17133,17'd17134,17'd17135,17'd13656,17'd11974,17'd17136,17'd17137,17'd17138,17'd11152,17'd133,17'd134,17'd130,17'd130,17'd132,17'd132,17'd133,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd357,17'd17139,17'd17140,17'd17141,17'd17142,17'd17143,17'd17144,17'd17145,17'd17146,17'd17147,17'd17148,17'd17149,17'd17150,17'd16948,17'd17151,17'd17152,17'd17153,17'd17154,17'd17155,17'd17156,17'd16936,17'd16824,17'd17157,17'd16104,17'd13548,17'd13398,17'd13668,17'd8769,17'd9642,17'd9912,17'd8917,17'd11987,17'd9767,17'd16472,17'd16473,17'd15084,17'd15213,17'd15841,17'd17158,17'd17047,17'd17159,17'd17160,17'd17161,17'd15975,17'd17162,17'd14844,17'd14709,17'd14710,17'd14561,17'd17163,17'd17163,17'd14415,17'd14159,17'd15082,17'd16834,17'd15714,17'd17164,17'd17049,17'd16597,17'd17165,17'd17166,17'd15842,17'd16111,17'd17167,17'd17167,17'd17167,17'd16944,17'd16728,17'd17055,17'd16355,17'd16835,17'd16360,17'd16360,17'd14416,17'd17168,17'd16600,17'd14562,17'd12604,17'd15596,17'd17169,17'd16603,17'd16949,17'd16606,17'd16244,17'd16608,17'd17170,17'd17060,17'd17061,17'd17062,17'd16843,17'd16843,17'd16246,17'd17171,17'd16844,17'd17063,17'd17063,17'd17064,17'd17172,17'd16845,17'd16370,17'd17171,17'd15852,17'd15723,17'd15093,17'd14570,17'd16247,17'd15988,17'd16121,17'd17065,17'd17065,17'd15725,17'd16956,17'd17173,17'd12622,17'd12468,17'd15611,17'd17174,17'd16957,17'd7671,17'd17175,17'd13170,17'd17069,17'd17176,17'd13286,17'd17071,17'd17072,17'd17177,17'd17178,17'd17179,17'd17180,17'd16492,17'd3896,17'd3895,17'd411,17'd1685,17'd1272,17'd203,17'd1669,17'd197,17'd417,17'd945,17'd2397,17'd2564,17'd6242,17'd6573,17'd6869,17'd6870,17'd7684,17'd14983,17'd8795,17'd8795,17'd10076,17'd10076,17'd9946,17'd10391,17'd11593,17'd12487,17'd11723,17'd11723,17'd13059,17'd13691,17'd15866,17'd15866,17'd16384,17'd16384,17'd17181,17'd16259,17'd17182,17'd16627,17'd16136,17'd15489,17'd16629,17'd16629,17'd16743,17'd16629,17'd16629,17'd15624,17'd17183,17'd15869,17'd17074,17'd8655,17'd10910,17'd8810,17'd9956,17'd9956,17'd11332,17'd15109,17'd12182,17'd12492,17'd11196,17'd9802,17'd17184,17'd2766,17'd1682,17'd17185,17'd1543,17'd17186
},
'{
17'd2422,17'd1831,17'd466,17'd1275,17'd2591,17'd4242,17'd4242,17'd2591,17'd465,17'd650,17'd3,17'd3430,17'd8971,17'd2423,17'd2591,17'd2591,17'd2933,17'd2933,17'd8814,17'd16747,17'd20,17'd21,17'd4,17'd6,17'd5205,17'd10658,17'd10915,17'd17077,17'd17078,17'd13296,17'd11063,17'd13062,17'd12782,17'd7059,17'd12782,17'd16390,17'd12649,17'd1413,17'd20,17'd10,17'd11,17'd18,17'd18,17'd17,17'd17,17'd17,17'd16,17'd16,17'd17187,17'd1415,17'd289,17'd4091,17'd5207,17'd5208,17'd4251,17'd2266,17'd1841,17'd2612,17'd2616,17'd17188,17'd17189,17'd17190,17'd17191,17'd17192,17'd16973,17'd16974,17'd17193,17'd14329,17'd14087,17'd13587,17'd16155,17'd17194,17'd17195,17'd17196,17'd17197,17'd17198,17'd17199,17'd17200,17'd17201,17'd15759,17'd16879,17'd16984,17'd16656,17'd16656,17'd17202,17'd17203,17'd13463,17'd13598,17'd13092,17'd13093,17'd13093,17'd13094,17'd12530,17'd13969,17'd13969,17'd12361,17'd14622,17'd14764,17'd12530,17'd12530,17'd12218,17'd12530,17'd11913,17'd11629,17'd17204,17'd17205,17'd17206,17'd17207,17'd15902,17'd16768,17'd14768,17'd14766,17'd17208,17'd17209,17'd16290,17'd16768,17'd15524,17'd16882,17'd17210,17'd17211,17'd17100,17'd15268,17'd15145,17'd17101,17'd16886,17'd16886,17'd17212,17'd16992,17'd16038,17'd17213,17'd14782,17'd14904,17'd12370,17'd16666,17'd16294,17'd15402,17'd16667,17'd17214,17'd17106,17'd17215,17'd17216,17'd16669,17'd17217,17'd16298,17'd17218,17'd15278,17'd17109,17'd17109,17'd17219,17'd15281,17'd15545,17'd15032,17'd16999,17'd17000,17'd17220,17'd10578,17'd17221,17'd17222,17'd17223,17'd16676,17'd17117,17'd16788,17'd12984,17'd16309,17'd14124,17'd13635,17'd17224,17'd14120,17'd13632,17'd17225,17'd12236,17'd12089,17'd17226,17'd17227,17'd17228,17'd17229,17'd11666,17'd13367,17'd11527,17'd10744,17'd17230,17'd8722,17'd17231,17'd14811,17'd17232,17'd15566,17'd12116,17'd10856,17'd17124,17'd10475,17'd11521,17'd14261,17'd11960,17'd16321,17'd16321,17'd12580,17'd14807,17'd14807,17'd16321,17'd16321,17'd12419,17'd12420,17'd11806,17'd13135,17'd12996,17'd16204,17'd13362,17'd13135,17'd11958,17'd12859,17'd14524,17'd14672,17'd16560,17'd17013,17'd17233,17'd17234,17'd16686,17'd17235,17'd16559,17'd15184,17'd17236,17'd11809,17'd17237,17'd10608,17'd7952,17'd17238,17'd17239,17'd17240,17'd17241,17'd14932,17'd14012,17'd12592,17'd13259,17'd16570,17'd10749,17'd14939,17'd17242,17'd17243,17'd17244,17'd12272,17'd17245,17'd17246,17'd11977,17'd10874,17'd15823,17'd132,17'd130,17'd129,17'd132,17'd132,17'd132,17'd131,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd133,17'd133,17'd133,17'd1197,17'd133,17'd135,17'd5593,17'd16579,17'd17247,17'd10192,17'd17248,17'd4981,17'd17249,17'd17250,17'd17251,17'd17252,17'd17253,17'd17254,17'd17169,17'd15833,17'd17255,17'd17256,17'd17257,17'd17258,17'd17259,17'd17041,17'd17260,17'd17042,17'd16104,17'd15973,17'd13546,17'd13546,17'd14839,17'd11832,17'd9642,17'd8917,17'd11987,17'd9767,17'd16472,17'd17261,17'd15324,17'd15325,17'd17262,17'd17263,17'd17264,17'd17265,17'd17266,17'd17267,17'd15715,17'd16238,17'd14844,17'd14710,17'd16113,17'd14561,17'd17268,17'd12445,17'd14561,17'd16599,17'd15085,17'd16594,17'd17269,17'd17049,17'd16721,17'd17270,17'd17271,17'd17272,17'd17273,17'd15974,17'd15975,17'd16945,17'd17274,17'd16832,17'd16728,17'd16728,17'd16355,17'd16355,17'd16355,17'd17275,17'd16360,17'd16360,17'd14416,17'd16601,17'd16239,17'd15980,17'd15596,17'd17169,17'd17276,17'd17277,17'd16606,17'd17278,17'd17279,17'd17279,17'd17280,17'd17281,17'd17282,17'd17283,17'd16118,17'd16370,17'd16370,17'd16246,17'd17063,17'd16844,17'd17171,17'd17171,17'd17171,17'd17171,17'd16118,17'd16118,17'd15603,17'd16119,17'd16371,17'd16121,17'd15988,17'd16247,17'd17065,17'd16247,17'd17066,17'd12761,17'd14050,17'd12468,17'd15477,17'd15991,17'd17284,17'd17285,17'd7672,17'd13170,17'd17286,17'd17287,17'd17288,17'd17289,17'd17290,17'd14057,17'd14857,17'd17291,17'd17292,17'd14858,17'd4883,17'd3391,17'd1823,17'd1111,17'd605,17'd204,17'd203,17'd421,17'd197,17'd943,17'd15234,17'd2565,17'd17293,17'd6408,17'd5502,17'd5502,17'd17073,17'd17294,17'd8491,17'd8795,17'd9405,17'd10076,17'd10076,17'd11722,17'd11593,17'd12487,17'd9110,17'd11723,17'd13059,17'd13425,17'd15866,17'd15866,17'd16384,17'd16493,17'd16135,17'd17181,17'd16626,17'd17295,17'd16136,17'd15489,17'd16629,17'd16628,17'd16629,17'd16629,17'd16743,17'd16630,17'd15624,17'd16260,17'd17296,17'd12182,17'd10910,17'd8810,17'd9956,17'd9956,17'd11332,17'd11332,17'd9120,17'd12492,17'd12493,17'd8504,17'd17297,17'd3097,17'd1682,17'd179,17'd17298,17'd649
},
'{
17'd3252,17'd1831,17'd2,17'd650,17'd977,17'd4242,17'd10260,17'd2591,17'd650,17'd1412,17'd2,17'd15745,17'd3430,17'd283,17'd651,17'd2933,17'd2933,17'd8814,17'd8814,17'd16747,17'd20,17'd21,17'd4,17'd7,17'd5205,17'd10915,17'd17077,17'd17299,17'd17078,17'd12648,17'd8510,17'd10916,17'd13063,17'd7059,17'd12782,17'd12782,17'd7375,17'd25,17'd2598,17'd20,17'd11,17'd19,17'd16,17'd16,17'd16,17'd16,17'd18,17'd18,17'd1277,17'd17187,17'd289,17'd289,17'd4091,17'd5208,17'd17300,17'd1423,17'd1285,17'd1710,17'd17301,17'd17302,17'd17303,17'd17304,17'd17305,17'd17306,17'd17307,17'd17086,17'd17308,17'd17088,17'd16274,17'd17309,17'd17310,17'd14458,17'd17311,17'd17092,17'd17312,17'd17313,17'd17314,17'd17315,17'd11472,17'd16654,17'd16879,17'd16984,17'd16656,17'd16515,17'd17316,17'd17203,17'd13463,17'd12678,17'd13093,17'd13093,17'd13094,17'd12218,17'd13969,17'd13969,17'd16658,17'd12361,17'd14764,17'd14764,17'd12530,17'd12530,17'd12218,17'd12680,17'd10815,17'd17317,17'd16766,17'd17318,17'd17319,17'd17320,17'd16033,17'd17321,17'd14892,17'd14766,17'd17208,17'd15521,17'd16290,17'd16987,17'd17322,17'd17323,17'd17324,17'd17099,17'd17325,17'd15268,17'd15145,17'd15776,17'd16037,17'd17326,17'd17327,17'd17328,17'd17329,17'd17330,17'd14904,17'd8853,17'd8703,17'd15274,17'd16044,17'd16891,17'd17214,17'd17331,17'd17332,17'd17216,17'd17333,17'd17334,17'd16534,17'd16536,17'd15408,17'd15409,17'd17109,17'd17109,17'd15410,17'd15157,17'd15031,17'd14236,17'd12967,17'd11773,17'd16052,17'd16897,17'd17113,17'd17335,17'd17336,17'd17337,17'd17338,17'd11377,17'd15420,17'd13502,17'd13355,17'd14252,17'd14922,17'd17339,17'd17340,17'd15674,17'd12088,17'd11650,17'd17341,17'd17342,17'd17008,17'd11805,17'd17343,17'd17344,17'd10169,17'd17345,17'd11402,17'd17346,17'd17347,17'd10173,17'd16549,17'd14928,17'd9739,17'd17124,17'd10475,17'd11395,17'd13646,17'd13761,17'd16321,17'd16321,17'd16321,17'd12580,17'd14807,17'd17348,17'd16321,17'd16321,17'd12420,17'd12420,17'd11806,17'd13135,17'd12996,17'd16204,17'd12996,17'd11958,17'd15570,17'd16559,17'd16915,17'd14524,17'd17013,17'd17013,17'd17233,17'd17349,17'd16560,17'd17235,17'd17350,17'd14261,17'd15176,17'd15807,17'd13002,17'd8101,17'd17351,17'd11968,17'd17352,17'd17353,17'd17354,17'd9890,17'd13528,17'd15695,17'd16806,17'd14142,17'd17355,17'd17356,17'd17357,17'd17358,17'd17359,17'd17360,17'd17361,17'd17362,17'd10874,17'd17363,17'd131,17'd134,17'd130,17'd132,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd132,17'd133,17'd133,17'd133,17'd1197,17'd133,17'd134,17'd5593,17'd11008,17'd17364,17'd17365,17'd17366,17'd17367,17'd17368,17'd17369,17'd17370,17'd17371,17'd17372,17'd17373,17'd17374,17'd17375,17'd17376,17'd17377,17'd17378,17'd17379,17'd17380,17'd17381,17'd17382,17'd16824,17'd17383,17'd16103,17'd17384,17'd17385,17'd17386,17'd8616,17'd9642,17'd16354,17'd11987,17'd9767,17'd16472,17'd17261,17'd15213,17'd15841,17'd17387,17'd17388,17'd17389,17'd17390,17'd17391,17'd17392,17'd15325,17'd16238,17'd14844,17'd17393,17'd16113,17'd14159,17'd15086,17'd14415,17'd14846,17'd16478,17'd15212,17'd17269,17'd17394,17'd17395,17'd16830,17'd17396,17'd17397,17'd17398,17'd17399,17'd17273,17'd17049,17'd17400,17'd17401,17'd17402,17'd17403,17'd16946,17'd15977,17'd16355,17'd16355,17'd16355,17'd15844,17'd16359,17'd15718,17'd15718,17'd14846,17'd14292,17'd12604,17'd15596,17'd16604,17'd17276,17'd16731,17'd17404,17'd16486,17'd17405,17'd17406,17'd17406,17'd17281,17'd17283,17'd16118,17'd16118,17'd16246,17'd16370,17'd16844,17'd16118,17'd16370,17'd17407,17'd17407,17'd17171,17'd17171,17'd16370,17'd15604,17'd15475,17'd16371,17'd16247,17'd15725,17'd15988,17'd16371,17'd16371,17'd16955,17'd16735,17'd16123,17'd14050,17'd17408,17'd15856,17'd17409,17'd17285,17'd7672,17'd17410,17'd17411,17'd12629,17'd17288,17'd17412,17'd17413,17'd14057,17'd17414,17'd17415,17'd17416,17'd17417,17'd14060,17'd3423,17'd1680,17'd1243,17'd1666,17'd425,17'd204,17'd1382,17'd1529,17'd198,17'd944,17'd2398,17'd17418,17'd6241,17'd5185,17'd5502,17'd6870,17'd17419,17'd8491,17'd8491,17'd9405,17'd10076,17'd10076,17'd12018,17'd10077,17'd12487,17'd10650,17'd9110,17'd12020,17'd13059,17'd15352,17'd15866,17'd16493,17'd16493,17'd15866,17'd17181,17'd16626,17'd17295,17'd16136,17'd15489,17'd16629,17'd16628,17'd16628,17'd16628,17'd16743,17'd16630,17'd15624,17'd17183,17'd17420,17'd11332,17'd8656,17'd8810,17'd9120,17'd9956,17'd11332,17'd11332,17'd9120,17'd12492,17'd12323,17'd8504,17'd17421,17'd9531,17'd1682,17'd17422,17'd770,17'd17423
},
'{
17'd14070,17'd1688,17'd1830,17'd650,17'd2591,17'd2933,17'd2591,17'd977,17'd283,17'd2,17'd15745,17'd15745,17'd13,17'd1275,17'd2591,17'd2591,17'd806,17'd806,17'd8814,17'd8814,17'd22,17'd23,17'd6,17'd7,17'd8190,17'd10658,17'd17424,17'd17425,17'd17299,17'd10658,17'd7727,17'd16142,17'd8520,17'd7059,17'd13063,17'd13062,17'd8,17'd23,17'd22,17'd20,17'd11,17'd18,17'd16,17'd16,17'd18,17'd18,17'd11,17'd19,17'd16,17'd16,17'd289,17'd4091,17'd5208,17'd5519,17'd2265,17'd2267,17'd993,17'd1148,17'd17426,17'd1718,17'd17427,17'd17428,17'd17429,17'd17430,17'd17431,17'd17432,17'd17433,17'd17434,17'd13587,17'd17435,17'd17436,17'd17437,17'd17438,17'd17439,17'd17440,17'd17313,17'd17441,17'd15638,17'd15133,17'd16654,17'd16879,17'd16879,17'd11624,17'd16655,17'd17442,17'd17443,17'd17444,17'd12954,17'd13093,17'd12955,17'd12218,17'd12530,17'd12361,17'd13969,17'd16658,17'd13969,17'd14764,17'd15137,17'd12218,17'd12218,17'd12680,17'd11913,17'd11629,17'd17204,17'd17205,17'd16410,17'd17445,17'd16411,17'd16987,17'd16768,17'd14892,17'd15260,17'd17209,17'd17446,17'd17447,17'd17448,17'd6299,17'd17449,17'd17450,17'd17451,17'd15145,17'd15268,17'd15776,17'd16036,17'd17326,17'd17452,17'd17453,17'd17454,17'd17455,17'd17456,17'd9017,17'd12370,17'd15537,17'd17457,17'd16996,17'd16996,17'd17331,17'd17106,17'd17216,17'd17458,17'd17333,17'd17459,17'd16670,17'd15155,17'd15409,17'd15923,17'd15279,17'd15279,17'd16185,17'd15156,17'd15032,17'd13863,17'd12968,17'd17460,17'd17461,17'd17462,17'd17222,17'd17463,17'd17464,17'd16543,17'd11377,17'd11785,17'd13503,17'd13356,17'd13635,17'd12842,17'd13873,17'd13242,17'd17225,17'd12236,17'd11937,17'd15936,17'd17465,17'd17466,17'd17467,17'd11395,17'd17468,17'd17469,17'd17470,17'd17471,17'd16553,17'd17472,17'd10174,17'd17473,17'd15566,17'd11277,17'd10164,17'd10740,17'd10737,17'd12861,17'd13761,17'd11959,17'd12419,17'd13519,17'd12106,17'd16321,17'd17348,17'd17474,17'd12106,17'd12106,17'd11960,17'd11806,17'd11962,17'd13362,17'd12422,17'd12422,17'd12996,17'd11958,17'd12418,17'd15571,17'd17475,17'd17235,17'd17235,17'd17013,17'd17476,17'd17477,17'd17013,17'd17235,17'd12253,17'd17478,17'd17479,17'd17480,17'd17481,17'd8104,17'd16566,17'd17482,17'd17483,17'd16691,17'd17484,17'd14682,17'd14678,17'd14271,17'd17485,17'd13142,17'd17486,17'd16211,17'd17487,17'd17488,17'd17489,17'd14273,17'd17490,17'd10873,17'd17363,17'd1045,17'd132,17'd132,17'd135,17'd135,17'd132,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd133,17'd133,17'd134,17'd132,17'd133,17'd134,17'd131,17'd5311,17'd3172,17'd10494,17'd17142,17'd17491,17'd17492,17'd17493,17'd17494,17'd17495,17'd17496,17'd17497,17'd17498,17'd17499,17'd17500,17'd17501,17'd17378,17'd17502,17'd17503,17'd17504,17'd17505,17'd17506,17'd17507,17'd17508,17'd17384,17'd14957,17'd12749,17'd8618,17'd17509,17'd17510,17'd9641,17'd8916,17'd11297,17'd17511,17'd15325,17'd17262,17'd16596,17'd17512,17'd17513,17'd17514,17'd17515,17'd17516,17'd15213,17'd14844,17'd14844,17'd14844,17'd16112,17'd15718,17'd14562,17'd15086,17'd14160,17'd15211,17'd15213,17'd15974,17'd17517,17'd17518,17'd17519,17'd17520,17'd17520,17'd17397,17'd17397,17'd17521,17'd17522,17'd17517,17'd17523,17'd17401,17'd17524,17'd17525,17'd17526,17'd17526,17'd17053,17'd16355,17'd16947,17'd16947,17'd15844,17'd16359,17'd15718,17'd17168,17'd14562,17'd12604,17'd15331,17'd16603,17'd17276,17'd16949,17'd17278,17'd17527,17'd17170,17'd16952,17'd17528,17'd17283,17'd16118,17'd15852,17'd16118,17'd16370,17'd16370,17'd16246,17'd16246,17'd17529,17'd17530,17'd17530,17'd17531,17'd17532,17'd15852,17'd15603,17'd16371,17'd16247,17'd16121,17'd15988,17'd17533,17'd17534,17'd16247,17'd16847,17'd17535,17'd12468,17'd17536,17'd17537,17'd16372,17'd17538,17'd7672,17'd13049,17'd17411,17'd17539,17'd13415,17'd17540,17'd17413,17'd17541,17'd17542,17'd17543,17'd17544,17'd17545,17'd17546,17'd5028,17'd624,17'd954,17'd1962,17'd1956,17'd17547,17'd1272,17'd1246,17'd420,17'd196,17'd1248,17'd2911,17'd6087,17'd5036,17'd3877,17'd5502,17'd6870,17'd14983,17'd8170,17'd8795,17'd8795,17'd10076,17'd12018,17'd10077,17'd12487,17'd10650,17'd9110,17'd11329,17'd12020,17'd15623,17'd15623,17'd15866,17'd16135,17'd16741,17'd16625,17'd16742,17'd17548,17'd16136,17'd15489,17'd16137,17'd17549,17'd17550,17'd16743,17'd16630,17'd16629,17'd14596,17'd13692,17'd16260,17'd11332,17'd10910,17'd10910,17'd9956,17'd9799,17'd9956,17'd12182,17'd9120,17'd12490,17'd8810,17'd8656,17'd8036,17'd2585,17'd17551,17'd17422,17'd15492,17'd17552
},
'{
17'd3252,17'd1689,17'd3749,17'd650,17'd465,17'd1275,17'd465,17'd465,17'd1,17'd466,17'd2594,17'd4247,17'd2,17'd283,17'd465,17'd2591,17'd806,17'd806,17'd8814,17'd8814,17'd22,17'd4,17'd6,17'd7,17'd10537,17'd10537,17'd17424,17'd17425,17'd10915,17'd10537,17'd12648,17'd12781,17'd12649,17'd13063,17'd10916,17'd5514,17'd4,17'd22,17'd22,17'd20,17'd11,17'd19,17'd16,17'd16,17'd18,17'd18,17'd11,17'd11,17'd18,17'd16,17'd289,17'd289,17'd3433,17'd4251,17'd1422,17'd17553,17'd17554,17'd17555,17'd1715,17'd17556,17'd17557,17'd17558,17'd17559,17'd17560,17'd17561,17'd17562,17'd16646,17'd17563,17'd16154,17'd15635,17'd17564,17'd17437,17'd17565,17'd14612,17'd17566,17'd17567,17'd17568,17'd15758,17'd17569,17'd17570,17'd16879,17'd16879,17'd16763,17'd16025,17'd17571,17'd17444,17'd12954,17'd12813,17'd12955,17'd12955,17'd12218,17'd12530,17'd13969,17'd13969,17'd16658,17'd13969,17'd14764,17'd15137,17'd12218,17'd12218,17'd12680,17'd10815,17'd17204,17'd16766,17'd17572,17'd17207,17'd15902,17'd16290,17'd16987,17'd17321,17'd14893,17'd15521,17'd17573,17'd17574,17'd17575,17'd5833,17'd17576,17'd17577,17'd16990,17'd16525,17'd15017,17'd17101,17'd15776,17'd15776,17'd16887,17'd16887,17'd17578,17'd17579,17'd17580,17'd14782,17'd9165,17'd16666,17'd17581,17'd17582,17'd16996,17'd17583,17'd17106,17'd17584,17'd17458,17'd17333,17'd17585,17'd17586,17'd17587,17'd15922,17'd15923,17'd15923,17'd15279,17'd16420,17'd15279,17'd17588,17'd16896,17'd17589,17'd11925,17'd17590,17'd17591,17'd17592,17'd17335,17'd17336,17'd10448,17'd15039,17'd12561,17'd17593,17'd12400,17'd13356,17'd15673,17'd12842,17'd14661,17'd11934,17'd12560,17'd12237,17'd17594,17'd17595,17'd17596,17'd17597,17'd17598,17'd12862,17'd17599,17'd15295,17'd17600,17'd10174,17'd16795,17'd15807,17'd17601,17'd15566,17'd12116,17'd11134,17'd10740,17'd10853,17'd12262,17'd11806,17'd11960,17'd16321,17'd13365,17'd13136,17'd12106,17'd12106,17'd17474,17'd17602,17'd17603,17'd12106,17'd13883,17'd11806,17'd11963,17'd12262,17'd17604,17'd12422,17'd15053,17'd16321,17'd14930,17'd15571,17'd17475,17'd17235,17'd17235,17'd17235,17'd17013,17'd16914,17'd17013,17'd17605,17'd15184,17'd12583,17'd17606,17'd17607,17'd8248,17'd7949,17'd17608,17'd14676,17'd8251,17'd17609,17'd16447,17'd14391,17'd10997,17'd14013,17'd17610,17'd14394,17'd17020,17'd17611,17'd17612,17'd17613,17'd17614,17'd17615,17'd17616,17'd13777,17'd133,17'd11541,17'd132,17'd132,17'd135,17'd132,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd132,17'd132,17'd132,17'd133,17'd134,17'd132,17'd133,17'd134,17'd131,17'd3811,17'd17617,17'd17618,17'd6201,17'd17619,17'd17620,17'd17621,17'd17622,17'd17623,17'd17624,17'd17625,17'd17626,17'd17627,17'd17628,17'd17629,17'd17630,17'd17631,17'd17632,17'd17633,17'd17634,17'd17635,17'd17636,17'd16470,17'd17637,17'd14957,17'd13399,17'd17638,17'd17639,17'd17640,17'd17510,17'd8917,17'd17641,17'd17162,17'd15325,17'd17044,17'd17642,17'd17643,17'd17644,17'd17645,17'd17515,17'd17516,17'd15714,17'd16599,17'd14844,17'd16599,17'd16112,17'd15718,17'd14562,17'd14562,17'd16478,17'd15212,17'd15842,17'd17646,17'd17518,17'd17647,17'd16942,17'd17045,17'd17648,17'd17648,17'd17397,17'd17397,17'd17521,17'd17522,17'd17649,17'd17517,17'd17650,17'd17524,17'd16832,17'd16727,17'd16944,17'd17053,17'd17053,17'd16947,17'd16947,17'd15844,17'd16725,17'd15718,17'd14846,17'd14562,17'd12604,17'd17651,17'd16586,17'd17652,17'd16606,17'd15983,17'd17527,17'd17170,17'd17528,17'd15093,17'd15724,17'd16118,17'd16118,17'd16246,17'd16370,17'd16370,17'd16953,17'd17529,17'd17530,17'd17531,17'd17653,17'd17530,17'd16246,17'd15723,17'd16371,17'd16247,17'd16121,17'd16121,17'd17533,17'd17654,17'd16371,17'd15606,17'd17655,17'd14423,17'd17656,17'd15611,17'd16372,17'd17657,17'd17175,17'd17410,17'd12628,17'd17288,17'd13415,17'd17540,17'd17413,17'd17658,17'd14173,17'd17659,17'd17291,17'd16854,17'd17660,17'd12483,17'd5629,17'd623,17'd626,17'd7512,17'd17661,17'd425,17'd952,17'd1382,17'd415,17'd418,17'd1386,17'd3228,17'd5503,17'd5036,17'd5502,17'd6869,17'd14983,17'd8170,17'd8795,17'd8795,17'd10076,17'd12018,17'd10077,17'd12019,17'd10650,17'd10650,17'd11051,17'd12020,17'd15623,17'd15623,17'd15866,17'd16135,17'd16741,17'd16625,17'd16742,17'd17548,17'd16627,17'd16136,17'd16137,17'd17549,17'd17550,17'd16743,17'd16630,17'd16629,17'd14596,17'd8325,17'd16260,17'd13939,17'd10910,17'd10910,17'd9120,17'd10256,17'd11332,17'd12182,17'd9120,17'd12642,17'd12493,17'd10910,17'd8036,17'd2774,17'd610,17'd1826,17'd402,17'd17185
},
'{
17'd4247,17'd15,17'd4884,17'd1412,17'd283,17'd1275,17'd1275,17'd3,17'd466,17'd4247,17'd4247,17'd466,17'd12,17'd1275,17'd2591,17'd2933,17'd806,17'd2423,17'd16747,17'd8814,17'd23,17'd6,17'd5205,17'd5205,17'd10795,17'd8340,17'd17662,17'd17663,17'd10913,17'd17664,17'd17665,17'd10796,17'd12925,17'd12925,17'd13062,17'd8,17'd22,17'd22,17'd22,17'd21,17'd11,17'd11,17'd19,17'd19,17'd11,17'd11,17'd20,17'd11,17'd19,17'd16,17'd289,17'd3595,17'd4249,17'd2265,17'd1136,17'd2788,17'd671,17'd17666,17'd17667,17'd17668,17'd17669,17'd17670,17'd17671,17'd17672,17'd17673,17'd17674,17'd17675,17'd17676,17'd17677,17'd17678,17'd17679,17'd17437,17'd16979,17'd17566,17'd17680,17'd17681,17'd17682,17'd15638,17'd17683,17'd17684,17'd17683,17'd16514,17'd17685,17'd16405,17'd17686,17'd17687,17'd17688,17'd17096,17'd13211,17'd12218,17'd12218,17'd12530,17'd13969,17'd13969,17'd15764,17'd14622,17'd14764,17'd14890,17'd12218,17'd13094,17'd12680,17'd11629,17'd17689,17'd16986,17'd17319,17'd17690,17'd16033,17'd16165,17'd16987,17'd17691,17'd17208,17'd15521,17'd17692,17'd17693,17'd17694,17'd17695,17'd17696,17'd17697,17'd16525,17'd15017,17'd17698,17'd17698,17'd16992,17'd17326,17'd16887,17'd16663,17'd17699,17'd17700,17'd17701,17'd15783,17'd12370,17'd8703,17'd17457,17'd17582,17'd17214,17'd16997,17'd17702,17'd17702,17'd17333,17'd17333,17'd17586,17'd17703,17'd17704,17'd15923,17'd17108,17'd15923,17'd16420,17'd17705,17'd17706,17'd14361,17'd12966,17'd17707,17'd17708,17'd10709,17'd17709,17'd17710,17'd16786,17'd17711,17'd15932,17'd11109,17'd12087,17'd14125,17'd13503,17'd17712,17'd12842,17'd14661,17'd12235,17'd16790,17'd12240,17'd11788,17'd17713,17'd17714,17'd12104,17'd12112,17'd11520,17'd17715,17'd9345,17'd16910,17'd8720,17'd17716,17'd15807,17'd17717,17'd17718,17'd10024,17'd17719,17'd17720,17'd16320,17'd14262,17'd12996,17'd11958,17'd16321,17'd16321,17'd13365,17'd13136,17'd12106,17'd12106,17'd17602,17'd17721,17'd17722,17'd13883,17'd11806,17'd13135,17'd13362,17'd12115,17'd12261,17'd17723,17'd12719,17'd13517,17'd16914,17'd17724,17'd17725,17'd17726,17'd17727,17'd17235,17'd17013,17'd16914,17'd17013,17'd13884,17'd13646,17'd12423,17'd17728,17'd17729,17'd9888,17'd17609,17'd9197,17'd17017,17'd17730,17'd7952,17'd16078,17'd17731,17'd8738,17'd7464,17'd15308,17'd17732,17'd17733,17'd17734,17'd17735,17'd13532,17'd17736,17'd17737,17'd13899,17'd131,17'd131,17'd134,17'd132,17'd132,17'd135,17'd132,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd134,17'd132,17'd3168,17'd12734,17'd7485,17'd17738,17'd17739,17'd17740,17'd17741,17'd17742,17'd17743,17'd17744,17'd17745,17'd17746,17'd17747,17'd17748,17'd17749,17'd17750,17'd17751,17'd17752,17'd17753,17'd17754,17'd17755,17'd17756,17'd17757,17'd17758,17'd12749,17'd8922,17'd13399,17'd8616,17'd11694,17'd10202,17'd9642,17'd16718,17'd17162,17'd15841,17'd17759,17'd17760,17'd17761,17'd17762,17'd17763,17'd17764,17'd17516,17'd16477,17'd17765,17'd15326,17'd14960,17'd16112,17'd15718,17'd14562,17'd15718,17'd15211,17'd15715,17'd17766,17'd17767,17'd17768,17'd17769,17'd17770,17'd16942,17'd17396,17'd17396,17'd16940,17'd17396,17'd16830,17'd17771,17'd17518,17'd17772,17'd17766,17'd17773,17'd17274,17'd16832,17'd16832,17'd16727,17'd16727,17'd16726,17'd17053,17'd15717,17'd15844,17'd16360,17'd14416,17'd16600,17'd14562,17'd12604,17'd12887,17'd16604,17'd17774,17'd16484,17'd17775,17'd17776,17'd17777,17'd16841,17'd15724,17'd17283,17'd16118,17'd16246,17'd16370,17'd17171,17'd17532,17'd17529,17'd17531,17'd17778,17'd17778,17'd17653,17'd17171,17'd15852,17'd17779,17'd16247,17'd16247,17'd16247,17'd15337,17'd15475,17'd17779,17'd16121,17'd15340,17'd14423,17'd17780,17'd15611,17'd15991,17'd14426,17'd17781,17'd16739,17'd17782,17'd13566,17'd17289,17'd13567,17'd17072,17'd17658,17'd17783,17'd14857,17'd17784,17'd17291,17'd17785,17'd13056,17'd17786,17'd1402,17'd2587,17'd233,17'd17787,17'd207,17'd644,17'd1685,17'd422,17'd194,17'd1106,17'd3080,17'd3398,17'd3877,17'd5366,17'd5502,17'd17419,17'd9945,17'd8795,17'd9253,17'd10076,17'd12018,17'd10077,17'd10077,17'd10650,17'd9110,17'd11329,17'd12020,17'd15238,17'd15623,17'd15866,17'd15866,17'd16741,17'd16625,17'd16742,17'd16626,17'd16627,17'd16136,17'd17549,17'd17549,17'd17550,17'd16629,17'd16630,17'd16629,17'd15624,17'd8325,17'd16260,17'd17788,17'd10910,17'd10910,17'd9120,17'd9799,17'd9956,17'd11332,17'd9120,17'd12490,17'd8810,17'd11196,17'd16495,17'd2774,17'd188,17'd17789,17'd402,17'd1826
},
'{
17'd466,17'd1412,17'd4884,17'd1412,17'd1,17'd1412,17'd1,17'd2,17'd2594,17'd2594,17'd4247,17'd2,17'd283,17'd465,17'd2933,17'd8814,17'd806,17'd2423,17'd16747,17'd2933,17'd4,17'd6,17'd5205,17'd5205,17'd10795,17'd10795,17'd17790,17'd17664,17'd10912,17'd17790,17'd17665,17'd10796,17'd12781,17'd13062,17'd7216,17'd23,17'd5518,17'd22,17'd22,17'd21,17'd20,17'd11,17'd11,17'd11,17'd11,17'd11,17'd20,17'd11,17'd19,17'd29,17'd289,17'd3595,17'd3105,17'd1840,17'd17553,17'd17791,17'd17792,17'd17793,17'd17794,17'd17795,17'd17796,17'd17797,17'd17798,17'd17799,17'd17800,17'd17674,17'd17675,17'd17801,17'd17802,17'd15255,17'd17803,17'd17804,17'd14883,17'd14612,17'd17805,17'd17806,17'd17807,17'd17200,17'd17201,17'd11355,17'd17683,17'd16514,17'd16405,17'd16162,17'd17808,17'd17687,17'd17809,17'd17096,17'd13094,17'd12218,17'd12530,17'd13840,17'd13969,17'd13969,17'd14622,17'd14764,17'd15137,17'd12814,17'd13094,17'd12957,17'd10815,17'd17317,17'd16986,17'd16289,17'd16519,17'd17810,17'd16987,17'd16290,17'd17811,17'd17208,17'd15643,17'd16165,17'd17447,17'd17448,17'd17812,17'd17813,17'd17814,17'd17815,17'd16525,17'd15017,17'd14481,17'd15776,17'd17326,17'd17326,17'd16775,17'd16529,17'd17816,17'd17817,17'd17105,17'd17818,17'd12071,17'd7428,17'd17457,17'd17214,17'd16997,17'd17819,17'd17702,17'd17820,17'd17821,17'd17822,17'd17703,17'd17823,17'd17824,17'd17824,17'd17108,17'd15923,17'd16420,17'd17705,17'd14361,17'd17825,17'd17826,17'd17827,17'd17828,17'd17829,17'd17830,17'd10139,17'd16899,17'd17337,17'd13629,17'd11786,17'd13504,17'd13504,17'd13502,17'd15169,17'd14661,17'd17831,17'd17832,17'd17833,17'd17834,17'd17835,17'd11508,17'd17836,17'd17837,17'd13366,17'd17838,17'd17839,17'd17840,17'd9038,17'd9039,17'd10174,17'd10334,17'd17841,17'd13522,17'd17842,17'd10326,17'd10740,17'd10737,17'd11963,17'd12719,17'd12106,17'd16321,17'd16321,17'd13136,17'd13136,17'd12106,17'd17603,17'd17721,17'd17721,17'd17722,17'd13883,17'd13135,17'd12996,17'd12262,17'd12115,17'd12261,17'd17843,17'd12106,17'd12417,17'd16560,17'd17844,17'd17845,17'd17846,17'd17727,17'd17727,17'd17235,17'd15687,17'd14672,17'd12414,17'd16068,17'd17847,17'd17848,17'd11967,17'd17849,17'd17850,17'd9197,17'd16333,17'd7785,17'd17851,17'd17852,17'd17853,17'd14393,17'd9893,17'd17854,17'd17855,17'd17856,17'd17857,17'd17858,17'd17859,17'd17860,17'd17861,17'd16090,17'd131,17'd132,17'd132,17'd132,17'd132,17'd135,17'd132,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd132,17'd132,17'd132,17'd134,17'd131,17'd15579,17'd4168,17'd17862,17'd17863,17'd17864,17'd17865,17'd17866,17'd17867,17'd17868,17'd17869,17'd17870,17'd17871,17'd17379,17'd17872,17'd17873,17'd17874,17'd17875,17'd17876,17'd17877,17'd17878,17'd17879,17'd17756,17'd17880,17'd13274,17'd17638,17'd17638,17'd8767,17'd11832,17'd10202,17'd9912,17'd17881,17'd15084,17'd17262,17'd17882,17'd17883,17'd17884,17'd17885,17'd17886,17'd17887,17'd17516,17'd15841,17'd17765,17'd14961,17'd14960,17'd16112,17'd15718,17'd15718,17'd15593,17'd15976,17'd15974,17'd17521,17'd16830,17'd17769,17'd17769,17'd17888,17'd17770,17'd16942,17'd17889,17'd17396,17'd17396,17'd17768,17'd17768,17'd16829,17'd17890,17'd17395,17'd17891,17'd17892,17'd17773,17'd16110,17'd16236,17'd16236,17'd16727,17'd16944,17'd15977,17'd17893,17'd17894,17'd17894,17'd15718,17'd14293,17'd14561,17'd12604,17'd12743,17'd17895,17'd17896,17'd17897,17'd17898,17'd17899,17'd17900,17'd17901,17'd15605,17'd15852,17'd15852,17'd16246,17'd17171,17'd17529,17'd17532,17'd17530,17'd17902,17'd17778,17'd17778,17'd17407,17'd16246,17'd17903,17'd16371,17'd16247,17'd16371,17'd15337,17'd15336,17'd17903,17'd17065,17'd17904,17'd15094,17'd17905,17'd17408,17'd17537,17'd15343,17'd17906,17'd16739,17'd13565,17'd17907,17'd17289,17'd13567,17'd17908,17'd17909,17'd17910,17'd17542,17'd17911,17'd17912,17'd17913,17'd13055,17'd17914,17'd4398,17'd628,17'd1546,17'd17915,17'd1097,17'd207,17'd803,17'd603,17'd2763,17'd948,17'd1387,17'd3399,17'd3877,17'd5366,17'd5366,17'd17073,17'd17916,17'd8795,17'd9253,17'd9405,17'd10076,17'd13690,17'd10077,17'd10650,17'd10650,17'd11051,17'd11329,17'd15238,17'd15238,17'd15866,17'd15866,17'd16741,17'd16625,17'd16742,17'd16626,17'd16627,17'd16136,17'd17549,17'd17549,17'd17550,17'd16629,17'd16630,17'd16629,17'd15624,17'd14596,17'd17183,17'd17296,17'd10910,17'd8656,17'd12322,17'd10256,17'd11332,17'd12182,17'd9120,17'd12642,17'd11196,17'd11196,17'd16495,17'd5192,17'd2112,17'd254,17'd934,17'd639
},
'{
17'd13,17'd283,17'd650,17'd1,17'd0,17'd1830,17'd15,17'd4247,17'd17917,17'd2594,17'd466,17'd0,17'd283,17'd465,17'd2933,17'd16747,17'd2423,17'd2423,17'd8814,17'd10260,17'd5,17'd7,17'd5205,17'd8040,17'd10912,17'd17790,17'd17664,17'd10912,17'd10913,17'd17790,17'd17662,17'd17918,17'd12648,17'd7216,17'd8,17'd22,17'd21,17'd21,17'd21,17'd21,17'd20,17'd20,17'd26,17'd26,17'd26,17'd26,17'd27,17'd27,17'd28,17'd4431,17'd3755,17'd3434,17'd2945,17'd17919,17'd2788,17'd671,17'd17920,17'd1571,17'd17921,17'd17922,17'd16971,17'd17923,17'd17924,17'd17925,17'd17926,17'd17674,17'd17675,17'd17927,17'd17928,17'd17929,17'd17930,17'd15000,17'd17931,17'd14090,17'd17932,17'd17681,17'd17933,17'd17200,17'd17201,17'd17934,17'd17569,17'd16762,17'd17935,17'd17936,17'd17937,17'd17938,17'd17939,17'd17940,17'd12218,17'd12530,17'd12530,17'd13840,17'd14891,17'd14764,17'd14764,17'd14621,17'd12814,17'd12814,17'd12218,17'd12680,17'd10815,17'd17941,17'd17206,17'd17319,17'd17320,17'd16033,17'd16290,17'd16987,17'd16987,17'd16165,17'd15769,17'd17321,17'd17942,17'd6132,17'd17943,17'd17577,17'd17944,17'd14631,17'd16773,17'd17325,17'd16036,17'd15776,17'd15392,17'd16530,17'd16177,17'd16995,17'd14639,17'd17105,17'd17818,17'd12370,17'd11920,17'd9313,17'd17583,17'd16997,17'd17945,17'd17946,17'd17947,17'd17820,17'd17948,17'd17949,17'd17950,17'd17704,17'd17824,17'd17951,17'd17952,17'd15409,17'd15279,17'd17705,17'd13738,17'd12546,17'd17953,17'd17954,17'd17955,17'd17956,17'd17957,17'd17002,17'd17958,17'd17338,17'd12395,17'd12568,17'd17959,17'd12709,17'd14372,17'd16308,17'd15420,17'd12560,17'd17833,17'd11940,17'd17960,17'd11383,17'd17961,17'd12409,17'd15679,17'd16068,17'd10478,17'd17962,17'd17840,17'd17963,17'd17964,17'd12117,17'd17965,17'd13522,17'd13369,17'd17966,17'd16320,17'd10853,17'd10989,17'd12996,17'd16321,17'd14807,17'd16321,17'd12106,17'd13519,17'd12259,17'd12719,17'd12581,17'd17967,17'd17967,17'd15053,17'd13883,17'd13135,17'd13362,17'd12115,17'd17968,17'd12261,17'd12581,17'd14807,17'd12415,17'd17476,17'd17969,17'd17970,17'd17971,17'd17727,17'd17727,17'd15571,17'd14524,17'd12997,17'd13363,17'd10476,17'd9479,17'd8885,17'd14812,17'd8252,17'd17128,17'd17016,17'd9197,17'd17972,17'd9623,17'd17019,17'd17356,17'd17856,17'd17973,17'd17974,17'd17975,17'd17976,17'd17977,17'd17978,17'd11976,17'd17490,17'd12275,17'd16090,17'd131,17'd134,17'd132,17'd133,17'd133,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd134,17'd131,17'd3812,17'd17979,17'd17980,17'd17981,17'd17982,17'd17983,17'd17984,17'd17985,17'd17986,17'd17987,17'd17988,17'd17989,17'd17989,17'd17990,17'd17991,17'd17992,17'd17993,17'd17994,17'd17995,17'd17996,17'd17748,17'd17997,17'd17998,17'd17999,17'd18000,17'd9772,17'd8618,17'd18001,17'd8917,17'd11162,17'd17261,17'd15713,17'd16939,17'd16831,17'd18002,17'd18003,17'd18004,17'd18005,17'd17887,17'd17392,17'd16939,17'd15083,17'd14961,17'd14961,17'd16112,17'd15718,17'd14294,17'd15717,17'd16110,17'd17646,17'd17396,17'd17888,17'd18006,17'd18006,17'd18006,17'd17888,17'd18007,17'd18008,17'd18007,17'd18007,17'd18009,17'd18010,17'd17768,17'd18011,17'd17890,17'd18012,17'd18013,17'd18014,17'd17892,17'd17773,17'd16110,17'd16236,17'd15715,17'd15976,17'd18015,17'd15717,17'd15717,17'd16359,17'd16362,17'd16113,17'd14710,17'd14158,17'd18016,17'd17150,17'd18017,17'd18018,17'd16486,17'd17059,17'd17281,17'd17281,17'd17282,17'd17283,17'd17063,17'd16845,17'd16370,17'd16246,17'd18019,17'd18020,17'd17778,17'd17778,17'd18020,17'd17171,17'd18021,17'd17654,17'd16119,17'd16119,17'd15337,17'd15337,17'd17534,17'd17779,17'd18022,17'd15340,17'd18023,17'd17780,17'd17537,17'd18024,17'd18025,17'd18026,17'd13565,17'd18027,17'd17289,17'd13567,17'd18028,17'd18029,17'd18030,17'd14173,17'd18031,17'd17784,17'd18032,17'd18033,17'd18034,17'd18035,17'd3874,17'd235,17'd1093,17'd2255,17'd459,17'd272,17'd1098,17'd2117,17'd13573,17'd1252,17'd3400,17'd3877,17'd5502,17'd5366,17'd7028,17'd17294,17'd11191,17'd11191,17'd8795,17'd10076,17'd13690,17'd10077,17'd12487,17'd10650,17'd11051,17'd11329,17'd12918,17'd15238,17'd15866,17'd15866,17'd16741,17'd16625,17'd16742,17'd16626,17'd16962,17'd16627,17'd17549,17'd17549,17'd16628,17'd16629,17'd16630,17'd16743,17'd16743,17'd16857,17'd14596,17'd16138,17'd14985,17'd15739,17'd8810,17'd9800,17'd11332,17'd12182,17'd8330,17'd14866,17'd5186,17'd9121,17'd16495,17'd3742,17'd2112,17'd460,17'd1403,17'd965
},
'{
17'd2423,17'd806,17'd3,17'd0,17'd14,17'd3249,17'd1689,17'd1831,17'd17917,17'd4247,17'd2,17'd3,17'd465,17'd1275,17'd8814,17'd2423,17'd12,17'd12,17'd1275,17'd2421,17'd6,17'd5205,17'd8040,17'd8340,17'd18036,17'd17790,17'd10913,17'd18036,17'd17664,17'd17790,17'd17790,17'd17918,17'd7374,17'd5206,17'd4,17'd23,17'd21,17'd21,17'd21,17'd21,17'd21,17'd21,17'd285,17'd285,17'd285,17'd26,17'd27,17'd28,17'd18037,17'd4431,17'd5208,17'd4250,17'd2606,17'd1284,17'd18038,17'd18039,17'd18040,17'd18041,17'd18042,17'd17669,17'd18043,17'd18044,17'd18045,17'd18046,17'd18047,17'd18048,17'd17675,17'd18049,17'd18050,17'd18051,17'd18052,17'd15507,17'd18053,17'd16979,17'd14333,17'd17440,17'd18054,17'd17315,17'd15257,17'd18055,17'd17201,17'd18056,17'd18057,17'd17937,17'd18058,17'd17939,17'd17940,17'd14470,17'd12530,17'd12530,17'd13840,17'd13840,17'd14891,17'd14764,17'd14621,17'd13211,17'd12814,17'd12218,17'd12680,17'd12531,17'd17204,17'd17205,17'd17319,17'd17320,17'd16411,17'd16033,17'd16987,17'd16290,17'd16290,17'd16165,17'd16290,17'd18059,17'd18060,17'd18061,17'd18062,17'd17577,17'd16990,17'd16526,17'd15017,17'd18063,17'd15776,17'd17326,17'd16530,17'd16178,17'd15781,17'd15272,17'd17456,17'd13104,17'd9165,17'd12071,17'd11920,17'd9313,17'd18064,17'd17819,17'd17946,17'd17946,17'd17702,17'd17702,17'd18065,17'd18066,17'd18067,17'd18068,17'd18069,17'd17951,17'd17952,17'd15409,17'd15279,17'd14909,17'd13488,17'd18070,17'd11101,17'd18071,17'd16539,17'd18072,17'd18073,17'd17115,17'd18074,17'd16195,17'd11936,17'd13637,17'd15671,17'd12567,17'd14372,17'd11934,17'd17593,17'd11936,17'd12850,17'd11790,17'd18075,17'd12991,17'd18076,17'd18077,17'd18078,17'd13886,17'd11136,17'd18079,17'd9344,17'd9344,17'd15180,17'd18080,17'd9741,17'd13522,17'd17966,17'd11398,17'd16068,17'd14262,17'd12262,17'd13135,17'd12580,17'd14807,17'd16321,17'd11958,17'd14002,17'd18081,17'd12581,17'd17843,17'd17967,17'd17603,17'd15053,17'd15053,17'd12996,17'd12262,17'd12115,17'd18082,17'd12421,17'd12106,17'd12254,17'd12860,17'd17969,17'd17969,17'd17475,17'd17727,17'd18083,17'd18084,17'd16558,17'd16559,17'd12413,17'd11666,17'd10479,17'd10335,17'd8412,17'd12426,17'd16691,17'd17850,17'd15056,17'd10860,17'd18085,17'd18086,17'd18087,17'd18088,17'd18089,17'd18090,17'd18091,17'd18092,17'd18093,17'd18094,17'd17859,17'd17860,17'd15821,17'd7980,17'd133,17'd11541,17'd134,17'd132,17'd133,17'd133,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd134,17'd132,17'd135,17'd132,17'd132,17'd132,17'd5311,17'd18095,17'd18096,17'd15314,17'd18097,17'd18098,17'd18099,17'd18100,17'd18101,17'd18102,17'd18103,17'd18104,17'd18105,17'd18105,17'd18106,17'd18107,17'd18108,17'd18109,17'd18110,17'd18111,17'd18112,17'd17879,17'd10051,17'd12892,17'd18000,17'd9772,17'd8767,17'd8616,17'd16354,17'd9374,17'd10768,17'd15713,17'd17387,17'd18113,17'd18114,17'd18115,17'd18116,17'd18117,17'd18118,17'd17392,17'd16596,17'd16594,17'd15085,17'd14961,17'd16112,17'd14294,17'd16359,17'd18015,17'd17891,17'd17767,17'd18119,17'd18120,17'd18121,17'd18121,17'd18122,17'd16941,17'd18123,17'd18124,17'd18123,17'd18123,17'd16941,17'd18009,17'd18125,17'd16829,17'd18126,17'd17890,17'd17890,17'd18127,17'd18013,17'd17891,17'd17766,17'd16110,17'd15842,17'd15715,17'd16944,17'd15716,17'd15716,17'd18128,17'd18128,17'd16362,17'd14293,17'd14710,17'd15329,17'd18129,17'd17895,17'd18017,17'd18130,17'd17527,17'd16952,17'd17062,17'd17281,17'd17282,17'd16843,17'd17063,17'd16246,17'd16246,17'd17171,17'd17407,17'd17653,17'd17778,17'd18020,17'd17407,17'd18131,17'd18132,17'd15475,17'd16119,17'd15337,17'd15337,17'd18133,17'd17534,17'd18134,17'd17904,17'd18135,17'd17905,17'd17656,17'd18024,17'd15859,17'd18136,17'd13565,17'd16621,17'd17289,17'd17412,17'd16853,17'd18137,17'd18138,17'd14308,17'd18139,17'd17911,17'd14433,17'd18140,17'd18141,17'd18142,17'd18143,17'd18144,17'd633,17'd1682,17'd965,17'd257,17'd645,17'd1686,17'd950,17'd18145,17'd3401,17'd3877,17'd5502,17'd5366,17'd5501,17'd17419,17'd11444,17'd11191,17'd8795,17'd9253,17'd13690,17'd13935,17'd12019,17'd12487,17'd11723,17'd11051,17'd18146,17'd15238,17'd16135,17'd15866,17'd16741,17'd16741,17'd18147,17'd16742,17'd17182,17'd16962,17'd18148,17'd17549,17'd16629,17'd16629,17'd16630,17'd16743,17'd16743,17'd16857,17'd14596,17'd15870,17'd15110,17'd13294,17'd8503,17'd7034,17'd12182,17'd12182,17'd8330,17'd9801,17'd18149,17'd13294,17'd9669,17'd2392,17'd1678,17'd2588,17'd965,17'd804
},
'{
17'd16499,17'd16747,17'd16636,17'd2,17'd14,17'd1689,17'd1688,17'd1831,17'd2594,17'd1127,17'd0,17'd283,17'd465,17'd2933,17'd8814,17'd16747,17'd16636,17'd806,17'd2591,17'd978,17'd6,17'd5205,17'd8040,17'd8340,17'd10912,17'd10913,17'd10912,17'd10912,17'd10913,17'd17664,17'd17664,17'd17664,17'd5205,17'd6,17'd4,17'd23,17'd21,17'd21,17'd21,17'd21,17'd22,17'd22,17'd1832,17'd1832,17'd285,17'd285,17'd27,17'd27,17'd6744,17'd5971,17'd5655,17'd4251,17'd1422,17'd18150,17'd18151,17'd18152,17'd18153,17'd18154,17'd18155,17'd18156,17'd18157,17'd18158,17'd18159,17'd18160,17'd18161,17'd18048,17'd18162,17'd18163,17'd18164,17'd14202,17'd18165,17'd15507,17'd16401,17'd13963,17'd18166,17'd18167,17'd18054,17'd17315,17'd15638,17'd15513,17'd16982,17'd18168,17'd18169,17'd18170,17'd18171,17'd18172,17'd18173,17'd14470,17'd12361,17'd13969,17'd13840,17'd13840,17'd14891,17'd14764,17'd13211,17'd13211,17'd13094,17'd12218,17'd12680,17'd12532,17'd17941,17'd18174,17'd17207,17'd17445,17'd16033,17'd16987,17'd16987,17'd16165,17'd16165,17'd16987,17'd18175,17'd17448,17'd17097,17'd14223,17'd18176,17'd17211,17'd14631,17'd15016,17'd18063,17'd18063,17'd17212,17'd17326,17'd16178,17'd16040,17'd18177,17'd18178,17'd18179,17'd12822,17'd12370,17'd8703,17'd10701,17'd9708,17'd9708,17'd9708,17'd18180,17'd18180,17'd17946,17'd17458,17'd17949,17'd18067,17'd18068,17'd18069,17'd17951,17'd18181,17'd17952,17'd15409,17'd15791,17'd14786,17'd18182,17'd18183,17'd18184,17'd10578,17'd18185,17'd18186,17'd18187,17'd18188,17'd13992,17'd13237,17'd13637,17'd18189,17'd13995,17'd12986,17'd14513,17'd12559,17'd12087,17'd12241,17'd13876,17'd13248,17'd18190,17'd18191,17'd18192,17'd12110,17'd11519,17'd10741,17'd18193,17'd9339,17'd9885,17'd13255,17'd18194,17'd18195,17'd18196,17'd10330,17'd11668,17'd11396,17'd13762,17'd12262,17'd12114,17'd12857,17'd12110,17'd12580,17'd12106,17'd12719,17'd18081,17'd18081,17'd17843,17'd12421,17'd18197,17'd18198,17'd15053,17'd16204,17'd13362,17'd12262,17'd12115,17'd17604,17'd17843,17'd16321,17'd12415,17'd17235,17'd18199,17'd18199,17'd17475,17'd17727,17'd18084,17'd18200,17'd12860,17'd13884,17'd12111,17'd10853,17'd10856,17'd9044,17'd18201,17'd18202,17'd16691,17'd18203,17'd11968,17'd18204,17'd13141,17'd18205,17'd15307,17'd15576,17'd17243,17'd18206,17'd18207,17'd18088,17'd18208,17'd11538,17'd18209,17'd18210,17'd18211,17'd1045,17'd132,17'd134,17'd1197,17'd133,17'd1481,17'd1481,17'd1481,17'd1481,17'd130,17'd130,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd135,17'd132,17'd133,17'd135,17'd3811,17'd18212,17'd18213,17'd18214,17'd16222,17'd18215,17'd18216,17'd18217,17'd18218,17'd18219,17'd18220,17'd18221,17'd17992,17'd18222,17'd18223,17'd18224,17'd18225,17'd18226,17'd18227,17'd18228,17'd17503,17'd18229,17'd9918,17'd10634,17'd18230,17'd12892,17'd8767,17'd8616,17'd16354,17'd16472,17'd16473,17'd15840,17'd17387,17'd18231,17'd18232,17'd17266,17'd18233,17'd18234,17'd18235,17'd18236,17'd18237,17'd15213,17'd15212,17'd15211,17'd16478,17'd16359,17'd15717,17'd18238,17'd18239,17'd18008,17'd18120,17'd18240,17'd18241,17'd18121,17'd18242,17'd18243,17'd18244,17'd18245,17'd18246,17'd18246,17'd16941,17'd18006,17'd18010,17'd17768,17'd16829,17'd18247,17'd16829,17'd17771,17'd17890,17'd18012,17'd17891,17'd18248,17'd16110,17'd17274,17'd15843,17'd18249,17'd18249,17'd18250,17'd18128,17'd15844,17'd16359,17'd16836,17'd16114,17'd18251,17'd18252,17'd16364,17'd18253,17'd18254,17'd17170,17'd18255,17'd17281,17'd17062,17'd17901,17'd18256,17'd17063,17'd16845,17'd17064,17'd17171,17'd17531,17'd17778,17'd18020,17'd18257,17'd18258,17'd18021,17'd15603,17'd15475,17'd16119,17'd15337,17'd15337,17'd17065,17'd18259,17'd18260,17'd18261,17'd18023,17'd14050,17'd18262,17'd18263,17'd18264,17'd16620,17'd16621,17'd13415,17'd17412,17'd16958,17'd18265,17'd18266,17'd14308,17'd14058,17'd18267,17'd18268,17'd18269,17'd18270,17'd5495,17'd18143,17'd3071,17'd634,17'd1683,17'd18271,17'd1684,17'd1268,17'd973,17'd9671,17'd18272,17'd1817,17'd4232,17'd5501,17'd5501,17'd5635,17'd17073,17'd11444,17'd11191,17'd8795,17'd8795,17'd12018,17'd12018,17'd12019,17'd12487,17'd11723,17'd12178,17'd12021,17'd12021,17'd16135,17'd15866,17'd16961,17'd16741,17'd18147,17'd16742,17'd17182,17'd16962,17'd18148,17'd17549,17'd16743,17'd16629,17'd16630,17'd16743,17'd16629,17'd16857,17'd14596,17'd8324,17'd18273,17'd13294,17'd8503,17'd7034,17'd12182,17'd12492,17'd14866,17'd7875,17'd5950,17'd6089,17'd9122,17'd4084,17'd189,17'd267,17'd2255,17'd2115
},
'{
17'd2423,17'd16636,17'd3430,17'd1127,17'd1689,17'd1688,17'd2422,17'd1831,17'd4247,17'd466,17'd3,17'd1275,17'd1275,17'd2933,17'd8814,17'd2423,17'd16636,17'd806,17'd977,17'd978,17'd3753,17'd3753,17'd8040,17'd8340,17'd10913,17'd18274,17'd10912,17'd17664,17'd10912,17'd10913,17'd17664,17'd7712,17'd5205,17'd6,17'd5,17'd23,17'd21,17'd21,17'd21,17'd21,17'd22,17'd22,17'd1832,17'd1832,17'd285,17'd286,17'd27,17'd28,17'd18037,17'd3910,17'd4579,17'd2947,17'd1704,17'd18275,17'd309,17'd18276,17'd18277,17'd18278,17'd18279,17'd18280,17'd18281,17'd18282,17'd18283,17'd18284,17'd18285,17'd18286,17'd18287,17'd18288,17'd14331,17'd18289,17'd17310,17'd15507,17'd15507,17'd18290,17'd18291,17'd18292,17'd10422,17'd18293,17'd15638,17'd18294,17'd16981,17'd18169,17'd18295,17'd18296,17'd18172,17'd18173,17'd14470,17'd14470,17'd13969,17'd13969,17'd13840,17'd13840,17'd14891,17'd14621,17'd12955,17'd13093,17'd13094,17'd12218,17'd11913,17'd11362,17'd17205,17'd17572,17'd17445,17'd17810,17'd15769,17'd16165,17'd16290,17'd16165,17'd15769,17'd16411,17'd17810,17'd18297,17'd18298,17'd18299,17'd18300,17'd18301,17'd18302,17'd18063,17'd18303,17'd15145,17'd17326,17'd17326,17'd16416,17'd18304,17'd18305,17'd18306,17'd9848,17'd9310,17'd16666,17'd8703,17'd9446,17'd18307,17'd18307,17'd9586,17'd17947,17'd18180,17'd17946,17'd17948,17'd18308,17'd18309,17'd18310,17'd18311,17'd18069,17'd17824,17'd17952,17'd15409,17'd15543,17'd13860,17'd18312,17'd18313,17'd18314,17'd10444,17'd18315,17'd18316,17'd10582,17'd18317,17'd18318,17'd12400,17'd18319,17'd15671,17'd12986,17'd12705,17'd18320,17'd17832,17'd12088,17'd17834,17'd12570,17'd13249,17'd18321,17'd18322,17'd12856,17'd13135,17'd16320,17'd18323,17'd18324,17'd16065,17'd10992,17'd10169,17'd9619,17'd18325,17'd15688,17'd11132,17'd18326,17'd18327,17'd12422,17'd18328,17'd12858,17'd12111,17'd12110,17'd16321,17'd17603,17'd12719,17'd12260,17'd18081,17'd17843,17'd18329,17'd18197,17'd18198,17'd15053,17'd12422,17'd13362,17'd12262,17'd12115,17'd18330,17'd12581,17'd13517,17'd16913,17'd17475,17'd17969,17'd18331,17'd17235,17'd17727,17'd16558,17'd16913,17'd12860,17'd13644,17'd11962,17'd10472,17'd18332,17'd12118,17'd13139,17'd8581,17'd17128,17'd11968,17'd17238,17'd8107,17'd15442,17'd8586,17'd18333,17'd18334,17'd18335,17'd18336,17'd16807,17'd18336,17'd18337,17'd18338,17'd17024,17'd15958,17'd11152,17'd133,17'd132,17'd132,17'd133,17'd133,17'd1481,17'd1481,17'd1481,17'd1481,17'd130,17'd130,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd2698,17'd132,17'd132,17'd135,17'd3168,17'd2863,17'd4817,17'd18339,17'd18340,17'd18341,17'd18342,17'd18343,17'd18344,17'd18345,17'd18346,17'd18347,17'd18348,17'd18349,17'd18350,17'd18351,17'd18352,17'd18226,17'd18353,17'd18354,17'd18355,17'd18356,17'd9510,17'd11425,17'd9512,17'd13027,17'd11992,17'd8616,17'd11832,17'd11988,17'd18357,17'd15840,17'd17387,17'd18358,17'd18232,17'd18359,17'd17265,17'd18234,17'd17160,17'd18360,17'd17044,17'd15213,17'd15212,17'd15211,17'd15593,17'd15593,17'd18015,17'd18361,17'd18126,17'd18124,17'd18362,17'd18240,17'd18121,17'd18121,17'd18363,17'd18010,17'd18125,17'd18364,17'd18365,17'd18246,17'd16941,17'd18122,17'd18010,17'd17769,17'd17768,17'd16829,17'd17768,17'd16829,17'd18011,17'd18126,17'd18366,17'd18367,17'd17891,17'd17773,17'd16945,17'd15466,17'd15466,17'd17526,17'd16355,17'd18368,17'd16363,17'd16360,17'd16113,17'd16239,17'd12604,17'd18252,17'd18369,17'd17897,17'd18370,17'd17899,17'd16952,17'd17062,17'd17901,17'd17283,17'd17063,17'd17064,17'd17064,17'd16246,17'd17531,17'd17653,17'd18371,17'd18020,17'd18372,17'd18131,17'd15723,17'd15475,17'd15475,17'd15336,17'd16120,17'd16371,17'd18373,17'd18374,17'd18375,17'd18261,17'd12622,17'd18262,17'd15992,17'd18376,17'd13682,17'd18377,17'd17071,17'd18378,17'd17072,17'd18265,17'd18379,17'd18380,17'd18381,17'd14058,17'd18268,17'd18382,17'd12317,17'd18383,17'd18384,17'd18385,17'd18386,17'd251,17'd17185,17'd18387,17'd263,17'd803,17'd1821,17'd13290,17'd1816,17'd4404,17'd5501,17'd5501,17'd4065,17'd17073,17'd9945,17'd11191,17'd8795,17'd8795,17'd12018,17'd12018,17'd10077,17'd12487,17'd11723,17'd12178,17'd12021,17'd12021,17'd16135,17'd15866,17'd16384,17'd16741,17'd18147,17'd16742,17'd18388,17'd17182,17'd18148,17'd17549,17'd15624,17'd16137,17'd15624,17'd16743,17'd16629,17'd16857,17'd14596,17'd15870,17'd18389,17'd16261,17'd9801,17'd8330,17'd12492,17'd12492,17'd8503,17'd9801,17'd18149,17'd13294,17'd8505,17'd4084,17'd641,17'd18390,17'd255,17'd2255
},
'{
17'd12647,17'd6419,17'd5196,17'd5196,17'd3250,17'd2422,17'd1831,17'd1831,17'd2595,17'd12,17'd1275,17'd806,17'd806,17'd806,17'd806,17'd16636,17'd21,17'd23,17'd4,17'd7,17'd5205,17'd8040,17'd8338,17'd8338,17'd13429,17'd8338,17'd8338,17'd8339,17'd8340,17'd8040,17'd5205,17'd5205,17'd3753,17'd5,17'd24,17'd24,17'd22,17'd22,17'd22,17'd23,17'd23,17'd22,17'd1832,17'd1832,17'd285,17'd286,17'd27,17'd6744,17'd3910,17'd3756,17'd2604,17'd1976,17'd18150,17'd18391,17'd18392,17'd18153,17'd18393,17'd18394,17'd18395,17'd16641,17'd18396,17'd18397,17'd18398,17'd18399,17'd18400,17'd18401,17'd18402,17'd18050,17'd14202,17'd17310,17'd18403,17'd18404,17'd15507,17'd18290,17'd18166,17'd18405,17'd10422,17'd18406,17'd17200,17'd18407,17'd18408,17'd18169,17'd18170,17'd18409,17'd18410,17'd18411,17'd14764,17'd12530,17'd13969,17'd13969,17'd15764,17'd14764,17'd14621,17'd12955,17'd12528,17'd12528,17'd12814,17'd12530,17'd11628,17'd18412,17'd18174,17'd17572,17'd17320,17'd15902,17'd16165,17'd16290,17'd17575,17'd18413,17'd17448,17'd18414,17'd15899,17'd18061,17'd18415,17'd18416,17'd18417,17'd18418,17'd18418,17'd14351,17'd14481,17'd15649,17'd17326,17'd16416,17'd15778,17'd15271,17'd14638,17'd13104,17'd9310,17'd18419,17'd15537,17'd18420,17'd18421,17'd18422,17'd18423,17'd10126,17'd18424,17'd18425,17'd17822,17'd18426,17'd18427,17'd18310,17'd18310,17'd18068,17'd17824,17'd17952,17'd18428,17'd16670,17'd15277,17'd13487,17'd18429,17'd18430,17'd18431,17'd18432,17'd18433,17'd18434,17'd18188,17'd14919,17'd11935,17'd12709,17'd18435,17'd18436,17'd13127,17'd17225,17'd18437,17'd13505,17'd13638,17'd11790,17'd18438,17'd15677,17'd18439,17'd12995,17'd18440,17'd16069,17'd18441,17'd18442,17'd16549,17'd16549,17'd9885,17'd12116,17'd17839,17'd10479,17'd10476,17'd14673,17'd13762,17'd12422,17'd18328,17'd12259,17'd15809,17'd13763,17'd16321,17'd17603,17'd18197,17'd17843,17'd18328,17'd18328,17'd17843,17'd17967,17'd17722,17'd17722,17'd18443,17'd18444,17'd15810,17'd18445,17'd18446,17'd18447,17'd13136,17'd14930,17'd17726,17'd18448,17'd17013,17'd16560,17'd17013,17'd17235,17'd18449,17'd15687,17'd12860,17'd18450,17'd14673,17'd11671,17'd9040,17'd17126,17'd15812,17'd17482,17'd17241,17'd7786,17'd18451,17'd18086,17'd15574,17'd18452,17'd18453,17'd18454,17'd10345,17'd18455,17'd16080,17'd18456,17'd11146,17'd17736,17'd18457,17'd18458,17'd542,17'd356,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd132,17'd134,17'd132,17'd2698,17'd5466,17'd18459,17'd18460,17'd18461,17'd18462,17'd18463,17'd18464,17'd18465,17'd18466,17'd18467,17'd18468,17'd18469,17'd18470,17'd18471,17'd18472,17'd18473,17'd18474,17'd18475,17'd18476,17'd18477,17'd18478,17'd18479,17'd9378,17'd11833,17'd11695,17'd9075,17'd11992,17'd18480,17'd11988,17'd10768,17'd15713,17'd18481,17'd18482,17'd18483,17'd18484,17'd18233,17'd17265,17'd18485,17'd18486,17'd17274,17'd15977,17'd16729,17'd15844,17'd16360,17'd17054,17'd18361,17'd18127,17'd18487,17'd18123,17'd18488,17'd18488,17'd18488,17'd18488,17'd18488,17'd16941,17'd18125,17'd18125,17'd18365,17'd18365,17'd18489,17'd18489,17'd18490,17'd18491,17'd18010,17'd18010,17'd18125,17'd16829,17'd16829,17'd18364,17'd18492,17'd18126,17'd17890,17'd18013,17'd17394,17'd15975,17'd15466,17'd18493,17'd18494,17'd16355,17'd16359,17'd16362,17'd16480,17'd18495,17'd18496,17'd16114,17'd13153,17'd15089,17'd18497,17'd17170,17'd16952,17'd16841,17'd15724,17'd15723,17'd16118,17'd16246,17'd16845,17'd17172,17'd16370,17'd17531,17'd17902,17'd17902,17'd17531,17'd16953,17'd15852,17'd15604,17'd15603,17'd15475,17'd16247,17'd16121,17'd18498,17'd18499,17'd18260,17'd18500,17'd18023,17'd15611,17'd18501,17'd18502,17'd18503,17'd18504,17'd17289,17'd17908,17'd15100,17'd18029,17'd18505,17'd18506,17'd18507,17'd18508,17'd18509,17'd18510,17'd18511,17'd18512,17'd8482,17'd18513,17'd18514,17'd18515,17'd18516,17'd17422,17'd456,17'd273,17'd603,17'd950,17'd1251,17'd5367,17'd18517,17'd14864,17'd4062,17'd4872,17'd8018,17'd8491,17'd9405,17'd9405,17'd11592,17'd11722,17'd11593,17'd12487,17'd11723,17'd12178,17'd12021,17'd12021,17'd15238,17'd15866,17'd16383,17'd16493,17'd16742,17'd16742,17'd18147,17'd16742,17'd16627,17'd15489,17'd15624,17'd15868,17'd15624,17'd15624,17'd15868,17'd15624,17'd8179,17'd8325,17'd10654,17'd10654,17'd9801,17'd8503,17'd8810,17'd7876,17'd9801,17'd11333,17'd8811,17'd12779,17'd8332,17'd5192,17'd271,17'd268,17'd266,17'd459
},
'{
17'd4886,17'd5196,17'd7711,17'd7711,17'd2422,17'd2422,17'd1831,17'd2594,17'd466,17'd3,17'd1275,17'd2933,17'd806,17'd806,17'd12,17'd2423,17'd21,17'd23,17'd6,17'd7,17'd5205,17'd8040,17'd8338,17'd8338,17'd13429,17'd13429,17'd8338,17'd8338,17'd8040,17'd8040,17'd5205,17'd3753,17'd5,17'd5,17'd24,17'd24,17'd22,17'd22,17'd23,17'd23,17'd23,17'd22,17'd1832,17'd285,17'd286,17'd286,17'd28,17'd288,17'd3754,17'd3435,17'd2946,17'd1704,17'd2788,17'd488,17'd18518,17'd1440,17'd18519,17'd18520,17'd18521,17'd18522,17'd18523,17'd18524,17'd18525,17'd14996,17'd16756,17'd18526,17'd18163,17'd14758,17'd18527,17'd17310,17'd18403,17'd13589,17'd15507,17'd13963,17'd16650,17'd18528,17'd18406,17'd18529,17'd18530,17'd17094,17'd18408,17'd18295,17'd18531,17'd18532,17'd15383,17'd14764,17'd12530,17'd12530,17'd13969,17'd13969,17'd15764,17'd14764,17'd14890,17'd12955,17'd12528,17'd12528,17'd12218,17'd11913,17'd11362,17'd18533,17'd17572,17'd17207,17'd16034,17'd15902,17'd16165,17'd16768,17'd18413,17'd18534,17'd18414,17'd17690,17'd6462,17'd18535,17'd18536,17'd18537,17'd18538,17'd18539,17'd18540,17'd14351,17'd17698,17'd15776,17'd17326,17'd15650,17'd15533,17'd18541,17'd18306,17'd14109,17'd18542,17'd18543,17'd15537,17'd18420,17'd18421,17'd18422,17'd13483,17'd10126,17'd18544,17'd18545,17'd17586,17'd18546,17'd18311,17'd18311,17'd18310,17'd18068,17'd17824,17'd17952,17'd17587,17'd17218,17'd18547,17'd18548,17'd18549,17'd18550,17'd18551,17'd18552,17'd17114,17'd18553,17'd17118,17'd12562,17'd13996,17'd12988,17'd18554,17'd13244,17'd12393,17'd12235,17'd17832,17'd12094,17'd12403,17'd18438,17'd18555,17'd13250,17'd15686,17'd13882,17'd13000,17'd11526,17'd13255,17'd10743,17'd15566,17'd18556,17'd12116,17'd11276,17'd12863,17'd11132,17'd11808,17'd11964,17'd16204,17'd18328,17'd12581,17'd13136,17'd13763,17'd13763,17'd16321,17'd17603,17'd18557,17'd12582,17'd17843,17'd17843,17'd18558,17'd17967,17'd18559,17'd18197,17'd18443,17'd13516,17'd18560,17'd18445,17'd18561,17'd12114,17'd12995,17'd14672,17'd18562,17'd18448,17'd17726,17'd17235,17'd17013,17'd16560,17'd18563,17'd15687,17'd18564,17'd18565,17'd12584,17'd17232,17'd8725,17'd18566,17'd12120,17'd10179,17'd12265,17'd15440,17'd18567,17'd18568,17'd18569,17'd18570,17'd17973,17'd18571,17'd10032,17'd18572,17'd18573,17'd18574,17'd18575,17'd18576,17'd18577,17'd7980,17'd8132,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd132,17'd134,17'd132,17'd1759,17'd18578,17'd4338,17'd18579,17'd18580,17'd18581,17'd18582,17'd18583,17'd18584,17'd18585,17'd18586,17'd18587,17'd18588,17'd18589,17'd18590,17'd18591,17'd18352,17'd18592,17'd18593,17'd18594,17'd18595,17'd18596,17'd18479,17'd9917,17'd10888,17'd11425,17'd11425,17'd11425,17'd9071,17'd11988,17'd18597,17'd15713,17'd18598,17'd18599,17'd18600,17'd18601,17'd18602,17'd17265,17'd18603,17'd18604,17'd16236,17'd17053,17'd16729,17'd15844,17'd15717,17'd18249,17'd18605,17'd18606,17'd18244,17'd18607,17'd18488,17'd18488,17'd18488,17'd18122,17'd16941,17'd16941,17'd18244,17'd18244,17'd18125,17'd18246,17'd18489,17'd18608,17'd18609,17'd18610,17'd18611,17'd18612,17'd18244,17'd18364,17'd18364,17'd18364,17'd18364,17'd18364,17'd18126,17'd17890,17'd18013,17'd17401,17'd18613,17'd15843,17'd15716,17'd15717,17'd15593,17'd16359,17'd18614,17'd18615,17'd18616,17'd18617,17'd15980,17'd14565,17'd15332,17'd18618,17'd17170,17'd16841,17'd15605,17'd17282,17'd15852,17'd16118,17'd17063,17'd17171,17'd17529,17'd17530,17'd17653,17'd17778,17'd17778,17'd17530,17'd16118,17'd15604,17'd15723,17'd15603,17'd16247,17'd16121,17'd18498,17'd18619,17'd18620,17'd17904,17'd18621,17'd17408,17'd17174,17'd18622,17'd18623,17'd18624,17'd17071,17'd17908,17'd15100,17'd18266,17'd18505,17'd18506,17'd18625,17'd18626,17'd18627,17'd18628,17'd12174,17'd18629,17'd6404,17'd18630,17'd18631,17'd18632,17'd18633,17'd1543,17'd965,17'd646,17'd1098,17'd601,17'd1390,17'd4066,17'd7521,17'd6575,17'd4232,17'd4872,17'd14983,17'd8491,17'd9405,17'd9405,17'd11592,17'd11722,17'd11593,17'd12487,17'd11723,17'd12178,17'd11873,17'd11873,17'd15238,17'd15623,17'd16383,17'd16493,17'd18147,17'd16742,17'd18147,17'd16742,17'd16962,17'd15489,17'd18634,17'd18635,17'd18634,17'd18634,17'd15868,17'd15624,17'd8325,17'd8325,17'd9668,17'd10654,17'd8503,17'd8503,17'd8810,17'd11333,17'd8656,17'd11333,17'd16002,17'd12779,17'd8035,17'd5192,17'd260,17'd271,17'd257,17'd266
},
'{
17'd7214,17'd7214,17'd7711,17'd7545,17'd2422,17'd3252,17'd1831,17'd2594,17'd0,17'd806,17'd2933,17'd2933,17'd806,17'd2423,17'd12,17'd2423,17'd25,17'd4,17'd6,17'd5205,17'd8040,17'd8040,17'd8338,17'd8338,17'd13429,17'd13429,17'd8338,17'd8338,17'd8040,17'd5793,17'd3753,17'd3753,17'd5,17'd5,17'd24,17'd24,17'd23,17'd23,17'd23,17'd23,17'd23,17'd22,17'd1832,17'd1832,17'd285,17'd286,17'd28,17'd4431,17'd3434,17'd4739,17'd2431,17'd1138,17'd995,17'd18636,17'd18637,17'd18638,17'd18639,17'd17427,17'd18640,17'd18641,17'd18642,17'd18643,17'd18644,17'd18645,17'd18646,17'd18647,17'd18648,17'd18649,17'd18650,17'd17435,17'd13448,17'd16509,17'd18651,17'd18652,17'd18653,17'd18406,17'd18529,17'd15895,17'd18530,17'd17094,17'd18654,17'd18170,17'd18531,17'd18532,17'd18173,17'd14622,17'd13969,17'd13969,17'd14891,17'd14764,17'd14764,17'd14621,17'd12955,17'd12955,17'd12955,17'd14890,17'd12361,17'd12532,17'd17941,17'd18655,17'd18656,17'd18657,17'd16034,17'd15902,17'd18413,17'd17692,17'd18534,17'd17448,17'd18414,17'd18658,17'd18061,17'd18659,17'd18660,17'd18661,17'd18540,17'd18662,17'd18662,17'd14900,17'd16176,17'd16886,17'd18663,17'd18664,17'd18541,17'd18665,17'd18666,17'd9164,17'd18542,17'd10127,17'd9313,17'd9166,17'd9850,17'd18667,17'd10126,17'd10292,17'd18425,17'd18545,17'd18426,17'd18427,17'd18668,17'd18668,17'd18311,17'd18068,17'd17952,17'd18428,17'd17587,17'd15277,17'd13739,17'd18669,17'd18430,17'd18670,17'd18671,17'd18672,17'd18673,17'd18674,17'd18675,17'd16309,17'd12848,17'd12709,17'd13501,17'd13127,17'd17225,17'd12235,17'd12236,17'd18676,17'd11945,17'd18677,17'd18678,17'd12854,17'd15808,17'd18679,17'd10475,17'd18680,17'd16683,17'd11277,17'd11277,17'd12116,17'd10479,17'd11528,17'd10991,17'd13886,17'd14673,17'd13762,17'd12996,17'd12719,17'd12420,17'd12419,17'd12110,17'd12419,17'd11958,17'd12581,17'd12582,17'd12582,17'd17843,17'd17843,17'd18197,17'd17722,17'd18197,17'd18557,17'd18681,17'd13516,17'd18682,17'd18560,17'd18683,17'd12259,17'd18684,17'd14524,17'd18685,17'd18448,17'd17726,17'd17235,17'd17013,17'd16914,17'd15811,17'd14672,17'd15434,17'd13646,17'd10330,17'd9743,17'd14675,17'd18686,17'd9622,17'd10179,17'd7786,17'd10180,17'd18086,17'd18687,17'd18688,17'd18689,17'd18690,17'd18691,17'd18692,17'd18693,17'd18694,17'd18695,17'd18696,17'd18697,17'd16578,17'd16090,17'd18698,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd132,17'd134,17'd132,17'd134,17'd6055,17'd18699,17'd18700,17'd18701,17'd18702,17'd18703,17'd18704,17'd18705,17'd18706,17'd18707,17'd18708,17'd18709,17'd18710,17'd18711,17'd18712,17'd18713,17'd18714,17'd18715,17'd18716,17'd18717,17'd18718,17'd18719,17'd9376,17'd9508,17'd9375,17'd9375,17'd9224,17'd18720,17'd11552,17'd18357,17'd15713,17'd18598,17'd18721,17'd17643,17'd18722,17'd18723,17'd18724,17'd18725,17'd18726,17'd17402,17'd17053,17'd17055,17'd17055,17'd18015,17'd18727,17'd18728,17'd18729,17'd18607,17'd18730,17'd18730,17'd18121,17'd18488,17'd18122,17'd18243,17'd18243,17'd18243,17'd18612,17'd18243,17'd18612,17'd18608,17'd18731,17'd18732,17'd18732,17'd18733,17'd18608,17'd18246,17'd18246,17'd18244,17'd18244,17'd18125,17'd18125,17'd18487,17'd18126,17'd18734,17'd18735,17'd18361,17'd18736,17'd15843,17'd15716,17'd18128,17'd18128,17'd18737,17'd18368,17'd18738,17'd18739,17'd15330,17'd8760,17'd18740,17'd16365,17'd17898,17'd17170,17'd17406,17'd17528,17'd17282,17'd16843,17'd16118,17'd16246,17'd17529,17'd17529,17'd17530,17'd17653,17'd17902,17'd17778,17'd16370,17'd15852,17'd15604,17'd15723,17'd16371,17'd16247,17'd18741,17'd18619,17'd18741,17'd18742,17'd18500,17'd18743,17'd15856,17'd18744,17'd18745,17'd18746,17'd18747,17'd17908,17'd18748,17'd18379,17'd18749,17'd18750,17'd18751,17'd18752,17'd18753,17'd18754,17'd11865,17'd18755,17'd18756,17'd18757,17'd18758,17'd18759,17'd435,17'd281,17'd402,17'd256,17'd645,17'd1821,17'd18272,17'd1817,17'd4404,17'd4062,17'd4232,17'd4717,17'd7684,17'd8170,17'd9405,17'd9405,17'd11592,17'd11592,17'd11593,17'd12487,17'd11723,17'd12178,17'd11873,17'd11873,17'd15238,17'd15623,17'd16384,17'd16384,17'd16493,17'd16742,17'd16742,17'd18147,17'd17548,17'd15489,17'd18634,17'd18635,17'd18634,17'd18634,17'd18635,17'd15624,17'd8325,17'd8325,17'd7199,17'd17074,17'd8810,17'd8810,17'd11196,17'd11333,17'd11333,17'd10793,17'd12779,17'd12779,17'd8035,17'd2774,17'd271,17'd646,17'd263,17'd266
},
'{
17'd7372,17'd7214,17'd7545,17'd7545,17'd3252,17'd2422,17'd1831,17'd4247,17'd1,17'd283,17'd1275,17'd2933,17'd806,17'd2423,17'd12,17'd806,17'd25,17'd4,17'd7,17'd5205,17'd8040,17'd8040,17'd8338,17'd8338,17'd13429,17'd8338,17'd8338,17'd8040,17'd8040,17'd5793,17'd3753,17'd3753,17'd5,17'd24,17'd24,17'd24,17'd23,17'd23,17'd23,17'd4,17'd23,17'd22,17'd1832,17'd285,17'd286,17'd286,17'd28,17'd3907,17'd3104,17'd1975,17'd2433,17'd827,17'd485,17'd1845,17'd18760,17'd18761,17'd18762,17'd18763,17'd18764,17'd18765,17'd18159,17'd18766,17'd18644,17'd18767,17'd18768,17'd18769,17'd16273,17'd17676,17'd18770,17'd16977,17'd13589,17'd16401,17'd17566,17'd18771,17'd18772,17'd18406,17'd15895,17'd17094,17'd16404,17'd18773,17'd18169,17'd17937,17'd18058,17'd18173,17'd14622,17'd15764,17'd13969,17'd13969,17'd14891,17'd14764,17'd14621,17'd12955,17'd13093,17'd13093,17'd12955,17'd12218,17'd12532,17'd17204,17'd18774,17'd18656,17'd17207,17'd17445,17'd15902,17'd15902,17'd17692,17'd18775,17'd18776,17'd18777,17'd16519,17'd18778,17'd18779,17'd18299,17'd18780,17'd18781,17'd18540,17'd18782,17'd18782,17'd17698,17'd16176,17'd16886,17'd16416,17'd18783,17'd18784,17'd18785,17'd9707,17'd9164,17'd18542,17'd10818,17'd9166,17'd9312,17'd9445,17'd9444,17'd18786,17'd18787,17'd18545,17'd17333,17'd18426,17'd18788,17'd18668,17'd18668,17'd18311,17'd18789,17'd18428,17'd18790,17'd16536,17'd14111,17'd18791,17'd11772,17'd18792,17'd18793,17'd18794,17'd18795,17'd18796,17'd18797,17'd13748,17'd18798,17'd12848,17'd12567,17'd12558,17'd11934,17'd12235,17'd12087,17'd18799,17'd18800,17'd18801,17'd18802,17'd18803,17'd18804,17'd18805,17'd11519,17'd10328,17'd18441,17'd10856,17'd16070,17'd14928,17'd11134,17'd15943,17'd10991,17'd13886,17'd14810,17'd11807,17'd12996,17'd12719,17'd16321,17'd12109,17'd12110,17'd12419,17'd12420,17'd12719,17'd17843,17'd12582,17'd12582,17'd17843,17'd12581,17'd17722,17'd17722,17'd18557,17'd18806,17'd18444,17'd13516,17'd17968,17'd12115,17'd11957,17'd13763,17'd18807,17'd16915,17'd18685,17'd18685,17'd17235,17'd17475,17'd17013,17'd15687,17'd15811,17'd13884,17'd14131,17'd16068,17'd9885,17'd9621,17'd18808,17'd8252,17'd11968,17'd15693,17'd15440,17'd10861,17'd18809,17'd15306,17'd14393,17'd18810,17'd18811,17'd12730,17'd18812,17'd18813,17'd18814,17'd18815,17'd18696,17'd16087,17'd7980,17'd1045,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd132,17'd134,17'd132,17'd132,17'd10492,17'd18816,17'd18817,17'd18818,17'd18819,17'd18703,17'd18820,17'd18821,17'd18822,17'd18823,17'd18824,17'd18825,17'd18826,17'd18827,17'd18828,17'd18829,17'd18830,17'd18831,17'd18832,17'd18833,17'd18718,17'd18719,17'd9376,17'd18834,17'd18834,17'd18835,17'd9914,17'd18836,17'd17641,17'd18357,17'd15840,17'd18598,17'd18837,17'd17643,17'd18003,17'd18838,17'd18839,17'd18840,17'd18486,17'd17773,17'd15976,17'd16728,17'd16728,17'd16832,17'd18841,17'd18842,17'd18611,17'd18843,17'd18844,17'd18241,17'd18241,17'd18730,17'd18730,17'd18611,17'd18612,17'd18612,17'd18612,17'd18608,17'd18608,17'd18608,17'd18608,17'd18733,17'd18733,17'd18732,17'd18732,17'd18731,17'd18845,17'd18365,17'd18246,17'd18244,17'd18244,17'd18846,17'd18487,17'd18487,17'd18734,17'd18735,17'd18361,17'd16945,17'd15843,17'd15592,17'd18128,17'd18128,17'd18368,17'd18738,17'd18847,17'd18848,17'd15330,17'd18016,17'd18740,17'd18849,17'd17898,17'd18850,17'd18851,17'd17528,17'd16843,17'd16118,17'd15604,17'd17532,17'd17532,17'd17529,17'd17653,17'd17902,17'd17778,17'd18019,17'd16118,17'd15604,17'd15723,17'd17065,17'd16247,17'd18741,17'd18498,17'd18741,17'd18134,17'd18852,17'd18853,17'd18854,17'd18855,17'd18856,17'd18857,17'd18858,17'd16958,17'd18748,17'd18379,17'd18859,17'd17909,17'd18860,17'd18861,17'd12769,17'd18862,17'd18863,17'd18864,17'd4054,17'd18865,17'd18866,17'd763,17'd18867,17'd18868,17'd401,17'd2255,17'd409,17'd2577,17'd1392,17'd1816,17'd4404,17'd4062,17'd4404,17'd4407,17'd7684,17'd8170,17'd9405,17'd10076,17'd10076,17'd11722,17'd11593,17'd12487,17'd11723,17'd11723,17'd11329,17'd11873,17'd15238,17'd15238,17'd16384,17'd16383,17'd16384,17'd16742,17'd16742,17'd18147,17'd16626,17'd16136,17'd18635,17'd18635,17'd18634,17'd18634,17'd18635,17'd18634,17'd8325,17'd16260,17'd18869,17'd17074,17'd8655,17'd8810,17'd11196,17'd11333,17'd11880,17'd11880,17'd12779,17'd12779,17'd8035,17'd5192,17'd260,17'd271,17'd256,17'd459
},
'{
17'd7372,17'd7214,17'd7711,17'd7545,17'd2422,17'd1831,17'd4247,17'd2,17'd283,17'd283,17'd1275,17'd1275,17'd806,17'd2423,17'd806,17'd2933,17'd4,17'd6,17'd5205,17'd5205,17'd8040,17'd8040,17'd8338,17'd8338,17'd8338,17'd8338,17'd8040,17'd8040,17'd8040,17'd3753,17'd3753,17'd3753,17'd24,17'd24,17'd24,17'd24,17'd23,17'd23,17'd4,17'd4,17'd23,17'd23,17'd1832,17'd1832,17'd285,17'd27,17'd4430,17'd3755,17'd3105,17'd14447,17'd14449,17'd2789,17'd308,17'd18870,17'd18871,17'd18872,17'd18873,17'd18874,17'd18875,17'd18876,17'd18159,17'd18877,17'd18161,17'd18878,17'd18769,17'd18879,17'd18880,17'd18881,17'd16647,17'd18882,17'd18883,17'd16875,17'd17440,17'd17933,17'd18293,17'd18406,17'd17094,17'd16878,17'd16404,17'd18773,17'd18170,17'd18058,17'd18532,17'd18173,17'd16027,17'd16163,17'd13969,17'd13969,17'd14764,17'd14890,17'd12955,17'd13093,17'd13093,17'd12955,17'd14621,17'd12361,17'd18884,17'd17689,17'd18655,17'd18656,17'd18657,17'd17445,17'd15902,17'd16290,17'd18413,17'd18775,17'd18885,17'd18886,17'd18887,17'd18888,17'd18889,17'd18890,17'd18891,17'd18892,17'd18782,17'd14481,17'd16885,17'd18893,17'd15269,17'd18894,17'd15654,17'd18895,17'd18666,17'd9707,17'd9583,17'd11631,17'd11095,17'd9311,17'd18896,17'd18896,17'd9445,17'd9445,17'd18897,17'd17947,17'd17333,17'd17822,17'd18427,17'd18668,17'd18898,17'd18898,17'd18899,17'd18900,17'd18790,17'd18901,17'd18902,17'd13859,17'd18903,17'd18904,17'd18905,17'd18906,17'd18907,17'd18908,17'd18909,17'd18910,17'd18911,17'd13355,17'd13355,17'd14372,17'd14661,17'd11934,17'd15674,17'd15423,17'd12243,17'd18912,17'd18913,17'd18914,17'd12258,17'd13364,17'd18915,17'd10741,17'd18916,17'd9740,17'd10479,17'd11134,17'd11134,17'd11528,17'd14518,17'd10739,17'd14931,17'd11520,17'd13520,17'd15053,17'd16321,17'd12109,17'd12414,17'd12109,17'd16321,17'd17603,17'd18917,17'd12582,17'd16204,17'd16204,17'd12582,17'd18917,17'd15053,17'd15053,17'd18806,17'd17604,17'd18082,17'd12115,17'd17968,17'd16204,17'd12420,17'd12256,17'd16798,17'd18918,17'd18685,17'd18685,17'd17235,17'd17235,17'd17726,17'd15687,17'd12860,17'd13644,17'd15175,17'd14518,17'd9339,17'd8410,17'd18919,17'd18203,17'd15693,17'd18920,17'd14681,17'd18921,17'd15305,17'd18922,17'd8429,17'd18923,17'd18924,17'd15196,17'd18925,17'd18926,17'd18927,17'd11540,17'd10756,17'd18928,17'd133,17'd134,17'd132,17'd11541,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd3168,17'd18929,17'd18930,17'd18931,17'd18932,17'd18933,17'd18934,17'd18935,17'd18936,17'd18937,17'd18938,17'd18939,17'd18940,17'd18941,17'd18942,17'd18943,17'd18944,17'd18945,17'd18946,17'd18947,17'd18948,17'd18949,17'd9376,17'd18950,17'd18950,17'd18951,17'd18835,17'd9507,17'd18597,17'd10768,17'd15840,17'd17387,17'd16831,17'd18002,17'd18952,17'd18005,17'd18953,17'd18840,17'd18486,17'd17401,17'd15715,17'd17525,17'd17167,17'd18954,17'd18735,17'd18729,17'd18955,17'd18956,17'd18956,17'd18955,17'd18957,17'd18957,17'd18957,17'd18957,17'd18733,17'd18958,17'd18958,17'd18732,17'd18733,17'd18733,17'd18958,17'd18733,17'd18733,17'd18732,17'd18732,17'd18959,17'd18960,17'd18732,17'd18733,17'd18958,17'd18612,17'd18243,17'd18961,17'd18846,17'd18962,17'd18734,17'd18735,17'd18361,17'd18736,17'd18963,17'd18964,17'd18737,17'd15593,17'd16362,17'd18965,17'd18966,17'd18848,17'd17057,17'd18967,17'd18968,17'd18969,17'd17775,17'd16951,17'd17280,17'd17282,17'd15604,17'd15852,17'd16118,17'd16246,17'd16370,17'd17407,17'd17778,17'd17653,17'd17530,17'd17532,17'd15852,17'd15604,17'd17534,17'd18133,17'd16121,17'd16247,17'd18741,17'd18741,17'd18970,17'd18971,17'd12163,17'd18972,17'd18502,17'd18973,17'd18974,17'd18975,17'd18265,17'd18379,17'd18976,17'd18505,17'd18977,17'd12314,17'd18978,17'd11584,17'd18979,17'd18980,17'd6081,17'd18981,17'd18982,17'd18983,17'd18984,17'd957,17'd17423,17'd186,17'd646,17'd18985,17'd12915,17'd18986,17'd3718,17'd4405,17'd4404,17'd4407,17'd7516,17'd8170,17'd8795,17'd10076,17'd10076,17'd11722,17'd11593,17'd12487,17'd9110,17'd11723,17'd11329,17'd11329,17'd15238,17'd15238,17'd16384,17'd18987,17'd16961,17'd18988,17'd18988,17'd16625,17'd16742,17'd17295,17'd15108,17'd18989,17'd18634,17'd17183,17'd18634,17'd18634,17'd8325,17'd16260,17'd18869,17'd18990,17'd12323,17'd11196,17'd11196,17'd11333,17'd9957,17'd10081,17'd16002,17'd12779,17'd8035,17'd2585,17'd271,17'd268,17'd266,17'd265
},
'{
17'd7372,17'd7214,17'd7711,17'd7711,17'd2422,17'd1688,17'd1127,17'd15,17'd1412,17'd283,17'd1275,17'd806,17'd2423,17'd2423,17'd806,17'd2591,17'd8,17'd6,17'd5205,17'd5205,17'd8040,17'd8040,17'd8338,17'd8338,17'd8338,17'd8338,17'd8040,17'd8040,17'd5205,17'd3753,17'd3753,17'd3753,17'd24,17'd24,17'd24,17'd24,17'd23,17'd4,17'd4,17'd4,17'd23,17'd23,17'd1691,17'd285,17'd286,17'd28,17'd4091,17'd3255,17'd2264,17'd1558,17'd18991,17'd2791,17'd491,17'd18992,17'd18993,17'd18994,17'd18995,17'd18996,17'd18997,17'd18876,17'd18283,17'd18998,17'd18999,17'd19000,17'd18769,17'd16273,17'd19001,17'd13446,17'd19002,17'd18882,17'd18883,17'd19003,17'd15894,17'd18772,17'd19004,17'd18528,17'd17094,17'd18773,17'd16651,17'd18408,17'd18531,17'd19005,17'd18173,17'd14622,17'd16163,17'd16163,17'd13969,17'd13840,17'd15137,17'd12529,17'd12679,17'd12679,17'd13093,17'd12955,17'd14764,17'd12361,17'd19006,17'd19007,17'd17206,17'd19008,17'd17445,17'd17320,17'd15524,17'd15769,17'd19009,17'd18776,17'd19010,17'd19011,17'd19012,17'd19013,17'd19014,17'd19015,17'd19016,17'd18892,17'd18782,17'd16036,17'd16992,17'd16886,17'd19017,17'd19018,17'd19019,17'd19020,17'd9707,17'd14109,17'd9310,17'd9310,17'd11095,17'd9311,17'd19021,17'd19022,17'd9445,17'd9311,17'd17947,17'd17702,17'd17333,17'd18426,17'd18311,17'd18898,17'd18898,17'd18898,17'd18069,17'd19023,17'd18790,17'd19024,17'd19025,17'd18312,17'd19026,17'd19027,17'd19028,17'd18672,17'd19029,17'd15929,17'd12984,17'd14661,17'd14124,17'd14662,17'd14372,17'd11934,17'd12704,17'd12397,17'd12236,17'd13638,17'd12403,17'd18801,17'd12715,17'd19030,17'd13882,17'd17125,17'd10991,17'd16683,17'd9885,17'd17599,17'd10479,17'd17719,17'd10479,17'd14518,17'd16320,17'd10737,17'd11395,17'd12861,17'd11960,17'd11959,17'd14807,17'd12253,17'd12253,17'd14807,17'd12106,17'd17967,17'd12582,17'd12582,17'd16204,17'd16204,17'd12582,17'd18917,17'd15053,17'd12996,17'd12422,17'd17968,17'd17968,17'd12115,17'd12422,17'd12719,17'd12856,17'd13884,17'd16915,17'd17475,17'd19031,17'd19031,17'd17235,17'd15571,17'd16327,17'd16558,17'd19032,17'd16443,17'd12720,17'd9740,17'd19033,17'd8247,17'd9888,17'd8734,17'd19034,17'd19035,17'd19036,17'd15442,17'd19037,17'd19038,17'd8739,17'd19039,17'd17854,17'd19040,17'd19041,17'd19042,17'd11819,17'd11150,17'd19043,17'd7979,17'd1197,17'd130,17'd132,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd357,17'd19044,17'd19045,17'd19046,17'd19047,17'd19048,17'd19049,17'd19050,17'd19051,17'd19052,17'd18586,17'd19053,17'd19054,17'd19055,17'd19056,17'd19057,17'd19058,17'd19059,17'd19060,17'd18716,17'd19061,17'd19062,17'd19063,17'd19062,17'd19064,17'd19065,17'd18951,17'd9643,17'd18357,17'd19066,17'd15840,17'd17387,17'd18113,17'd19067,17'd17160,17'd18117,17'd18839,17'd19068,17'd18486,17'd17401,17'd16111,17'd16236,17'd17274,17'd18841,17'd19069,17'd18958,17'd19070,17'd19071,17'd19072,17'd19070,17'd19073,17'd19074,17'd19074,17'd19074,17'd19073,17'd19075,17'd18732,17'd18733,17'd18733,17'd18733,17'd18732,17'd18732,17'd18732,17'd18732,17'd18732,17'd18959,17'd18959,17'd18959,17'd18960,17'd18732,17'd18958,17'd18612,17'd18612,17'd18961,17'd18961,17'd18962,17'd19076,17'd19077,17'd18841,17'd19078,17'd15843,17'd19079,17'd14964,17'd19080,17'd16363,17'd16836,17'd18966,17'd19081,17'd19082,17'd19083,17'd19084,17'd19085,17'd16367,17'd17280,17'd19086,17'd15093,17'd15852,17'd15604,17'd15852,17'd16246,17'd17171,17'd17531,17'd17531,17'd17531,17'd17530,17'd16118,17'd15852,17'd18132,17'd17654,17'd16247,17'd16247,17'd18741,17'd18741,17'd19087,17'd19088,17'd14051,17'd19089,17'd19090,17'd19091,17'd19092,17'd15480,17'd19093,17'd18379,17'd17658,17'd18505,17'd19094,17'd19095,17'd19096,17'd19097,17'd19098,17'd5350,17'd6719,17'd3217,17'd19099,17'd19100,17'd19101,17'd18867,17'd1398,17'd19102,17'd255,17'd190,17'd2921,17'd19103,17'd13422,17'd19104,17'd4404,17'd4062,17'd7343,17'd14983,17'd8491,17'd8795,17'd10076,17'd12018,17'd10391,17'd11593,17'd9110,17'd9110,17'd11329,17'd11329,17'd15238,17'd15623,17'd16493,17'd16961,17'd16961,17'd16625,17'd18988,17'd16625,17'd16742,17'd17548,17'd15108,17'd19105,17'd18634,17'd17183,17'd18634,17'd18634,17'd8325,17'd16260,17'd19106,17'd18990,17'd19107,17'd11196,17'd10910,17'd11333,17'd10393,17'd10081,17'd12779,17'd13427,17'd19108,17'd3742,17'd426,17'd207,17'd262,17'd265
},
'{
17'd5508,17'd7545,17'd3250,17'd3250,17'd1831,17'd1688,17'd14,17'd0,17'd283,17'd3,17'd806,17'd806,17'd16747,17'd16747,17'd2933,17'd2421,17'd6,17'd5205,17'd5205,17'd5205,17'd8040,17'd8040,17'd8338,17'd8338,17'd8338,17'd8338,17'd8040,17'd8040,17'd3753,17'd3753,17'd5,17'd5,17'd24,17'd24,17'd24,17'd24,17'd24,17'd5,17'd5,17'd5,17'd5,17'd23,17'd1691,17'd467,17'd7061,17'd6744,17'd4091,17'd3434,17'd1974,17'd1136,17'd481,17'd69,17'd19109,17'd19110,17'd19111,17'd19112,17'd1996,17'd19113,17'd19114,17'd4108,17'd19115,17'd15124,17'd19116,17'd19117,17'd19118,17'd19119,17'd18881,17'd19120,17'd19002,17'd19121,17'd13590,17'd14203,17'd17933,17'd19004,17'd17199,17'd19122,17'd19123,17'd18773,17'd19124,17'd18170,17'd19125,17'd14621,17'd14622,17'd15764,17'd16163,17'd16658,17'd13969,17'd12530,17'd12529,17'd19126,17'd19127,17'd19127,17'd12528,17'd14621,17'd12361,17'd16658,17'd19128,17'd19007,17'd18656,17'd17207,17'd17445,17'd17320,17'd18534,17'd17694,17'd19129,17'd19130,17'd19131,17'd19132,17'd19133,17'd19134,17'd19135,17'd19136,17'd19016,17'd18781,17'd16885,17'd15909,17'd16416,17'd16416,17'd19137,17'd19138,17'd18665,17'd19139,17'd9582,17'd9016,17'd9310,17'd9311,17'd9445,17'd9445,17'd19022,17'd19022,17'd11095,17'd9446,17'd17702,17'd17333,17'd19140,17'd19141,17'd18668,17'd18898,17'd18898,17'd18668,17'd18068,17'd19142,17'd17587,17'd19143,17'd19144,17'd19145,17'd19146,17'd19147,17'd19148,17'd19149,17'd19150,17'd18797,17'd12981,17'd14372,17'd14920,17'd13501,17'd19151,17'd16546,17'd11934,17'd12560,17'd13506,17'd12572,17'd19152,17'd19153,17'd19154,17'd12413,17'd17125,17'd16687,17'd12116,17'd10743,17'd11671,17'd19155,17'd10330,17'd10166,17'd10991,17'd19156,17'd10853,17'd19157,17'd12861,17'd12857,17'd12580,17'd12579,17'd12579,17'd12108,17'd12579,17'd17348,17'd18197,17'd18557,17'd18806,17'd16204,17'd19158,17'd19158,17'd18917,17'd18917,17'd18917,17'd16204,17'd12115,17'd17968,17'd17968,17'd17604,17'd12719,17'd12580,17'd12415,17'd17605,17'd17475,17'd17235,17'd17013,17'd17013,17'd17013,17'd15687,17'd18449,17'd16558,17'd19032,17'd15175,17'd10991,17'd9337,17'd19159,17'd13003,17'd8103,17'd8254,17'd15692,17'd13377,17'd18921,17'd14392,17'd17020,17'd7629,17'd18810,17'd19160,17'd19161,17'd19162,17'd19163,17'd19164,17'd19165,17'd19166,17'd12874,17'd17363,17'd133,17'd130,17'd132,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd19167,17'd19168,17'd19169,17'd19170,17'd19171,17'd19172,17'd19173,17'd19174,17'd19175,17'd19176,17'd19177,17'd19178,17'd19179,17'd19180,17'd19181,17'd19182,17'd19183,17'd19184,17'd18591,17'd19185,17'd19186,17'd19062,17'd19187,17'd19188,17'd19189,17'd19190,17'd19191,17'd10887,17'd19192,17'd16826,17'd19193,17'd18231,17'd19067,17'd19194,17'd19195,17'd19196,17'd19197,17'd19198,17'd19199,17'd17402,17'd17773,17'd17773,17'd18735,17'd19200,17'd18732,17'd19201,17'd19202,17'd19202,17'd19201,17'd19203,17'd19203,17'd19204,17'd19205,17'd19205,17'd19206,17'd19206,17'd19207,17'd19208,17'd19208,17'd19208,17'd19075,17'd19073,17'd19075,17'd19075,17'd19208,17'd19209,17'd19074,17'd19074,17'd19073,17'd18957,17'd18733,17'd18958,17'd19210,17'd18961,17'd19211,17'd19212,17'd19212,17'd19213,17'd18014,17'd17274,17'd15716,17'd19214,17'd19214,17'd16480,17'd16362,17'd19215,17'd19216,17'd19217,17'd19218,17'd17033,17'd19219,17'd19220,17'd15984,17'd16369,17'd15091,17'd16610,17'd15723,17'd15723,17'd15852,17'd16246,17'd17171,17'd17407,17'd17531,17'd17531,17'd17532,17'd16846,17'd15604,17'd15603,17'd18133,17'd19221,17'd16121,17'd18134,17'd19087,17'd19222,17'd19223,17'd15478,17'd19224,17'd19225,17'd19226,17'd19227,17'd19228,17'd18748,17'd19229,17'd18750,17'd19230,17'd19231,17'd19232,17'd19233,17'd19234,17'd19235,17'd6080,17'd19236,17'd19237,17'd19238,17'd19239,17'd19240,17'd399,17'd19241,17'd965,17'd641,17'd8316,17'd4230,17'd2401,17'd19242,17'd3575,17'd4232,17'd4872,17'd7684,17'd8018,17'd8491,17'd10076,17'd12018,17'd10391,17'd11593,17'd9110,17'd9110,17'd11329,17'd11329,17'd15238,17'd15866,17'd19243,17'd19243,17'd16741,17'd16741,17'd16625,17'd18988,17'd16742,17'd16626,17'd15489,17'd15489,17'd18989,17'd14437,17'd14437,17'd14437,17'd12920,17'd13938,17'd19106,17'd18990,17'd18990,17'd11196,17'd10910,17'd8504,17'd12643,17'd9957,17'd13427,17'd8658,17'd19108,17'd2585,17'd207,17'd268,17'd459,17'd265
},
'{
17'd5508,17'd7545,17'd3250,17'd3250,17'd1831,17'd1688,17'd14,17'd0,17'd283,17'd3,17'd2423,17'd806,17'd16747,17'd16747,17'd2933,17'd978,17'd6,17'd5205,17'd5205,17'd5205,17'd8040,17'd8040,17'd8338,17'd8338,17'd8338,17'd8040,17'd8040,17'd3753,17'd3753,17'd3594,17'd5,17'd5,17'd24,17'd24,17'd24,17'd24,17'd24,17'd5,17'd5,17'd5,17'd5,17'd4,17'd467,17'd1833,17'd6902,17'd4431,17'd3755,17'd3104,17'd1702,17'd19244,17'd14871,17'd839,17'd19245,17'd18871,17'd19246,17'd19247,17'd19248,17'd2281,17'd19249,17'd18642,17'd18643,17'd18399,17'd19116,17'd18878,17'd19250,17'd17434,17'd13446,17'd19120,17'd19251,17'd13198,17'd19252,17'd17806,17'd17933,17'd19004,17'd19123,17'd19123,17'd19123,17'd16651,17'd19253,17'd18531,17'd19005,17'd14621,17'd14622,17'd15764,17'd16658,17'd16658,17'd13969,17'd12530,17'd12529,17'd19126,17'd19254,17'd19127,17'd12955,17'd12530,17'd16658,17'd18884,17'd18774,17'd17206,17'd19255,17'd17207,17'd17320,17'd16519,17'd18060,17'd19256,17'd19257,17'd19258,17'd19259,17'd19133,17'd19260,17'd19261,17'd19262,17'd19263,17'd19136,17'd18662,17'd18893,17'd15909,17'd16038,17'd16416,17'd19264,17'd19265,17'd19266,17'd19267,17'd9164,17'd16042,17'd18542,17'd9311,17'd9584,17'd9445,17'd19022,17'd9165,17'd10818,17'd18897,17'd17821,17'd17949,17'd19268,17'd19269,17'd18898,17'd19270,17'd18898,17'd18668,17'd18068,17'd17823,17'd16670,17'd14644,17'd12545,17'd19271,17'd18071,17'd19272,17'd19273,17'd18553,17'd19274,17'd14919,17'd14252,17'd13634,17'd13498,17'd13243,17'd13126,17'd12704,17'd12397,17'd12088,17'd12094,17'd19275,17'd19276,17'd19277,17'd15686,17'd15054,17'd11523,17'd19278,17'd9480,17'd19279,17'd19155,17'd19280,17'd19281,17'd19282,17'd10604,17'd10735,17'd18560,17'd11957,17'd12111,17'd12419,17'd14807,17'd12579,17'd12254,17'd12108,17'd14807,17'd17474,17'd18557,17'd18806,17'd12422,17'd16204,17'd19158,17'd15185,17'd18917,17'd18917,17'd16204,17'd12262,17'd18560,17'd18682,17'd12115,17'd17604,17'd12106,17'd12579,17'd16913,17'd17727,17'd17235,17'd17235,17'd17014,17'd17014,17'd17013,17'd15687,17'd16913,17'd19283,17'd19284,17'd13137,17'd9739,17'd19285,17'd19286,17'd13005,17'd7949,17'd12589,17'd19287,17'd19288,17'd17852,17'd15574,17'd14818,17'd17732,17'd18810,17'd8264,17'd19289,17'd18925,17'd19290,17'd19291,17'd15313,17'd19292,17'd10873,17'd16090,17'd1481,17'd721,17'd132,17'd5593,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd19293,17'd19294,17'd19295,17'd19296,17'd19297,17'd19298,17'd19299,17'd19300,17'd19301,17'd19302,17'd19303,17'd19304,17'd19305,17'd19306,17'd19307,17'd19308,17'd19309,17'd19310,17'd19311,17'd18595,17'd19312,17'd19313,17'd19314,17'd19315,17'd19316,17'd19317,17'd19318,17'd19319,17'd19320,17'd19321,17'd19193,17'd19322,17'd19323,17'd19324,17'd19325,17'd19326,17'd19327,17'd18606,17'd19328,17'd17402,17'd19329,17'd18248,17'd19330,17'd19331,17'd19073,17'd19332,17'd19333,17'd19333,17'd19203,17'd19204,17'd19204,17'd19334,17'd19335,17'd19336,17'd19336,17'd19336,17'd19205,17'd19206,17'd19337,17'd19208,17'd19208,17'd19073,17'd19073,17'd19209,17'd19338,17'd19208,17'd19074,17'd19339,17'd19074,17'd19075,17'd18732,17'd18733,17'd19340,17'd19210,17'd18961,17'd19211,17'd19341,17'd19212,17'd19077,17'd18248,17'd17167,17'd15716,17'd19342,17'd19343,17'd19344,17'd18738,17'd19345,17'd19217,17'd13023,17'd19346,17'd14718,17'd11177,17'd15471,17'd16951,17'd19347,17'd15091,17'd15724,17'd15603,17'd15603,17'd15852,17'd17171,17'd17407,17'd17653,17'd17531,17'd17529,17'd16953,17'd15852,17'd15723,17'd17654,17'd18133,17'd16121,17'd16121,17'd18741,17'd19222,17'd18375,17'd13559,17'd19348,17'd17906,17'd19349,17'd19350,17'd19351,17'd19352,17'd18750,17'd19353,17'd19354,17'd19355,17'd4383,17'd4702,17'd19356,17'd19357,17'd19358,17'd19359,17'd19360,17'd19361,17'd19362,17'd788,17'd615,17'd19363,17'd1826,17'd772,17'd3090,17'd3087,17'd1953,17'd19364,17'd3575,17'd4232,17'd4717,17'd7516,17'd14983,17'd8170,17'd9405,17'd10076,17'd10391,17'd10077,17'd10650,17'd9110,17'd11329,17'd11329,17'd15238,17'd15623,17'd16135,17'd19243,17'd16741,17'd16741,17'd16625,17'd18988,17'd16742,17'd16742,17'd15489,17'd19105,17'd18989,17'd14437,17'd18989,17'd14437,17'd12920,17'd19365,17'd19366,17'd18990,17'd18990,17'd11196,17'd10910,17'd8504,17'd16631,17'd10393,17'd8658,17'd8658,17'd7534,17'd2585,17'd207,17'd268,17'd266,17'd459
},
'{
17'd2422,17'd2422,17'd1831,17'd1831,17'd4247,17'd14,17'd1,17'd1412,17'd3,17'd3,17'd2423,17'd16636,17'd16500,17'd2933,17'd4,17'd4,17'd7,17'd5205,17'd8040,17'd8340,17'd8340,17'd8340,17'd8340,17'd8040,17'd8040,17'd8040,17'd8040,17'd5205,17'd3753,17'd6,17'd5,17'd5,17'd24,17'd24,17'd5,17'd5,17'd5,17'd5,17'd5,17'd5,17'd4,17'd23,17'd467,17'd286,17'd18037,17'd3907,17'd4249,17'd2602,17'd1557,17'd827,17'd304,17'd491,17'd18992,17'd19367,17'd17556,17'd19368,17'd2136,17'd19369,17'd18876,17'd18159,17'd19370,17'd19371,17'd19372,17'd19373,17'd19001,17'd19374,17'd19120,17'd19002,17'd13081,17'd19375,17'd19376,17'd19377,17'd19377,17'd18771,17'd19378,17'd19379,17'd19380,17'd19381,17'd18296,17'd19005,17'd14890,17'd12814,17'd12530,17'd13969,17'd16658,17'd16765,17'd14622,17'd14890,17'd12679,17'd19127,17'd19126,17'd19126,17'd12814,17'd12530,17'd16658,17'd19382,17'd18655,17'd18656,17'd19383,17'd19383,17'd16289,17'd19384,17'd19384,17'd16289,17'd19385,17'd16986,17'd19386,17'd19387,17'd19388,17'd19389,17'd19390,17'd19390,17'd18781,17'd14225,17'd19391,17'd16886,17'd16416,17'd18664,17'd19392,17'd19393,17'd19394,17'd9847,17'd13732,17'd18542,17'd11095,17'd9311,17'd9445,17'd9310,17'd11095,17'd10818,17'd18787,17'd17820,17'd18065,17'd19395,17'd19269,17'd19396,17'd19270,17'd18898,17'd18668,17'd19397,17'd18067,17'd19398,17'd15154,17'd19399,17'd12378,17'd19400,17'd19401,17'd19402,17'd18073,17'd19403,17'd19404,17'd19405,17'd15421,17'd14123,17'd19406,17'd15171,17'd19151,17'd17225,17'd12087,17'd13877,17'd12245,17'd18801,17'd18678,17'd12410,17'd13363,17'd11521,17'd12863,17'd17965,17'd11809,17'd16680,17'd11135,17'd11526,17'd11669,17'd10854,17'd10853,17'd14262,17'd12999,17'd12998,17'd13365,17'd12856,17'd12253,17'd18564,17'd12254,17'd19407,17'd19408,17'd19409,17'd19410,17'd19411,17'd16326,17'd15185,17'd15185,17'd15185,17'd16325,17'd16442,17'd12422,17'd12115,17'd18682,17'd18682,17'd19412,17'd12719,17'd12417,17'd12416,17'd15571,17'd17726,17'd17475,17'd17235,17'd16686,17'd13642,17'd19413,17'd16560,17'd17475,17'd19414,17'd15299,17'd14518,17'd19415,17'd19416,17'd19417,17'd19418,17'd12265,17'd15440,17'd10861,17'd13654,17'd19419,17'd8428,17'd8739,17'd11815,17'd19420,17'd19421,17'd18091,17'd19422,17'd19423,17'd17360,17'd19166,17'd18458,17'd17363,17'd133,17'd133,17'd130,17'd132,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd19293,17'd19424,17'd19425,17'd19426,17'd4656,17'd19427,17'd19428,17'd19429,17'd19430,17'd19431,17'd19432,17'd19433,17'd19434,17'd19435,17'd19436,17'd19437,17'd19438,17'd19439,17'd18945,17'd19440,17'd18354,17'd18948,17'd18354,17'd19441,17'd19442,17'd19314,17'd19443,17'd19444,17'd19445,17'd17043,17'd17271,17'd18358,17'd19323,17'd19446,17'd19447,17'd19448,17'd18121,17'd19449,17'd19450,17'd19451,17'd18248,17'd18735,17'd19452,17'd19453,17'd19454,17'd19455,17'd19456,17'd19456,17'd19457,17'd19458,17'd19459,17'd19459,17'd19460,17'd19461,17'd19462,17'd19463,17'd19463,17'd19464,17'd19460,17'd19465,17'd19466,17'd19467,17'd19468,17'd19469,17'd19469,17'd19470,17'd19207,17'd19337,17'd19454,17'd19454,17'd19209,17'd18609,17'd19471,17'd19471,17'd19472,17'd19472,17'd19200,17'd19473,17'd19212,17'd19213,17'd19474,17'd16356,17'd18964,17'd18614,17'd19343,17'd16836,17'd16114,17'd19475,17'd14965,17'd18740,17'd14833,17'd19476,17'd9387,17'd19477,17'd16368,17'd19347,17'd17528,17'd15605,17'd15605,17'd17282,17'd16118,17'd17171,17'd17531,17'd17653,17'd17530,17'd17532,17'd16118,17'd15852,17'd19478,17'd18133,17'd17533,17'd17533,17'd18741,17'd19479,17'd19480,17'd19481,17'd19482,17'd18622,17'd19483,17'd19484,17'd19485,17'd19486,17'd19353,17'd19353,17'd19354,17'd19487,17'd7019,17'd4211,17'd19488,17'd4218,17'd4049,17'd4051,17'd19489,17'd19490,17'd19491,17'd19492,17'd177,17'd178,17'd17185,17'd255,17'd19493,17'd19494,17'd19495,17'd3718,17'd3575,17'd3575,17'd4407,17'd4872,17'd14983,17'd8795,17'd9534,17'd13810,17'd10391,17'd10077,17'd10650,17'd9110,17'd11329,17'd10078,17'd12918,17'd12918,17'd17181,17'd16135,17'd19243,17'd19243,17'd19243,17'd19496,17'd16742,17'd16626,17'd16962,17'd19105,17'd14437,17'd19497,17'd19497,17'd19365,17'd12920,17'd12920,17'd19106,17'd18990,17'd18990,17'd12323,17'd11196,17'd9802,17'd17421,17'd8657,17'd7701,17'd7701,17'd19498,17'd2765,17'd258,17'd257,17'd266,17'd459
},
'{
17'd2422,17'd2422,17'd1831,17'd1831,17'd4247,17'd14,17'd1,17'd1412,17'd3,17'd3,17'd2423,17'd16636,17'd16747,17'd2933,17'd4,17'd6,17'd5205,17'd5205,17'd8040,17'd8340,17'd8340,17'd8340,17'd8340,17'd8040,17'd8040,17'd8040,17'd5205,17'd3753,17'd6,17'd5,17'd5,17'd24,17'd24,17'd5,17'd5,17'd5,17'd5,17'd5,17'd5,17'd5,17'd4,17'd25,17'd286,17'd287,17'd9554,17'd3754,17'd2944,17'd2266,17'd19499,17'd482,17'd19500,17'd19501,17'd18760,17'd19502,17'd19503,17'd1996,17'd19504,17'd19505,17'd19506,17'd18159,17'd19507,17'd19371,17'd18999,17'd19508,17'd19509,17'd13959,17'd19120,17'd16400,17'd16275,17'd13590,17'd14203,17'd15894,17'd15894,17'd17440,17'd14090,17'd17312,17'd19510,17'd18654,17'd18058,17'd12955,17'd12814,17'd12360,17'd12530,17'd13969,17'd12361,17'd12361,17'd14621,17'd12955,17'd12679,17'd19127,17'd19126,17'd12528,17'd12218,17'd11913,17'd19006,17'd17689,17'd19511,17'd18656,17'd18656,17'd18656,17'd16164,17'd19384,17'd16164,17'd17319,17'd19383,17'd16986,17'd19512,17'd19513,17'd19514,17'd19389,17'd19515,17'd19516,17'd19517,17'd14225,17'd16885,17'd16886,17'd15777,17'd19518,17'd19519,17'd19266,17'd10567,17'd9847,17'd19520,17'd18542,17'd19521,17'd9311,17'd9310,17'd11095,17'd19521,17'd10818,17'd18787,17'd19522,17'd19523,17'd19269,17'd19396,17'd19396,17'd19396,17'd18898,17'd18311,17'd18309,17'd17950,17'd19524,17'd19525,17'd19526,17'd10953,17'd18431,17'd19527,17'd18672,17'd16899,17'd19528,17'd12563,17'd13502,17'd14662,17'd14123,17'd15171,17'd13874,17'd12086,17'd15674,17'd18799,17'd12402,17'd19529,17'd18913,17'd19530,17'd15808,17'd11667,17'd11399,17'd9884,17'd9742,17'd19531,17'd16070,17'd10479,17'd19532,17'd11130,17'd19533,17'd13516,17'd13362,17'd12857,17'd13365,17'd12995,17'd13517,17'd12579,17'd12254,17'd12254,17'd19407,17'd18559,17'd18197,17'd18806,17'd18806,17'd16326,17'd15185,17'd15185,17'd15185,17'd16325,17'd19158,17'd12262,17'd12115,17'd18682,17'd17968,17'd18328,17'd11958,17'd12418,17'd19534,17'd16327,17'd17726,17'd17235,17'd15571,17'd13642,17'd13642,17'd16914,17'd15687,17'd16559,17'd19284,17'd13000,17'd9883,17'd9044,17'd19535,17'd8101,17'd12120,17'd15188,17'd10180,17'd19536,17'd19537,17'd14683,17'd7626,17'd13772,17'd19538,17'd19539,17'd15062,17'd19540,17'd19541,17'd14821,17'd10350,17'd19542,17'd13899,17'd16090,17'd133,17'd133,17'd133,17'd132,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd358,17'd3812,17'd19543,17'd18579,17'd19544,17'd19545,17'd19546,17'd19547,17'd19548,17'd19549,17'd19550,17'd19551,17'd19552,17'd19553,17'd19554,17'd19555,17'd19556,17'd19557,17'd19184,17'd19558,17'd19559,17'd19185,17'd19560,17'd18717,17'd19561,17'd19441,17'd19562,17'd19563,17'd19444,17'd17387,17'd17263,17'd19067,17'd19323,17'd19564,17'd19565,17'd19566,17'd18121,17'd19567,17'd18248,17'd19568,17'd19569,17'd19077,17'd19452,17'd19570,17'd19571,17'd19455,17'd19206,17'd19205,17'd19458,17'd19459,17'd19459,17'd19572,17'd19462,17'd19463,17'd19573,17'd19574,17'd19575,17'd19576,17'd19575,17'd19577,17'd19578,17'd19465,17'd19465,17'd19469,17'd19579,17'd19580,17'd19468,17'd19571,17'd19454,17'd19454,17'd19454,17'd19581,17'd19582,17'd19340,17'd19583,17'd19583,17'd19200,17'd19200,17'd19212,17'd19069,17'd19584,17'd19474,17'd18736,17'd19585,17'd19586,17'd19587,17'd15846,17'd15215,17'd13153,17'd14717,17'd19588,17'd14719,17'd19589,17'd15220,17'd15983,17'd16951,17'd17061,17'd15093,17'd15605,17'd15724,17'd15604,17'd16246,17'd17530,17'd17531,17'd17530,17'd17529,17'd16246,17'd16118,17'd19478,17'd17654,17'd19221,17'd19221,17'd16121,17'd19590,17'd18022,17'd19223,17'd14425,17'd19224,17'd19591,17'd19592,17'd19593,17'd19594,17'd19353,17'd19595,17'd19596,17'd4859,17'd4210,17'd4210,17'd6233,17'd19597,17'd19598,17'd4221,17'd19599,17'd19600,17'd19601,17'd19602,17'd177,17'd215,17'd17423,17'd254,17'd19603,17'd19494,17'd19495,17'd13422,17'd3575,17'd3575,17'd4062,17'd4872,17'd14983,17'd8795,17'd8796,17'd9534,17'd10391,17'd10077,17'd10650,17'd9110,17'd11329,17'd10078,17'd12918,17'd12918,17'd17181,17'd17181,17'd16135,17'd19243,17'd19496,17'd19496,17'd16742,17'd18388,17'd19604,17'd19105,17'd19497,17'd19497,17'd19497,17'd19365,17'd12920,17'd19605,17'd19606,17'd18990,17'd18389,17'd19107,17'd11196,17'd9802,17'd17297,17'd7533,17'd7701,17'd8035,17'd19498,17'd19607,17'd256,17'd257,17'd459,17'd459
},
'{
17'd2422,17'd2422,17'd1831,17'd1831,17'd1127,17'd2,17'd3,17'd283,17'd3,17'd3,17'd2423,17'd2423,17'd20,17'd23,17'd6,17'd6,17'd5205,17'd8040,17'd8040,17'd8340,17'd8340,17'd8340,17'd8040,17'd8040,17'd8040,17'd8040,17'd5205,17'd3753,17'd6,17'd5,17'd5,17'd24,17'd5,17'd5,17'd5,17'd5,17'd5,17'd5,17'd5,17'd5,17'd23,17'd21,17'd286,17'd18037,17'd11210,17'd3435,17'd2602,17'd19608,17'd19609,17'd483,17'd19610,17'd19611,17'd19612,17'd19613,17'd19614,17'd19615,17'd19616,17'd19114,17'd16014,17'd18159,17'd18643,17'd19371,17'd18047,17'd19617,17'd19618,17'd19619,17'd19002,17'd13081,17'd16509,17'd16875,17'd14203,17'd15894,17'd17440,17'd14090,17'd14090,17'd17312,17'd18773,17'd18170,17'd19005,17'd12814,17'd12814,17'd12360,17'd12530,17'd13840,17'd12530,17'd12218,17'd13211,17'd13093,17'd13092,17'd13209,17'd12679,17'd12528,17'd12530,17'd11764,17'd19382,17'd18655,17'd19620,17'd19511,17'd18174,17'd17205,17'd11231,17'd11231,17'd17206,17'd19383,17'd18174,17'd16766,17'd19621,17'd19622,17'd19623,17'd19624,17'd19625,17'd19626,17'd19517,17'd18782,17'd16885,17'd19391,17'd19264,17'd19627,17'd19266,17'd10566,17'd10567,17'd9582,17'd9309,17'd11631,17'd11095,17'd9311,17'd9017,17'd9165,17'd10818,17'd10701,17'd18787,17'd19522,17'd19628,17'd19629,17'd19630,17'd19630,17'd19396,17'd18668,17'd18427,17'd17950,17'd19631,17'd19632,17'd19633,17'd12225,17'd17954,17'd18551,17'd19634,17'd19635,17'd19636,17'd19637,17'd13503,17'd19638,17'd13995,17'd14123,17'd15171,17'd12234,17'd12559,17'd14374,17'd19639,17'd18912,17'd14127,17'd19640,17'd19641,17'd18805,17'd16320,17'd16796,17'd16912,17'd10170,17'd11135,17'd19642,17'd11528,17'd19282,17'd11275,17'd19643,17'd16326,17'd13883,17'd12419,17'd12995,17'd12856,17'd12417,17'd12579,17'd12253,17'd16203,17'd19408,17'd18557,17'd18557,17'd12582,17'd12582,17'd12582,17'd12582,17'd18917,17'd18917,17'd15185,17'd16326,17'd12115,17'd17968,17'd19644,17'd18330,17'd14002,17'd12995,17'd12860,17'd16558,17'd17726,17'd17726,17'd15571,17'd15571,17'd14672,17'd14672,17'd15571,17'd14672,17'd19032,17'd19645,17'd10476,17'd10744,17'd11403,17'd14135,17'd7947,17'd9622,17'd10746,17'd14531,17'd19646,17'd19647,17'd19648,17'd8263,17'd15696,17'd11815,17'd19649,17'd19650,17'd16451,17'd19651,17'd19652,17'd19653,17'd19654,17'd19655,17'd16090,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd357,17'd5311,17'd19656,17'd19657,17'd17364,17'd18580,17'd19658,17'd19659,17'd19660,17'd19661,17'd19662,17'd19663,17'd19664,17'd19665,17'd19666,17'd19667,17'd19668,17'd19669,17'd19670,17'd19671,17'd19672,17'd19559,17'd19559,17'd18833,17'd19673,17'd18717,17'd19674,17'd19675,17'd19444,17'd16827,17'd17512,17'd19676,17'd18002,17'd19564,17'd19677,17'd19678,17'd19679,17'd19680,17'd19681,17'd19568,17'd19682,17'd19069,17'd19683,17'd19684,17'd19337,17'd19685,17'd19469,17'd19686,17'd19572,17'd19687,17'd19461,17'd19462,17'd19688,17'd19689,17'd19690,17'd19691,17'd19692,17'd19693,17'd19694,17'd19693,17'd19695,17'd19696,17'd19697,17'd19698,17'd19699,17'd19699,17'd19700,17'd19469,17'd19468,17'd19470,17'd19701,17'd19702,17'd19703,17'd19704,17'd19705,17'd19706,17'd19707,17'd19200,17'd19473,17'd19076,17'd19708,17'd19709,17'd19710,17'd18963,17'd19711,17'd19712,17'd19713,17'd15215,17'd8611,17'd14565,17'd14718,17'd15457,17'd14832,17'd19589,17'd19220,17'd16245,17'd18851,17'd17061,17'd17061,17'd17528,17'd15724,17'd17283,17'd16370,17'd18019,17'd17531,17'd17529,17'd16370,17'd16246,17'd16118,17'd15723,17'd15475,17'd18133,17'd16121,17'd19590,17'd18742,17'd19714,17'd19715,17'd19716,17'd19717,17'd19718,17'd19719,17'd19720,17'd19721,17'd19722,17'd19723,17'd10243,17'd4211,17'd19724,17'd19725,17'd19726,17'd19727,17'd3557,17'd19728,17'd19729,17'd19730,17'd19731,17'd788,17'd215,17'd400,17'd17789,17'd189,17'd19732,17'd19495,17'd1816,17'd4064,17'd4408,17'd4062,17'd4717,17'd7684,17'd8170,17'd8954,17'd9534,17'd9946,17'd10391,17'd10650,17'd9110,17'd11329,17'd10078,17'd12918,17'd12918,17'd12918,17'd17181,17'd17181,17'd17181,17'd17181,17'd17181,17'd16259,17'd16259,17'd12640,17'd12777,17'd10079,17'd9952,17'd9952,17'd9951,17'd8962,17'd8962,17'd4072,17'd19733,17'd19733,17'd19734,17'd19735,17'd8182,17'd17297,17'd7359,17'd7533,17'd7533,17'd9663,17'd2924,17'd1242,17'd801,17'd460,17'd456
},
'{
17'd2422,17'd2422,17'd1831,17'd4247,17'd466,17'd0,17'd3,17'd3,17'd12,17'd12,17'd2423,17'd2423,17'd21,17'd23,17'd6,17'd3753,17'd8040,17'd8040,17'd8040,17'd8340,17'd8340,17'd8340,17'd8040,17'd8040,17'd8040,17'd8040,17'd5205,17'd3753,17'd6,17'd5,17'd24,17'd24,17'd5,17'd5,17'd5,17'd5,17'd5,17'd5,17'd5,17'd5,17'd23,17'd21,17'd27,17'd18037,17'd11210,17'd3258,17'd2263,17'd1557,17'd57,17'd14872,17'd19736,17'd19737,17'd19738,17'd19739,17'd19740,17'd19615,17'd19741,17'd19742,17'd16014,17'd19743,17'd19115,17'd19744,17'd19745,17'd19746,17'd19747,17'd19748,17'd12940,17'd13081,17'd13449,17'd19003,17'd14203,17'd19749,17'd18652,17'd14090,17'd19750,17'd19751,17'd19752,17'd18531,17'd14890,17'd12360,17'd12360,17'd12530,17'd12530,17'd12530,17'd12530,17'd12065,17'd13093,17'd12813,17'd13092,17'd13209,17'd12955,17'd12814,17'd11913,17'd11362,17'd19753,17'd19511,17'd19511,17'd18655,17'd17205,17'd16766,17'd11231,17'd11231,17'd17206,17'd19383,17'd16766,17'd19754,17'd19755,17'd19756,17'd19757,17'd19758,17'd19515,17'd13850,17'd14105,17'd17102,17'd19391,17'd19759,17'd19760,17'd19761,17'd10698,17'd10121,17'd9847,17'd9582,17'd9309,17'd9310,17'd11095,17'd11095,17'd9017,17'd9165,17'd9446,17'd9446,17'd18787,17'd19523,17'd19762,17'd19629,17'd19630,17'd19763,17'd19764,17'd18311,17'd18546,17'd19765,17'd19766,17'd19767,17'd19768,17'd19769,17'd19770,17'd19771,17'd19772,17'd15550,17'd18910,17'd13636,17'd15555,17'd17959,17'd13995,17'd13127,17'd13632,17'd19773,17'd19774,17'd19775,17'd19776,17'd19777,17'd19778,17'd19641,17'd15046,17'd10735,17'd10023,17'd10992,17'd10170,17'd19779,17'd11401,17'd11670,17'd11133,17'd10739,17'd10989,17'd16326,17'd16442,17'd14130,17'd12580,17'd12856,17'd12417,17'd12417,17'd12579,17'd12579,17'd19408,17'd18559,17'd19410,17'd19410,17'd12582,17'd12582,17'd12582,17'd18917,17'd18917,17'd18917,17'd19158,17'd13516,17'd17968,17'd17968,17'd18330,17'd18328,17'd13136,17'd12575,17'd16559,17'd17727,17'd17726,17'd17726,17'd15571,17'd15687,17'd14672,17'd14672,17'd14524,17'd13884,17'd14131,17'd16069,17'd17719,17'd17600,17'd9744,17'd19780,17'd17241,17'd15188,17'd19781,17'd14938,17'd14387,17'd19782,17'd19783,17'd19784,17'd8429,17'd9893,17'd17610,17'd16212,17'd14272,17'd11818,17'd9754,17'd19785,17'd13899,17'd15823,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd10492,17'd19786,17'd19787,17'd19788,17'd19789,17'd19790,17'd19791,17'd19792,17'd19793,17'd19794,17'd19795,17'd19796,17'd19797,17'd19798,17'd19799,17'd19800,17'd19801,17'd19802,17'd19803,17'd19804,17'd19672,17'd19805,17'd19806,17'd19807,17'd18594,17'd19808,17'd19809,17'd19810,17'd19811,17'd17643,17'd19812,17'd17267,17'd19813,17'd19814,17'd19815,17'd19679,17'd19680,17'd19816,17'd19817,17'd19818,17'd19708,17'd19819,17'd19820,17'd19470,17'd19821,17'd19822,17'd19823,17'd19824,17'd19825,17'd19462,17'd19688,17'd19826,17'd19827,17'd19692,17'd19828,17'd19829,17'd19830,17'd19831,17'd19832,17'd19833,17'd19834,17'd19695,17'd19835,17'd19836,17'd19837,17'd19837,17'd19838,17'd19686,17'd19580,17'd19702,17'd19702,17'd19839,17'd19703,17'd19840,17'd19705,17'd19841,17'd19707,17'd19200,17'd19473,17'd19842,17'd19708,17'd19818,17'd19710,17'd15843,17'd19843,17'd19844,17'd15595,17'd9640,17'd8148,17'd14551,17'd14719,17'd14832,17'd14832,17'd19845,17'd15471,17'd19846,17'd19086,17'd17061,17'd17061,17'd15093,17'd15724,17'd16118,17'd17171,17'd17531,17'd17530,17'd18019,17'd17171,17'd16246,17'd15604,17'd15603,17'd16119,17'd16121,17'd15988,17'd18260,17'd19847,17'd19848,17'd19849,17'd19850,17'd19851,17'd19852,17'd19853,17'd19854,17'd19722,17'd19855,17'd19856,17'd19857,17'd4211,17'd19858,17'd7679,17'd19859,17'd19860,17'd19861,17'd19862,17'd19863,17'd763,17'd788,17'd19864,17'd17186,17'd15626,17'd2588,17'd19865,17'd8016,17'd1388,17'd4064,17'd4064,17'd4062,17'd4717,17'd7516,17'd8170,17'd8954,17'd8796,17'd9946,17'd10391,17'd9254,17'd9110,17'd11329,17'd11329,17'd12918,17'd12918,17'd12918,17'd12918,17'd12918,17'd17181,17'd17181,17'd17181,17'd17181,17'd12776,17'd19866,17'd9795,17'd19867,17'd9952,17'd9952,17'd9951,17'd8962,17'd8649,17'd19868,17'd19869,17'd19733,17'd19869,17'd19870,17'd19871,17'd17184,17'd17421,17'd7533,17'd19872,17'd4078,17'd19873,17'd255,17'd801,17'd456,17'd456
},
'{
17'd3250,17'd2422,17'd1831,17'd4247,17'd2,17'd12,17'd806,17'd806,17'd2423,17'd2423,17'd2423,17'd8814,17'd23,17'd4,17'd6,17'd5205,17'd8040,17'd8040,17'd8340,17'd8340,17'd8340,17'd8040,17'd8040,17'd8040,17'd8040,17'd8040,17'd3753,17'd3753,17'd5,17'd5,17'd24,17'd24,17'd7383,17'd7383,17'd5,17'd5,17'd5,17'd5,17'd5,17'd5,17'd23,17'd285,17'd6744,17'd9554,17'd12335,17'd3105,17'd19874,17'd1135,17'd61,17'd69,17'd19875,17'd19876,17'd19877,17'd19878,17'd19879,17'd19880,17'd19881,17'd19882,17'd19883,17'd19884,17'd19885,17'd15251,17'd19886,17'd19887,17'd12939,17'd19888,17'd13197,17'd16275,17'd16649,17'd15128,17'd19889,17'd17566,17'd14883,17'd19750,17'd19751,17'd19124,17'd18170,17'd18532,17'd19890,17'd15137,17'd12530,17'd12530,17'd12530,17'd12530,17'd14890,17'd12528,17'd13092,17'd13092,17'd13599,17'd13599,17'd13211,17'd12362,17'd12532,17'd17941,17'd18174,17'd19891,17'd18774,17'd19892,17'd17689,17'd19893,17'd16766,17'd18174,17'd18656,17'd18656,17'd19893,17'd19512,17'd7746,17'd19894,17'd19389,17'd19758,17'd19895,17'd19896,17'd19897,17'd14632,17'd19759,17'd13975,17'd19898,17'd19899,17'd10698,17'd9989,17'd19900,17'd13732,17'd11631,17'd9310,17'd9017,17'd9017,17'd9165,17'd9165,17'd18307,17'd19901,17'd19902,17'd19903,17'd19762,17'd19904,17'd19905,17'd19906,17'd19907,17'd18310,17'd18546,17'd19631,17'd15919,17'd19908,17'd19909,17'd19910,17'd19911,17'd19912,17'd16054,17'd14510,17'd14373,17'd19913,17'd17959,17'd13129,17'd13501,17'd12393,17'd19773,17'd15675,17'd19914,17'd12098,17'd19915,17'd19916,17'd19530,17'd18804,17'd19917,17'd10325,17'd19918,17'd9885,17'd19779,17'd19919,17'd11400,17'd19532,17'd10855,17'd10852,17'd14262,17'd12996,17'd19920,17'd15184,17'd12995,17'd14809,17'd12418,17'd12418,17'd12253,17'd14807,17'd18198,17'd18557,17'd19921,17'd18681,17'd19158,17'd15185,17'd18917,17'd18917,17'd18197,17'd18917,17'd11964,17'd13516,17'd19922,17'd17968,17'd18328,17'd12719,17'd12856,17'd12997,17'd14524,17'd17235,17'd15571,17'd15571,17'd15687,17'd15687,17'd12860,17'd12860,17'd12860,17'd13644,17'd15175,17'd10991,17'd9346,17'd12118,17'd19923,17'd17128,17'd10860,17'd10180,17'd10747,17'd12429,17'd19924,17'd15306,17'd19784,17'd19925,17'd12593,17'd19926,17'd18092,17'd19927,17'd18094,17'd19928,17'd19929,17'd19930,17'd10874,17'd131,17'd131,17'd132,17'd133,17'd133,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd2861,17'd6691,17'd19931,17'd19932,17'd19933,17'd19934,17'd19935,17'd19936,17'd19937,17'd19938,17'd19939,17'd19940,17'd19941,17'd19942,17'd19943,17'd19944,17'd19945,17'd19946,17'd19947,17'd19948,17'd19949,17'd19950,17'd18947,17'd19951,17'd18947,17'd19808,17'd19809,17'd19810,17'd17642,17'd19952,17'd19953,17'd18483,17'd19954,17'd19677,17'd19565,17'd18121,17'd19955,17'd18735,17'd19817,17'd19708,17'd19200,17'd19956,17'd19957,17'd19821,17'd19578,17'd19700,17'd19699,17'd19463,17'd19463,17'd19688,17'd19826,17'd19958,17'd19959,17'd19960,17'd19961,17'd19962,17'd19963,17'd19964,17'd19965,17'd19965,17'd19966,17'd19967,17'd19968,17'd19969,17'd19969,17'd19969,17'd19970,17'd19971,17'd19837,17'd19700,17'd19972,17'd19701,17'd19973,17'd19974,17'd19453,17'd19975,17'd19841,17'd19707,17'd19707,17'd19473,17'd19976,17'd19708,17'd19709,17'd19977,17'd15716,17'd19978,17'd19979,17'd15210,17'd14716,17'd13544,17'd14718,17'd14952,17'd19980,17'd19981,17'd19982,17'd19983,17'd19984,17'd17060,17'd17061,17'd14570,17'd15093,17'd15604,17'd16246,17'd18019,17'd17407,17'd17407,17'd17171,17'd16370,17'd15852,17'd17282,17'd15605,17'd19221,17'd16121,17'd18260,17'd19985,17'd19986,17'd19987,17'd19988,17'd19989,17'd19990,17'd19991,17'd19992,17'd19722,17'd19721,17'd19596,17'd19232,17'd4701,17'd7844,17'd7508,17'd19993,17'd19994,17'd19995,17'd19996,17'd19997,17'd19998,17'd19999,17'd20000,17'd20001,17'd213,17'd255,17'd20002,17'd20003,17'd2106,17'd4064,17'd4064,17'd7031,17'd7193,17'd7346,17'd7856,17'd9252,17'd8796,17'd8955,17'd10526,17'd9255,17'd9110,17'd11329,17'd18146,17'd12918,17'd12918,17'd20004,17'd12918,17'd12776,17'd12776,17'd17181,17'd17181,17'd12918,17'd12776,17'd19866,17'd11192,17'd20005,17'd10079,17'd9952,17'd9951,17'd9951,17'd8649,17'd4412,17'd3726,17'd20006,17'd20006,17'd20007,17'd4874,17'd19498,17'd19498,17'd19872,17'd19872,17'd5786,17'd1239,17'd20008,17'd403,17'd20009,17'd20009
},
'{
17'd3250,17'd2422,17'd1831,17'd4247,17'd2,17'd3,17'd806,17'd806,17'd806,17'd2423,17'd2423,17'd2933,17'd23,17'd5,17'd3753,17'd5205,17'd8040,17'd8340,17'd8340,17'd8340,17'd8040,17'd8040,17'd8040,17'd8040,17'd8040,17'd8040,17'd3753,17'd3753,17'd5,17'd5,17'd24,17'd24,17'd7383,17'd7383,17'd5,17'd5,17'd5,17'd5,17'd5,17'd5,17'd23,17'd285,17'd6744,17'd3907,17'd12335,17'd2264,17'd1839,17'd991,17'd65,17'd840,17'd20010,17'd20011,17'd17667,17'd20012,17'd19879,17'd19880,17'd20013,17'd20014,17'd20015,17'd20016,17'd20017,17'd20018,17'd20019,17'd20020,17'd12664,17'd19888,17'd13197,17'd16275,17'd16649,17'd15128,17'd16875,17'd13963,17'd14883,17'd19750,17'd20021,17'd20022,17'd18058,17'd15383,17'd18411,17'd14891,17'd13969,17'd12361,17'd12530,17'd12814,17'd12528,17'd12679,17'd13092,17'd13092,17'd13599,17'd17809,17'd14470,17'd16765,17'd19006,17'd18533,17'd20023,17'd18174,17'd17689,17'd19128,17'd19893,17'd19893,17'd17205,17'd19891,17'd18656,17'd18656,17'd17689,17'd19387,17'd20024,17'd20025,17'd20026,17'd20027,17'd20028,17'd20029,17'd14632,17'd20030,17'd13975,17'd20031,17'd13330,17'd20032,17'd10698,17'd9847,17'd19900,17'd9309,17'd11631,17'd9310,17'd9017,17'd9017,17'd9165,17'd9018,17'd18307,17'd20033,17'd19523,17'd20034,17'd20035,17'd19904,17'd19906,17'd20036,17'd18311,17'd18546,17'd20037,17'd20038,17'd20039,17'd11367,17'd20040,17'd10301,17'd20041,17'd20042,17'd18797,17'd15420,17'd17959,17'd20043,17'd17959,17'd13130,17'd14253,17'd12235,17'd12559,17'd13506,17'd18800,17'd11796,17'd19276,17'd12992,17'd12574,17'd12718,17'd10735,17'd20044,17'd9341,17'd12116,17'd20045,17'd20046,17'd11525,17'd14263,17'd10738,17'd10736,17'd15186,17'd12861,17'd18565,17'd15184,17'd12417,17'd13643,17'd12418,17'd12418,17'd12579,17'd19408,17'd18197,17'd20047,17'd18681,17'd18681,17'd19158,17'd15185,17'd18917,17'd18917,17'd18557,17'd12582,17'd11964,17'd11965,17'd17968,17'd12422,17'd12719,17'd16321,17'd12418,17'd12860,17'd15571,17'd15571,17'd15571,17'd15687,17'd15687,17'd15811,17'd12860,17'd12860,17'd12418,17'd14131,17'd12720,17'd9473,17'd11402,17'd8573,17'd19780,17'd8734,17'd20048,17'd19781,17'd15442,17'd20049,17'd20050,17'd18922,17'd20051,17'd13142,17'd20052,17'd20053,17'd19040,17'd20054,17'd20055,17'd20056,17'd20057,17'd20058,17'd16090,17'd132,17'd132,17'd132,17'd131,17'd133,17'd130,17'd136,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd3168,17'd2866,17'd20059,17'd20060,17'd19296,17'd20061,17'd20062,17'd20063,17'd20064,17'd20065,17'd20066,17'd20067,17'd20068,17'd20069,17'd20070,17'd20071,17'd20072,17'd20073,17'd20074,17'd20075,17'd20076,17'd20077,17'd19807,17'd20078,17'd19807,17'd20079,17'd19317,17'd19810,17'd20080,17'd20081,17'd20082,17'd20083,17'd20084,17'd20085,17'd19565,17'd18241,17'd18846,17'd19077,17'd19077,17'd19212,17'd19331,17'd20086,17'd20087,17'd19824,17'd19699,17'd20088,17'd20089,17'd20090,17'd19573,17'd19689,17'd19827,17'd19959,17'd20091,17'd20092,17'd20093,17'd20094,17'd20094,17'd20095,17'd20096,17'd20097,17'd20098,17'd19966,17'd20099,17'd20100,17'd20101,17'd20102,17'd20102,17'd19971,17'd19971,17'd19823,17'd19822,17'd20103,17'd19702,17'd19973,17'd19974,17'd20104,17'd19975,17'd20105,17'd20105,17'd19331,17'd20106,17'd18962,17'd19069,17'd19817,17'd18727,17'd20107,17'd18965,17'd17056,17'd20108,17'd9372,17'd20109,17'd15456,17'd20110,17'd20111,17'd20112,17'd20113,17'd20114,17'd18851,17'd17060,17'd19086,17'd15093,17'd15603,17'd15852,17'd16370,17'd18019,17'd18019,17'd18019,17'd16370,17'd16118,17'd17283,17'd15724,17'd18133,17'd17533,17'd18134,17'd18742,17'd20115,17'd19715,17'd20116,17'd20117,17'd11857,17'd20118,17'd20119,17'd19486,17'd20120,17'd20121,17'd11438,17'd5768,17'd6400,17'd20122,17'd7846,17'd20123,17'd20124,17'd20125,17'd20126,17'd20127,17'd763,17'd765,17'd434,17'd251,17'd2115,17'd19493,17'd3580,17'd1954,17'd4720,17'd4064,17'd7031,17'd6243,17'd6724,17'd7856,17'd9252,17'd9534,17'd8955,17'd9946,17'd9254,17'd11051,17'd18146,17'd18146,17'd12918,17'd12918,17'd20004,17'd18146,17'd12776,17'd12776,17'd12776,17'd17181,17'd12918,17'd12776,17'd19866,17'd9948,17'd20128,17'd10079,17'd9952,17'd9952,17'd9951,17'd8649,17'd4411,17'd3726,17'd20007,17'd20006,17'd20006,17'd5186,17'd4236,17'd19498,17'd19872,17'd6412,17'd4877,17'd2108,17'd1094,17'd17551,17'd278,17'd278
},
'{
17'd3250,17'd1831,17'd2594,17'd2595,17'd13,17'd3,17'd806,17'd806,17'd806,17'd16636,17'd2423,17'd2933,17'd4,17'd6,17'd3753,17'd8040,17'd8040,17'd8340,17'd8340,17'd8340,17'd8040,17'd8040,17'd8040,17'd8040,17'd8040,17'd5793,17'd3753,17'd3753,17'd3594,17'd3594,17'd24,17'd24,17'd7554,17'd7383,17'd5,17'd5,17'd5,17'd5,17'd5,17'd5,17'd1832,17'd27,17'd4430,17'd3755,17'd3258,17'd2122,17'd1282,17'd666,17'd20129,17'd843,17'd20130,17'd20131,17'd20132,17'd20012,17'd20133,17'd20134,17'd20135,17'd20136,17'd18876,17'd20137,17'd20138,17'd20139,17'd20140,17'd20141,17'd20142,17'd20143,17'd18882,17'd16275,17'd16649,17'd16649,17'd20144,17'd20145,17'd14883,17'd16876,17'd19752,17'd20146,17'd19005,17'd18411,17'd18411,17'd20147,17'd15764,17'd14622,17'd14621,17'd12955,17'd13209,17'd14469,17'd14469,17'd13092,17'd13599,17'd19005,17'd14470,17'd16658,17'd19382,17'd18774,17'd17205,17'd17205,17'd19893,17'd20148,17'd19893,17'd19893,17'd17206,17'd20149,17'd20149,17'd18656,17'd17689,17'd20150,17'd20151,17'd20152,17'd20153,17'd20154,17'd20155,17'd14775,17'd20030,17'd20156,17'd20157,17'd20158,17'd20159,17'd13096,17'd10698,17'd9847,17'd13732,17'd11631,17'd9309,17'd9309,17'd14109,17'd9017,17'd9018,17'd9311,17'd10126,17'd20160,17'd20161,17'd20162,17'd20035,17'd19904,17'd19906,17'd20163,17'd18310,17'd20164,17'd17950,17'd19766,17'd20165,17'd19909,17'd18431,17'd18671,17'd20166,17'd20167,17'd20168,17'd12242,17'd20169,17'd20169,17'd12709,17'd14513,17'd17225,17'd12235,17'd13996,17'd20170,17'd19776,17'd20171,17'd20172,17'd20173,17'd13365,17'd12996,17'd10472,17'd20174,17'd9885,17'd17469,17'd19155,17'd13647,17'd11669,17'd11130,17'd14262,17'd16797,17'd17598,17'd18679,17'd15183,17'd14130,17'd12253,17'd12418,17'd12418,17'd12417,17'd16321,17'd18198,17'd12582,17'd19921,17'd19158,17'd19158,17'd19158,17'd15185,17'd15053,17'd15053,17'd18557,17'd18806,17'd13516,17'd11965,17'd17968,17'd16204,17'd12420,17'd12109,17'd12859,17'd16559,17'd15571,17'd15571,17'd15687,17'd15687,17'd19534,17'd19534,17'd19534,17'd12860,17'd12579,17'd11806,17'd10472,17'd20175,17'd20176,17'd8578,17'd17352,17'd20177,17'd20178,17'd15436,17'd20179,17'd20180,17'd20181,17'd10483,17'd14394,17'd14534,17'd20182,17'd20183,17'd20184,17'd20185,17'd20186,17'd20187,17'd16577,17'd20188,17'd133,17'd130,17'd130,17'd132,17'd131,17'd132,17'd136,17'd136,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd135,17'd20189,17'd20190,17'd18817,17'd20191,17'd19047,17'd20192,17'd20193,17'd20194,17'd20195,17'd20196,17'd20197,17'd20198,17'd20199,17'd20200,17'd20201,17'd20202,17'd20203,17'd20204,17'd20205,17'd20206,17'd20207,17'd19807,17'd20207,17'd19951,17'd20208,17'd19674,17'd20209,17'd20210,17'd20211,17'd20212,17'd20213,17'd20214,17'd19325,17'd20215,17'd20216,17'd19210,17'd19069,17'd19069,17'd19200,17'd20217,17'd20218,17'd19700,17'd19837,17'd20090,17'd20219,17'd20219,17'd20220,17'd20221,17'd19827,17'd20222,17'd20091,17'd20223,17'd20224,17'd20225,17'd20226,17'd20226,17'd20227,17'd20228,17'd20229,17'd20229,17'd20230,17'd20231,17'd20232,17'd20233,17'd19695,17'd20234,17'd20102,17'd20102,17'd19971,17'd19838,17'd20235,17'd20236,17'd20237,17'd20238,17'd20239,17'd20086,17'd20240,17'd19975,17'd19975,17'd19331,17'd19473,17'd19708,17'd19709,17'd20241,17'd20242,17'd20243,17'd19345,17'd20244,17'd8609,17'd20245,17'd20246,17'd20247,17'd19982,17'd20112,17'd20248,17'd20249,17'd19984,17'd18851,17'd19086,17'd14570,17'd15475,17'd15603,17'd15852,17'd16370,17'd18019,17'd17171,17'd16370,17'd16246,17'd16843,17'd17282,17'd15475,17'd19221,17'd18741,17'd20250,17'd20251,17'd20252,17'd20253,17'd20254,17'd20255,17'd12311,17'd20256,17'd20257,17'd19353,17'd19722,17'd20258,17'd5174,17'd6861,17'd20259,17'd20260,17'd3371,17'd20261,17'd20262,17'd19862,17'd20263,17'd20264,17'd20265,17'd20266,17'd613,17'd1682,17'd10073,17'd3410,17'd19495,17'd4064,17'd4064,17'd7031,17'd6243,17'd6576,17'd8169,17'd9252,17'd9534,17'd8797,17'd8798,17'd9255,17'd11051,17'd18146,17'd18146,17'd12918,17'd12918,17'd20004,17'd18146,17'd19866,17'd12640,17'd12776,17'd12918,17'd12918,17'd12776,17'd9948,17'd9948,17'd20128,17'd19867,17'd9952,17'd9952,17'd9951,17'd12179,17'd4412,17'd3726,17'd7522,17'd3881,17'd8025,17'd20267,17'd20268,17'd20269,17'd6412,17'd6412,17'd4877,17'd20270,17'd1095,17'd1095,17'd181,17'd20271
},
'{
17'd3250,17'd1831,17'd2594,17'd466,17'd12,17'd3,17'd806,17'd806,17'd806,17'd16636,17'd2423,17'd2933,17'd8,17'd3753,17'd5793,17'd8040,17'd8040,17'd8340,17'd8340,17'd8340,17'd8040,17'd8040,17'd8040,17'd8040,17'd5793,17'd3753,17'd3753,17'd3594,17'd3594,17'd5,17'd24,17'd24,17'd7554,17'd7554,17'd5,17'd5,17'd5,17'd5,17'd5,17'd4,17'd285,17'd27,17'd4430,17'd3255,17'd3105,17'd1702,17'd1134,17'd58,17'd20272,17'd493,17'd20273,17'd20274,17'd20275,17'd20276,17'd20277,17'd20278,17'd20279,17'd20280,17'd20281,17'd20282,17'd4909,17'd20283,17'd20284,17'd20285,17'd19888,17'd13197,17'd20286,17'd20287,17'd16649,17'd16649,17'd13589,17'd20288,17'd20289,17'd20290,17'd20291,17'd17939,17'd14621,17'd14764,17'd14622,17'd14622,17'd15764,17'd14622,17'd14890,17'd12679,17'd14469,17'd14469,17'd14469,17'd13092,17'd12955,17'd13211,17'd16765,17'd20292,17'd19382,17'd18774,17'd17205,17'd16766,17'd17689,17'd20148,17'd19893,17'd19754,17'd17206,17'd20293,17'd20293,17'd19383,17'd16986,17'd8214,17'd20294,17'd20295,17'd20153,17'd20296,17'd18661,17'd14775,17'd19759,17'd20297,17'd20031,17'd13330,17'd13096,17'd11916,17'd9988,17'd9581,17'd9309,17'd11631,17'd9309,17'd9309,17'd14109,17'd14109,17'd19022,17'd9584,17'd18423,17'd20298,17'd20162,17'd20299,17'd20299,17'd20035,17'd19764,17'd19907,17'd20164,17'd17950,17'd20300,17'd20301,17'd10573,17'd20302,17'd18793,17'd20303,17'd18796,17'd11109,17'd20304,17'd20305,17'd20306,17'd20307,17'd13995,17'd14513,17'd20308,17'd12087,17'd20309,17'd20310,17'd11657,17'd19916,17'd20311,17'd12856,17'd13883,17'd11275,17'd10327,17'd18916,17'd9884,17'd19155,17'd20312,17'd11525,17'd11130,17'd11129,17'd11963,17'd12861,17'd20313,17'd16322,17'd16443,17'd11959,17'd12859,17'd12859,17'd12418,17'd14807,17'd20314,17'd17722,17'd18443,17'd18444,17'd15185,17'd19158,17'd19158,17'd12996,17'd15053,17'd15053,17'd18557,17'd19921,17'd10989,17'd11965,17'd17604,17'd12581,17'd12580,17'd12418,17'd12415,17'd14672,17'd14524,17'd14524,17'd15687,17'd16913,17'd19534,17'd19534,17'd12415,17'd15434,17'd13882,17'd14673,17'd9473,17'd20315,17'd19535,17'd9484,17'd8734,17'd20316,17'd20317,17'd20318,17'd20319,17'd20320,17'd14271,17'd7629,17'd7629,17'd20321,17'd20322,17'd20323,17'd20324,17'd20325,17'd20326,17'd20327,17'd20328,17'd13901,17'd16090,17'd134,17'd134,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd133,17'd134,17'd6531,17'd14146,17'd20329,17'd3030,17'd20330,17'd20331,17'd20332,17'd20333,17'd20334,17'd20335,17'd20336,17'd20337,17'd20338,17'd20339,17'd20340,17'd20341,17'd20342,17'd20343,17'd20344,17'd20345,17'd20346,17'd19951,17'd20346,17'd20347,17'd20208,17'd20348,17'd20349,17'd19674,17'd20350,17'd20351,17'd18359,17'd20352,17'd19325,17'd20353,17'd20354,17'd18610,17'd19473,17'd18962,17'd19707,17'd19841,17'd20238,17'd20355,17'd20102,17'd20102,17'd19970,17'd20356,17'd20221,17'd19827,17'd20357,17'd20358,17'd20223,17'd20359,17'd20360,17'd20361,17'd20362,17'd20227,17'd20363,17'd20364,17'd20365,17'd20365,17'd20366,17'd20367,17'd20230,17'd19966,17'd20368,17'd20100,17'd20369,17'd20101,17'd20370,17'd20371,17'd19838,17'd20235,17'd20236,17'd20237,17'd20238,17'd20239,17'd20372,17'd20240,17'd19975,17'd19706,17'd19707,17'd20373,17'd20374,17'd20375,17'd20376,17'd20377,17'd20378,17'd20379,17'd20380,17'd9372,17'd20381,17'd14832,17'd19982,17'd20382,17'd20383,17'd20113,17'd19846,17'd18851,17'd19086,17'd19086,17'd15093,17'd15475,17'd15723,17'd16118,17'd17171,17'd17171,17'd16370,17'd16246,17'd16118,17'd15604,17'd15475,17'd16119,17'd16247,17'd18134,17'd20384,17'd20385,17'd20386,17'd19224,17'd20387,17'd11859,17'd12477,17'd20388,17'd18977,17'd19353,17'd20389,17'd20390,17'd4700,17'd20391,17'd20392,17'd20393,17'd20394,17'd20395,17'd20396,17'd20397,17'd20398,17'd20399,17'd20400,17'd433,17'd186,17'd409,17'd20401,17'd1819,17'd6249,17'd4064,17'd7031,17'd7031,17'd6576,17'd8169,17'd9252,17'd8796,17'd8797,17'd9946,17'd9254,17'd11051,17'd18146,17'd18146,17'd18146,17'd18146,17'd20402,17'd18146,17'd9948,17'd9948,17'd19866,17'd19866,17'd12918,17'd12776,17'd9948,17'd9948,17'd20403,17'd19867,17'd10079,17'd9952,17'd9951,17'd12179,17'd4412,17'd3726,17'd3726,17'd3881,17'd8025,17'd5640,17'd20268,17'd20269,17'd6412,17'd5951,17'd4574,17'd20270,17'd2420,17'd181,17'd252,17'd252
},
'{
17'd1831,17'd1831,17'd4247,17'd466,17'd12,17'd3,17'd806,17'd806,17'd20404,17'd20404,17'd20,17'd4,17'd6,17'd3753,17'd8040,17'd8339,17'd8339,17'd8339,17'd8040,17'd8040,17'd8040,17'd8040,17'd8040,17'd5793,17'd3753,17'd3753,17'd3753,17'd6,17'd5,17'd24,17'd5,17'd5,17'd6,17'd3753,17'd6,17'd6,17'd1690,17'd1690,17'd1691,17'd1691,17'd7385,17'd7060,17'd4431,17'd3255,17'd13066,17'd20405,17'd825,17'd65,17'd20406,17'd20407,17'd20408,17'd20409,17'd20410,17'd20411,17'd20134,17'd20412,17'd20413,17'd20414,17'd20415,17'd20416,17'd14607,17'd20417,17'd20418,17'd20419,17'd19002,17'd18882,17'd16275,17'd20420,17'd13199,17'd20144,17'd20421,17'd17091,17'd16876,17'd19752,17'd18531,17'd15383,17'd15137,17'd12530,17'd12361,17'd14622,17'd14764,17'd14890,17'd13599,17'd13092,17'd13597,17'd12357,17'd13092,17'd12527,17'd13094,17'd12361,17'd12681,17'd20422,17'd20422,17'd20423,17'd12681,17'd12532,17'd20424,17'd18884,17'd17689,17'd17205,17'd18656,17'd20425,17'd17207,17'd17318,17'd20426,17'd20427,17'd20294,17'd20428,17'd20429,17'd20430,17'd20431,17'd20432,17'd20433,17'd19898,17'd20434,17'd12067,17'd20435,17'd20436,17'd9581,17'd9582,17'd14109,17'd14109,17'd14109,17'd14109,17'd9309,17'd9583,17'd9444,17'd18423,17'd20437,17'd20438,17'd20439,17'd20439,17'd19762,17'd19269,17'd19269,17'd18310,17'd20440,17'd20441,17'd15790,17'd20442,17'd19769,17'd20443,17'd10446,17'd19029,17'd18318,17'd12089,17'd20444,17'd20445,17'd20446,17'd15671,17'd12986,17'd12086,17'd15674,17'd13506,17'd18800,17'd11797,17'd20447,17'd20448,17'd13763,17'd11959,17'd11274,17'd10167,17'd18441,17'd17719,17'd11528,17'd11527,17'd14134,17'd19282,17'd14931,17'd10989,17'd11963,17'd11961,17'd12718,17'd12577,17'd12109,17'd13517,17'd12256,17'd12418,17'd12417,17'd12107,17'd20449,17'd20450,17'd18681,17'd16326,17'd11963,17'd13362,17'd13135,17'd13883,17'd18917,17'd12582,17'd19158,17'd13516,17'd20451,17'd10989,17'd13135,17'd16321,17'd12416,17'd14672,17'd16799,17'd16799,17'd16799,17'd12997,17'd12860,17'd12254,17'd20452,17'd18564,17'd13884,17'd12577,17'd11521,17'd12585,17'd8874,17'd20453,17'd20454,17'd7946,17'd13006,17'd10341,17'd20455,17'd20456,17'd15438,17'd19648,17'd17132,17'd17132,17'd20457,17'd20181,17'd20458,17'd20459,17'd20460,17'd20461,17'd20462,17'd20463,17'd20464,17'd20465,17'd5593,17'd131,17'd132,17'd133,17'd133,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd1481,17'd1481,17'd130,17'd130,17'd132,17'd132,17'd131,17'd131,17'd134,17'd132,17'd130,17'd130,17'd1481,17'd1481,17'd134,17'd131,17'd132,17'd134,17'd130,17'd130,17'd130,17'd136,17'd136,17'd136,17'd136,17'd138,17'd128,17'd134,17'd134,17'd20466,17'd1197,17'd132,17'd3168,17'd20467,17'd19045,17'd20468,17'd20469,17'd20470,17'd20471,17'd20472,17'd20473,17'd20474,17'd20475,17'd20476,17'd20477,17'd20478,17'd20479,17'd20480,17'd20481,17'd20203,17'd20482,17'd20345,17'd20483,17'd20484,17'd20485,17'd20486,17'd19561,17'd19316,17'd20487,17'd20488,17'd20489,17'd20490,17'd18233,17'd20491,17'd20492,17'd20493,17'd20494,17'd20495,17'd18610,17'd19706,17'd20496,17'd20372,17'd20497,17'd20498,17'd20499,17'd20500,17'd20221,17'd20501,17'd20502,17'd20503,17'd20504,17'd20505,17'd20359,17'd20506,17'd20507,17'd20226,17'd20227,17'd20508,17'd20509,17'd20510,17'd20511,17'd20512,17'd20513,17'd20513,17'd20514,17'd20515,17'd20516,17'd20517,17'd20518,17'd20519,17'd20370,17'd20520,17'd20521,17'd19837,17'd20522,17'd19822,17'd20523,17'd20524,17'd20525,17'd20526,17'd20104,17'd20104,17'd20527,17'd19452,17'd20528,17'd20529,17'd20530,17'd20376,17'd19342,17'd19080,17'd20531,17'd11295,17'd20532,17'd20533,17'd20534,17'd20535,17'd20536,17'd20537,17'd20538,17'd20539,17'd20540,17'd20541,17'd20541,17'd16247,17'd17779,17'd20542,17'd16246,17'd17171,17'd17171,17'd16370,17'd16613,17'd15986,17'd15474,17'd15724,17'd16371,17'd19087,17'd20543,17'd20544,17'd20545,17'd20546,17'd20547,17'd20548,17'd20549,17'd20550,17'd20551,17'd20552,17'd20553,17'd20554,17'd11438,17'd20555,17'd20392,17'd20556,17'd20557,17'd20558,17'd20559,17'd20126,17'd20560,17'd20561,17'd20562,17'd20563,17'd1683,17'd457,17'd20564,17'd20565,17'd5039,17'd3082,17'd4063,17'd4405,17'd4718,17'd11189,17'd9109,17'd9109,17'd8796,17'd8955,17'd9254,17'd11723,17'd12020,17'd10078,17'd19866,17'd18146,17'd12918,17'd12776,17'd10078,17'd20566,17'd9794,17'd9794,17'd11329,17'd11724,17'd11874,17'd10249,17'd20403,17'd20005,17'd20567,17'd11053,17'd9540,17'd8323,17'd7861,17'd3406,17'd3883,17'd3724,17'd7350,17'd6876,17'd20568,17'd4416,17'd4725,17'd4877,17'd3093,17'd2584,17'd2420,17'd1683,17'd252,17'd20569
},
'{
17'd1688,17'd1688,17'd1127,17'd2,17'd12,17'd3,17'd806,17'd806,17'd20404,17'd1128,17'd21,17'd4,17'd6,17'd3753,17'd8040,17'd8339,17'd8339,17'd8339,17'd8040,17'd8040,17'd8040,17'd8040,17'd8040,17'd5793,17'd3753,17'd3753,17'd6,17'd5,17'd5,17'd24,17'd4,17'd5,17'd3753,17'd3753,17'd6,17'd6,17'd1690,17'd1690,17'd1691,17'd1691,17'd20570,17'd7060,17'd4091,17'd3104,17'd1840,17'd20571,17'd58,17'd15366,17'd674,17'd20572,17'd18870,17'd20573,17'd20574,17'd20575,17'd20278,17'd20576,17'd20577,17'd18876,17'd20578,17'd15250,17'd20579,17'd20140,17'd20580,17'd19748,17'd16400,17'd16275,17'd20581,17'd20581,17'd16021,17'd20582,17'd20288,17'd20583,17'd20584,17'd20022,17'd18532,17'd14890,17'd12360,17'd12530,17'd12361,17'd12361,17'd14621,17'd14890,17'd13209,17'd13092,17'd13597,17'd14469,17'd12527,17'd11626,17'd12956,17'd11913,17'd11362,17'd19753,17'd20423,17'd12681,17'd16658,17'd16765,17'd20424,17'd17317,17'd16766,17'd17205,17'd17572,17'd20425,17'd20585,17'd15766,17'd7083,17'd20586,17'd20587,17'd20428,17'd20429,17'd20588,17'd20589,17'd20590,17'd20591,17'd13475,17'd20032,17'd20435,17'd9845,17'd9706,17'd9581,17'd9164,17'd9164,17'd9164,17'd14109,17'd14109,17'd9309,17'd9583,17'd9444,17'd13483,17'd20592,17'd20593,17'd20594,17'd20594,17'd20595,17'd20596,17'd19269,17'd18546,17'd15660,17'd15542,17'd20597,17'd11486,17'd20598,17'd20599,17'd20600,17'd15667,17'd20601,17'd12406,17'd20445,17'd20445,17'd20602,17'd13247,17'd15674,17'd12235,17'd20603,17'd12094,17'd11946,17'd20604,17'd20605,17'd20606,17'd11960,17'd17478,17'd11400,17'd16912,17'd20607,17'd11276,17'd11527,17'd11527,17'd10476,17'd10854,17'd11965,17'd11964,17'd11806,17'd13761,17'd12109,17'd12109,17'd12417,17'd12417,17'd13512,17'd12418,17'd14807,17'd19408,17'd20608,17'd20609,17'd18681,17'd16326,17'd11963,17'd13362,17'd11958,17'd11958,17'd18917,17'd19158,17'd11396,17'd11808,17'd11129,17'd12262,17'd11958,17'd14807,17'd12416,17'd15687,17'd14672,17'd16799,17'd13512,17'd12859,17'd16685,17'd18564,17'd12254,17'd16685,17'd12578,17'd11806,17'd20610,17'd9742,17'd15297,17'd11137,17'd20611,17'd20612,17'd15440,17'd15439,17'd20455,17'd20613,17'd14266,17'd20614,17'd20615,17'd7627,17'd20616,17'd20617,17'd16571,17'd17022,17'd20618,17'd20619,17'd20620,17'd20621,17'd20622,17'd5593,17'd5593,17'd131,17'd133,17'd133,17'd133,17'd133,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd131,17'd131,17'd11541,17'd131,17'd131,17'd131,17'd11541,17'd11541,17'd11541,17'd20466,17'd20623,17'd20624,17'd20625,17'd20626,17'd20627,17'd20628,17'd20629,17'd20630,17'd20631,17'd20632,17'd20633,17'd19295,17'd20634,17'd20635,17'd20636,17'd20637,17'd20638,17'd20639,17'd20640,17'd20641,17'd20642,17'd20642,17'd20643,17'd20644,17'd20645,17'd19947,17'd19948,17'd19804,17'd19558,17'd20483,17'd20346,17'd18594,17'd20646,17'd17875,17'd20647,17'd20648,17'd18601,17'd20649,17'd20650,17'd20651,17'd20493,17'd20652,17'd20653,17'd20654,17'd18608,17'd20655,17'd20656,17'd20657,17'd20658,17'd20659,17'd20660,17'd20661,17'd20662,17'd20663,17'd20664,17'd20665,17'd20666,17'd20667,17'd20360,17'd20226,17'd20228,17'd20668,17'd20669,17'd20670,17'd20671,17'd20672,17'd20672,17'd20673,17'd20673,17'd20674,17'd20675,17'd20676,17'd20677,17'd20678,17'd20679,17'd20680,17'd20101,17'd20681,17'd20682,17'd20683,17'd19698,17'd20236,17'd20237,17'd20684,17'd20685,17'd20372,17'd20104,17'd20527,17'd20373,17'd20374,17'd20686,17'd20687,17'd19977,17'd20688,17'd18737,17'd14294,17'd20689,17'd20245,17'd20690,17'd20691,17'd20692,17'd20693,17'd20537,17'd20538,17'd20539,17'd20694,17'd20540,17'd20695,17'd20695,17'd17065,17'd17903,17'd15852,17'd16370,17'd17171,17'd17171,17'd20696,17'd16613,17'd16611,17'd17282,17'd16371,17'd18741,17'd19087,17'd20697,17'd13926,17'd20253,17'd20698,17'd20699,17'd20700,17'd20701,17'd20702,17'd18977,17'd20553,17'd13172,17'd19230,17'd19233,17'd20703,17'd20704,17'd20705,17'd20706,17'd20707,17'd20708,17'd20709,17'd20710,17'd20711,17'd20563,17'd213,17'd20712,17'd8485,17'd20713,17'd2755,17'd2756,17'd4563,17'd19104,17'd4718,17'd11189,17'd10248,17'd10248,17'd8796,17'd9534,17'd9793,17'd9110,17'd11329,17'd10078,17'd20714,17'd19866,17'd12918,17'd12776,17'd10078,17'd20566,17'd20715,17'd20716,17'd11329,17'd11724,17'd11874,17'd10249,17'd20403,17'd20005,17'd20567,17'd20567,17'd9540,17'd8323,17'd7861,17'd4721,17'd3883,17'd4411,17'd20717,17'd6876,17'd20718,17'd20719,17'd5953,17'd4877,17'd3242,17'd2416,17'd639,17'd1826,17'd252,17'd20720
},
'{
17'd1688,17'd1127,17'd2,17'd0,17'd3,17'd3,17'd806,17'd2423,17'd1128,17'd1128,17'd21,17'd4,17'd6,17'd5793,17'd8338,17'd8339,17'd8340,17'd8340,17'd8040,17'd8040,17'd8040,17'd8040,17'd5205,17'd3753,17'd3753,17'd3753,17'd6,17'd5,17'd24,17'd24,17'd5,17'd5,17'd3753,17'd3753,17'd6,17'd6,17'd1690,17'd1691,17'd1691,17'd1832,17'd20570,17'd4430,17'd5208,17'd2944,17'd1702,17'd991,17'd303,17'd19500,17'd20721,17'd1564,17'd20722,17'd20723,17'd20724,17'd20725,17'd20726,17'd20727,17'd19249,17'd20728,17'd20729,17'd20730,17'd20731,17'd20140,17'd20580,17'd13080,17'd13081,17'd16275,17'd20581,17'd20581,17'd13589,17'd20145,17'd17091,17'd20732,17'd20733,17'd20734,17'd18532,17'd18411,17'd15137,17'd12530,17'd12361,17'd12361,17'd14621,17'd12955,17'd13209,17'd13092,17'd13462,17'd13462,17'd13209,17'd13093,17'd12530,17'd11764,17'd11362,17'd11362,17'd12681,17'd12532,17'd12361,17'd16765,17'd12531,17'd19006,17'd17689,17'd18174,17'd17572,17'd17319,17'd16164,17'd20735,17'd20736,17'd18535,17'd20587,17'd20428,17'd20737,17'd20738,17'd20738,17'd13849,17'd13605,17'd13097,17'd12067,17'd20435,17'd9845,17'd9706,17'd20739,17'd20740,17'd9582,17'd9582,17'd9582,17'd9707,17'd9848,17'd9849,17'd9992,17'd13483,17'd20741,17'd20742,17'd20743,17'd20743,17'd20744,17'd20745,17'd18427,17'd18426,17'd20746,17'd14494,17'd10821,17'd20747,17'd10137,17'd20748,17'd20749,17'd11109,17'd19914,17'd20750,17'd20751,17'd20306,17'd13359,17'd20752,17'd20753,17'd20603,17'd13506,17'd18800,17'd19915,17'd19916,17'd14376,17'd15294,17'd11395,17'd11131,17'd20754,17'd20755,17'd16796,17'd20756,17'd10477,17'd10991,17'd10739,17'd10990,17'd10989,17'd11807,17'd13363,17'd12110,17'd12995,17'd13517,17'd12417,17'd12859,17'd12418,17'd12417,17'd14807,17'd18198,17'd14258,17'd19921,17'd16326,17'd19158,17'd12996,17'd18917,17'd11958,17'd12106,17'd18917,17'd12422,17'd10989,17'd11808,17'd10989,17'd11963,17'd12420,17'd12579,17'd12416,17'd14672,17'd16799,17'd16799,17'd14523,17'd13643,17'd12415,17'd12415,17'd18564,17'd15434,17'd12419,17'd11395,17'd11135,17'd20757,17'd15179,17'd11137,17'd7946,17'd7788,17'd10180,17'd10861,17'd14682,17'd19646,17'd19648,17'd14142,17'd13772,17'd15062,17'd17019,17'd15061,17'd15063,17'd20758,17'd20759,17'd20760,17'd20761,17'd717,17'd133,17'd131,17'd131,17'd131,17'd1481,17'd20762,17'd20762,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd132,17'd134,17'd128,17'd128,17'd134,17'd11541,17'd11541,17'd16090,17'd16090,17'd1759,17'd134,17'd131,17'd131,17'd11683,17'd11821,17'd20763,17'd20764,17'd20765,17'd20766,17'd20767,17'd20768,17'd20769,17'd20770,17'd20771,17'd20772,17'd20773,17'd20774,17'd20775,17'd20776,17'd20777,17'd20778,17'd20779,17'd20780,17'd20781,17'd20782,17'd20783,17'd20784,17'd20785,17'd20199,17'd20786,17'd20787,17'd20788,17'd20789,17'd20790,17'd20791,17'd20792,17'd20793,17'd20794,17'd19558,17'd20483,17'd20795,17'd19951,17'd18594,17'd20647,17'd20796,17'd20797,17'd20798,17'd20799,17'd20800,17'd20801,17'd20802,17'd20803,17'd20804,17'd20805,17'd18957,17'd20806,17'd20807,17'd20808,17'd20809,17'd20810,17'd20811,17'd20812,17'd20813,17'd20814,17'd20815,17'd20667,17'd20506,17'd20360,17'd20360,17'd20816,17'd20817,17'd20818,17'd20819,17'd20670,17'd20672,17'd20820,17'd20821,17'd20822,17'd20823,17'd20824,17'd20825,17'd20826,17'd20827,17'd20828,17'd20829,17'd20830,17'd20831,17'd20100,17'd20832,17'd19695,17'd19696,17'd20355,17'd20833,17'd20834,17'd20525,17'd20372,17'd20656,17'd20685,17'd20835,17'd20836,17'd20837,17'd20838,17'd20839,17'd20840,17'd18368,17'd15718,17'd20841,17'd20842,17'd13911,17'd20691,17'd20843,17'd20844,17'd20536,17'd20538,17'd20845,17'd20846,17'd20694,17'd20695,17'd20695,17'd16371,17'd17065,17'd15723,17'd16118,17'd16370,17'd17171,17'd16370,17'd16246,17'd16842,17'd17283,17'd17654,17'd20847,17'd19087,17'd20848,17'd20849,17'd19987,17'd20850,17'd20851,17'd20852,17'd11861,17'd20853,17'd20120,17'd20854,17'd20855,17'd19230,17'd20856,17'd7678,17'd20857,17'd20858,17'd20859,17'd20860,17'd20861,17'd20397,17'd20862,17'd20863,17'd20563,17'd251,17'd966,17'd20002,17'd20864,17'd6578,17'd2756,17'd6249,17'd3718,17'd4719,17'd11189,17'd10248,17'd7687,17'd8954,17'd8797,17'd9536,17'd9110,17'd11329,17'd11874,17'd9948,17'd9948,17'd12918,17'd12776,17'd10078,17'd9796,17'd9406,17'd12919,17'd11329,17'd10078,17'd11874,17'd11874,17'd11192,17'd20005,17'd20567,17'd11053,17'd8801,17'd8323,17'd7861,17'd4721,17'd3883,17'd3724,17'd7350,17'd6876,17'd7040,17'd5953,17'd5953,17'd20865,17'd20866,17'd20867,17'd1683,17'd17422,17'd20868,17'd20868
},
'{
17'd1688,17'd1127,17'd2,17'd0,17'd3,17'd3,17'd806,17'd2423,17'd1128,17'd11,17'd25,17'd4,17'd6,17'd5205,17'd8340,17'd8339,17'd8340,17'd8340,17'd8040,17'd8040,17'd8040,17'd8040,17'd3753,17'd3753,17'd3753,17'd3753,17'd5,17'd5,17'd24,17'd24,17'd5,17'd5,17'd5205,17'd3753,17'd6,17'd6,17'd1690,17'd1691,17'd1832,17'd285,17'd7060,17'd4431,17'd3434,17'd2602,17'd1282,17'd825,17'd20869,17'd20870,17'd20721,17'd18518,17'd20871,17'd20872,17'd1851,17'd20873,17'd20874,17'd20875,17'd16268,17'd5069,17'd20876,17'd20877,17'd20731,17'd20878,17'd20879,17'd20880,17'd13081,17'd16275,17'd20581,17'd16509,17'd13589,17'd20288,17'd20881,17'd20882,17'd20883,17'd20884,17'd18173,17'd14764,17'd13840,17'd12530,17'd12530,17'd12218,17'd12955,17'd13093,17'd13092,17'd13092,17'd13462,17'd13209,17'd12528,17'd12955,17'd13840,17'd11764,17'd11362,17'd11629,17'd12532,17'd12531,17'd12362,17'd20885,17'd20886,17'd17204,17'd17205,17'd17206,17'd16289,17'd16289,17'd19384,17'd20887,17'd20586,17'd18535,17'd20888,17'd20428,17'd20737,17'd20737,17'd20889,17'd20031,17'd20434,17'd12067,17'd10120,17'd9845,17'd9706,17'd9706,17'd20739,17'd20740,17'd9582,17'd9582,17'd9582,17'd9582,17'd9848,17'd9849,17'd9992,17'd20890,17'd20891,17'd20892,17'd20594,17'd20744,17'd20744,17'd20745,17'd18546,17'd17459,17'd20893,17'd13107,17'd20894,17'd20895,17'd20896,17'd18187,17'd14119,17'd13627,17'd20897,17'd20898,17'd20751,17'd20899,17'd20900,17'd20901,17'd20902,17'd20903,17'd20305,17'd20904,17'd20905,17'd20906,17'd20907,17'd20908,17'd10603,17'd17124,17'd20909,17'd16912,17'd10479,17'd10478,17'd14518,17'd11132,17'd10854,17'd11274,17'd11964,17'd11806,17'd12110,17'd12414,17'd12417,17'd12417,17'd12418,17'd12859,17'd12418,17'd14807,17'd18198,17'd18917,17'd18681,17'd18444,17'd16326,17'd15185,17'd18917,17'd17722,17'd12106,17'd12106,17'd18917,17'd12422,17'd11965,17'd20910,17'd19157,17'd12858,17'd12580,17'd12253,17'd12415,17'd12860,17'd12997,17'd14523,17'd14523,17'd13643,17'd12416,17'd12416,17'd12579,17'd13882,17'd12861,17'd13886,17'd9620,17'd8883,17'd20176,17'd12865,17'd12120,17'd10180,17'd15439,17'd20455,17'd18921,17'd12429,17'd14533,17'd8429,17'd8739,17'd17485,17'd20911,17'd16570,17'd20912,17'd20913,17'd9355,17'd20914,17'd20915,17'd717,17'd133,17'd134,17'd131,17'd132,17'd1481,17'd20762,17'd20762,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd131,17'd132,17'd130,17'd130,17'd130,17'd132,17'd131,17'd131,17'd20622,17'd20622,17'd11541,17'd11541,17'd11683,17'd20916,17'd20917,17'd20769,17'd20918,17'd20919,17'd20920,17'd20921,17'd20922,17'd20923,17'd20924,17'd20925,17'd20926,17'd20926,17'd20927,17'd20928,17'd20929,17'd20930,17'd20931,17'd20932,17'd20933,17'd20934,17'd20935,17'd20936,17'd20937,17'd20938,17'd20939,17'd20940,17'd20941,17'd20942,17'd20943,17'd20944,17'd20945,17'd20946,17'd20947,17'd20948,17'd20949,17'd20950,17'd20483,17'd20951,17'd20795,17'd20952,17'd20208,17'd20953,17'd20954,17'd20955,17'd20956,17'd20957,17'd20958,17'd20959,17'd20960,17'd20961,17'd20962,17'd20963,17'd20964,17'd20965,17'd20355,17'd19695,17'd19961,17'd20966,17'd20967,17'd20967,17'd20664,17'd20815,17'd20667,17'd20360,17'd20360,17'd20968,17'd20363,17'd20969,17'd20669,17'd20970,17'd20971,17'd20972,17'd20973,17'd20974,17'd20975,17'd20976,17'd20977,17'd20977,17'd20978,17'd20979,17'd20980,17'd20981,17'd20829,17'd20982,17'd20983,17'd20984,17'd20985,17'd19969,17'd20089,17'd20986,17'd20987,17'd20834,17'd20525,17'd20684,17'd20988,17'd20685,17'd20989,17'd20837,17'd20838,17'd20990,17'd20991,17'd15717,17'd14416,17'd20992,17'd20993,17'd20994,17'd20995,17'd20996,17'd20997,17'd20693,17'd20998,17'd20999,17'd21000,17'd20846,17'd21001,17'd20695,17'd16371,17'd16371,17'd15475,17'd15604,17'd16246,17'd17171,17'd16370,17'd16246,17'd21002,17'd16842,17'd15603,17'd18133,17'd18741,17'd19479,17'd18852,17'd19715,17'd21003,17'd21004,17'd21005,17'd21006,17'd21007,17'd20389,17'd21008,17'd20855,17'd21009,17'd20258,17'd6075,17'd21010,17'd21011,17'd21012,17'd21013,17'd21014,17'd21015,17'd21016,17'd1086,17'd20563,17'd250,17'd460,17'd21017,17'd21018,17'd6252,17'd2757,17'd3404,17'd13291,17'd5033,17'd11189,17'd10248,17'd7687,17'd8954,17'd8797,17'd9536,17'd9110,17'd11329,17'd11874,17'd11192,17'd9948,17'd12776,17'd12640,17'd9947,17'd9796,17'd9406,17'd21019,17'd9947,17'd10078,17'd11874,17'd10249,17'd20403,17'd20005,17'd20567,17'd20567,17'd9540,17'd8648,17'd7861,17'd4721,17'd3883,17'd4411,17'd21020,17'd6876,17'd6882,17'd5951,17'd4725,17'd3093,17'd21021,17'd20867,17'd1683,17'd1548,17'd15626,17'd15355
},
'{
17'd4247,17'd1127,17'd2,17'd0,17'd3,17'd12,17'd2423,17'd2423,17'd11,17'd10,17'd9,17'd8,17'd7,17'd8040,17'd8339,17'd8339,17'd8340,17'd8340,17'd8040,17'd8040,17'd8040,17'd8040,17'd3753,17'd3753,17'd3594,17'd3594,17'd5,17'd24,17'd24,17'd24,17'd5,17'd3594,17'd8040,17'd5793,17'd3753,17'd6,17'd1690,17'd1691,17'd7385,17'd7060,17'd4430,17'd3755,17'd3104,17'd1973,17'd1134,17'd57,17'd21022,17'd21023,17'd19501,17'd21024,17'd21025,17'd21026,17'd1852,17'd21027,17'd21028,17'd20135,17'd21029,17'd21030,17'd14994,17'd21031,17'd21032,17'd21033,17'd21034,17'd19002,17'd13198,17'd20581,17'd16155,17'd13448,17'd18165,17'd14089,17'd19751,17'd20021,17'd21035,17'd21036,17'd20147,17'd14764,17'd13840,17'd12530,17'd14621,17'd14621,17'd13093,17'd13093,17'd13092,17'd13092,17'd13092,17'd13209,17'd12528,17'd14890,17'd13840,17'd13969,17'd12532,17'd12531,17'd12531,17'd20424,17'd12362,17'd12361,17'd12532,17'd17941,17'd17205,17'd17206,17'd16289,17'd16164,17'd21037,17'd21038,17'd20586,17'd18535,17'd21039,17'd21040,17'd20889,17'd13848,17'd21041,17'd13474,17'd21042,17'd11916,17'd10120,17'd20435,17'd20436,17'd9706,17'd20739,17'd20740,17'd9846,17'd9846,17'd9990,17'd10288,17'd10122,17'd10568,17'd13731,17'd21043,17'd21044,17'd21044,17'd20594,17'd19629,17'd19396,17'd18311,17'd18426,17'd16297,17'd21045,17'd10950,17'd21046,17'd19771,17'd21047,17'd18909,17'd12395,17'd19639,17'd21048,17'd21049,17'd20306,17'd18189,17'd13505,17'd21050,17'd21051,17'd21052,17'd21053,17'd21054,17'd19778,17'd21055,17'd15047,17'd10605,17'd9618,17'd9341,17'd21056,17'd9883,17'd10478,17'd10478,17'd11132,17'd11399,17'd11274,17'd11964,17'd13135,17'd11960,17'd12110,17'd12109,17'd12418,17'd12415,17'd12415,17'd12416,17'd12108,17'd17348,17'd15053,17'd16204,17'd11964,17'd13516,17'd19158,17'd16325,17'd17722,17'd20314,17'd20314,17'd17722,17'd12582,17'd12115,17'd11965,17'd10989,17'd12114,17'd12420,17'd12109,17'd12253,17'd15434,17'd12859,17'd12859,17'd12418,17'd14525,17'd21057,17'd14003,17'd12253,17'd15184,17'd13764,17'd14810,17'd17839,17'd19033,17'd8724,17'd8409,17'd14384,17'd15948,17'd21058,17'd16078,17'd18921,17'd21059,17'd14678,17'd10031,17'd18810,17'd7629,17'd21060,17'd21061,17'd16807,17'd21062,17'd21063,17'd21064,17'd21065,17'd21066,17'd541,17'd130,17'd129,17'd132,17'd132,17'd1481,17'd20762,17'd20762,17'd20762,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd136,17'd130,17'd132,17'd131,17'd131,17'd131,17'd130,17'd130,17'd136,17'd130,17'd130,17'd132,17'd11541,17'd131,17'd133,17'd13777,17'd21067,17'd21068,17'd21069,17'd20773,17'd21070,17'd21071,17'd21072,17'd21073,17'd21074,17'd21075,17'd21076,17'd21076,17'd21077,17'd21078,17'd21078,17'd21079,17'd21080,17'd21081,17'd21082,17'd21083,17'd21084,17'd21085,17'd21086,17'd21087,17'd21088,17'd21089,17'd21090,17'd21091,17'd21092,17'd21093,17'd21094,17'd21095,17'd21096,17'd21097,17'd21098,17'd20946,17'd21099,17'd21100,17'd21101,17'd20483,17'd20483,17'd21102,17'd21103,17'd21104,17'd18109,17'd21105,17'd17875,17'd20211,17'd21106,17'd21107,17'd21108,17'd21109,17'd21110,17'd20960,17'd21111,17'd21112,17'd19074,17'd21113,17'd19699,17'd19691,17'd20505,17'd20966,17'd20967,17'd20663,17'd20505,17'd21114,17'd21115,17'd20360,17'd20816,17'd20817,17'd20668,17'd20669,17'd20514,17'd21116,17'd20825,17'd21117,17'd21118,17'd21119,17'd21120,17'd21121,17'd21122,17'd21123,17'd21124,17'd21125,17'd21125,17'd20979,17'd20827,17'd21126,17'd21127,17'd21128,17'd21129,17'd20985,17'd19835,17'd21130,17'd20833,17'd21131,17'd21132,17'd21133,17'd21134,17'd21135,17'd21136,17'd21137,17'd21138,17'd20990,17'd21139,17'd21140,17'd21141,17'd21142,17'd21143,17'd21144,17'd21145,17'd21146,17'd21147,17'd20844,17'd20537,17'd20538,17'd21000,17'd20846,17'd21001,17'd20695,17'd16371,17'd16371,17'd16119,17'd15723,17'd16118,17'd16246,17'd16246,17'd16246,17'd21002,17'd16843,17'd18132,17'd17654,17'd16371,17'd18620,17'd21148,17'd19986,17'd21149,17'd21150,17'd21151,17'd11582,17'd11861,17'd21007,17'd20389,17'd19486,17'd13172,17'd21152,17'd21153,17'd21154,17'd21155,17'd20557,17'd21156,17'd21157,17'd21158,17'd21159,17'd21160,17'd786,17'd249,17'd1095,17'd21161,17'd8485,17'd21162,17'd2755,17'd3404,17'd13291,17'd4063,17'd8318,17'd10248,17'd8490,17'd9252,17'd8797,17'd9536,17'd11594,17'd11873,17'd11874,17'd11192,17'd9948,17'd12776,17'd12640,17'd9794,17'd21163,17'd21019,17'd8646,17'd9111,17'd9111,17'd11874,17'd11874,17'd9256,17'd9796,17'd21163,17'd11053,17'd9407,17'd8648,17'd4567,17'd3233,17'd3726,17'd3724,17'd8025,17'd6876,17'd21164,17'd5044,17'd5642,17'd3242,17'd4417,17'd2110,17'd182,17'd17422,17'd21165,17'd21165
},
'{
17'd4247,17'd1127,17'd2,17'd0,17'd12,17'd12,17'd2423,17'd2423,17'd11,17'd25,17'd4,17'd6,17'd5205,17'd8190,17'd8340,17'd8339,17'd8340,17'd8340,17'd8040,17'd8040,17'd8040,17'd8040,17'd3753,17'd3753,17'd3594,17'd3594,17'd5,17'd24,17'd24,17'd24,17'd5,17'd6,17'd3753,17'd3753,17'd6,17'd5,17'd1691,17'd285,17'd7061,17'd6744,17'd4431,17'd3754,17'd2601,17'd2121,17'd990,17'd58,17'd21166,17'd21167,17'd21168,17'd20871,17'd20872,17'd21169,17'd21170,17'd21171,17'd20874,17'd21172,17'd3768,17'd21173,17'd21174,17'd21175,17'd21176,17'd21177,17'd21178,17'd19002,17'd21179,17'd20581,17'd16155,17'd13704,17'd21180,17'd21181,17'd21182,17'd21183,17'd21036,17'd18173,17'd14622,17'd14622,17'd13969,17'd12530,17'd14621,17'd12955,17'd13093,17'd12813,17'd13092,17'd13092,17'd13092,17'd21184,17'd14890,17'd15137,17'd13840,17'd13840,17'd11764,17'd12531,17'd20424,17'd20424,17'd12361,17'd12531,17'd17204,17'd18774,17'd17206,17'd21185,17'd16289,17'd19384,17'd20887,17'd21186,17'd20736,17'd21187,17'd20294,17'd20295,17'd21188,17'd21041,17'd21189,17'd13604,17'd21190,17'd10119,17'd10120,17'd9845,17'd9706,17'd9706,17'd20739,17'd20739,17'd9846,17'd9846,17'd10288,17'd10288,17'd10122,17'd10568,17'd13731,17'd14779,17'd21191,17'd21192,17'd20439,17'd21193,17'd19764,17'd18310,17'd17703,17'd21194,17'd21195,17'd21196,17'd21197,17'd21198,17'd19636,17'd21199,17'd11937,17'd21200,17'd21048,17'd21201,17'd13359,17'd13506,17'd13505,17'd20903,17'd12406,17'd21202,17'd19915,17'd20447,17'd21203,17'd21204,17'd12720,17'd10479,17'd9344,17'd9191,17'd9885,17'd11527,17'd21205,17'd15176,17'd21206,17'd11808,17'd11964,17'd15185,17'd13761,17'd15184,17'd12414,17'd12579,17'd12416,17'd12860,17'd12415,17'd14003,17'd19407,17'd20314,17'd12582,17'd12262,17'd14262,17'd11964,17'd19158,17'd16325,17'd18559,17'd20314,17'd18559,17'd18557,17'd12422,17'd12115,17'd10989,17'd13362,17'd13519,17'd12995,17'd12414,17'd12253,17'd15434,17'd15434,17'd12253,17'd12417,17'd21207,17'd21207,17'd12416,17'd15434,17'd19645,17'd12862,17'd10164,17'd9342,17'd8882,17'd8574,17'd21208,17'd21209,17'd21210,17'd21211,17'd21058,17'd19288,17'd14392,17'd20616,17'd15951,17'd21212,17'd16569,17'd21213,17'd21214,17'd21215,17'd21216,17'd21217,17'd21218,17'd10757,17'd21219,17'd1196,17'd128,17'd132,17'd132,17'd132,17'd130,17'd1481,17'd1481,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd136,17'd136,17'd130,17'd132,17'd132,17'd132,17'd130,17'd130,17'd720,17'd128,17'd130,17'd134,17'd131,17'd131,17'd19655,17'd21220,17'd21221,17'd21222,17'd21223,17'd21224,17'd21225,17'd21226,17'd21227,17'd21228,17'd21229,17'd21230,17'd21231,17'd21232,17'd21233,17'd21234,17'd21235,17'd21236,17'd21237,17'd21238,17'd21239,17'd21240,17'd21241,17'd21242,17'd21243,17'd21244,17'd21245,17'd21246,17'd21247,17'd21248,17'd21249,17'd21250,17'd21251,17'd21252,17'd21253,17'd21254,17'd21255,17'd21256,17'd21257,17'd21258,17'd21259,17'd19804,17'd21260,17'd21261,17'd21262,17'd21263,17'd18947,17'd20647,17'd17875,17'd21264,17'd21265,17'd21266,17'd21267,17'd21268,17'd21269,17'd21110,17'd21270,17'd21271,17'd19332,17'd21272,17'd19463,17'd19691,17'd20966,17'd21273,17'd21274,17'd20664,17'd20665,17'd21275,17'd20225,17'd21276,17'd20817,17'd20969,17'd20669,17'd20970,17'd21277,17'd20972,17'd21278,17'd20977,17'd20976,17'd21279,17'd21280,17'd21281,17'd21282,17'd21283,17'd21283,17'd21284,17'd21285,17'd21286,17'd21287,17'd21288,17'd21289,17'd21290,17'd21128,17'd21291,17'd20369,17'd20089,17'd21130,17'd21292,17'd21293,17'd21294,17'd21295,17'd21296,17'd21297,17'd21298,17'd21137,17'd21138,17'd21299,17'd21300,17'd21301,17'd21302,17'd21143,17'd10360,17'd21303,17'd21304,17'd21305,17'd21306,17'd20693,17'd20998,17'd21307,17'd20846,17'd21001,17'd21001,17'd16247,17'd16247,17'd16119,17'd15603,17'd15604,17'd16118,17'd16118,17'd16118,17'd21308,17'd17063,17'd15604,17'd17534,17'd17065,17'd16247,17'd21309,17'd21310,17'd21311,17'd21312,17'd21313,17'd21314,17'd11714,17'd21315,17'd21316,17'd19854,17'd20553,17'd12768,17'd21317,17'd7679,17'd21318,17'd21319,17'd21320,17'd21321,17'd21322,17'd2091,17'd21323,17'd21324,17'd21325,17'd634,17'd772,17'd20002,17'd21326,17'd6578,17'd3404,17'd13291,17'd4063,17'd8318,17'd7687,17'd8490,17'd8794,17'd9109,17'd9406,17'd11594,17'd11873,17'd11874,17'd11192,17'd9948,17'd12640,17'd9948,17'd9794,17'd20567,17'd12321,17'd12321,17'd8956,17'd9111,17'd10249,17'd10249,17'd20716,17'd9796,17'd21163,17'd21163,17'd9665,17'd9540,17'd4413,17'd21327,17'd21328,17'd4411,17'd21020,17'd6876,17'd21164,17'd5187,17'd5642,17'd3242,17'd4417,17'd2771,17'd181,17'd17422,17'd179,17'd17075
},
'{
17'd1127,17'd1127,17'd2,17'd0,17'd12,17'd12,17'd2423,17'd2423,17'd20,17'd25,17'd8,17'd6,17'd5205,17'd8190,17'd10795,17'd8340,17'd8340,17'd8340,17'd8040,17'd8040,17'd5205,17'd5205,17'd3753,17'd3594,17'd5,17'd5,17'd24,17'd24,17'd24,17'd24,17'd5,17'd6,17'd3753,17'd3753,17'd7554,17'd7383,17'd1691,17'd285,17'd7060,17'd6744,17'd3755,17'd3431,17'd2263,17'd1282,17'd825,17'd21329,17'd15248,17'd19610,17'd21330,17'd20871,17'd21331,17'd21332,17'd21333,17'd21334,17'd21335,17'd2628,17'd21336,17'd21337,17'd21338,17'd21339,17'd21340,17'd21341,17'd19619,17'd16400,17'd20581,17'd20287,17'd13448,17'd15635,17'd21342,17'd21343,17'd21344,17'd20884,17'd20147,17'd14622,17'd14622,17'd12361,17'd12361,17'd12530,17'd12955,17'd12679,17'd13209,17'd13092,17'd13092,17'd13092,17'd13209,17'd21184,17'd15137,17'd16286,17'd13840,17'd13840,17'd11913,17'd11913,17'd20424,17'd12531,17'd12531,17'd12532,17'd17941,17'd18774,17'd17206,17'd21185,17'd16164,17'd18658,17'd21345,17'd6768,17'd20586,17'd18659,17'd20294,17'd21039,17'd21346,17'd21346,17'd13329,17'd9003,17'd21190,17'd10119,17'd10120,17'd9845,17'd9706,17'd9580,17'd9580,17'd9580,17'd9988,17'd9989,17'd10948,17'd11092,17'd11483,17'd21347,17'd13854,17'd14779,17'd13730,17'd21348,17'd21193,17'd21349,17'd18899,17'd18789,17'd21350,17'd21351,17'd21352,17'd21353,17'd20599,17'd21354,17'd13872,17'd11648,17'd21355,17'd21356,17'd21357,17'd21358,17'd20902,17'd15676,17'd20900,17'd19914,17'd12407,17'd21359,17'd14924,17'd12573,17'd21360,17'd11520,17'd11133,17'd10992,17'd10335,17'd10335,17'd16070,17'd10478,17'd10477,17'd11132,17'd10854,17'd11274,17'd19158,17'd13883,17'd12110,17'd12578,17'd12859,17'd14003,17'd12416,17'd12415,17'd19534,17'd13515,17'd19407,17'd18197,17'd17604,17'd13516,17'd14262,17'd13762,17'd16442,17'd21361,17'd21362,17'd21363,17'd18197,17'd18806,17'd12115,17'd18560,17'd15810,17'd11957,17'd21364,17'd13518,17'd12575,17'd12414,17'd18450,17'd12414,17'd12253,17'd12417,17'd21207,17'd21207,17'd12416,17'd12578,17'd13764,17'd10477,17'd10743,17'd16910,17'd12118,17'd9349,17'd8581,17'd8256,17'd15949,17'd21365,17'd15303,17'd21366,17'd8586,17'd14393,17'd21367,17'd21368,17'd21369,17'd21370,17'd21371,17'd21372,17'd21373,17'd21374,17'd10617,17'd7812,17'd717,17'd1197,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd136,17'd136,17'd136,17'd136,17'd130,17'd130,17'd130,17'd130,17'd130,17'd132,17'd21375,17'd21376,17'd21377,17'd21222,17'd21378,17'd21379,17'd21380,17'd21381,17'd21382,17'd21383,17'd21384,17'd21385,17'd21385,17'd21386,17'd21387,17'd21388,17'd21389,17'd21390,17'd21391,17'd21233,17'd21392,17'd21393,17'd21394,17'd21395,17'd21396,17'd21397,17'd21398,17'd21399,17'd21400,17'd21401,17'd21402,17'd21403,17'd21404,17'd21405,17'd21406,17'd21407,17'd21252,17'd21097,17'd21408,17'd21409,17'd21410,17'd21411,17'd21412,17'd19671,17'd21413,17'd21413,17'd21414,17'd21415,17'd19951,17'd20208,17'd17875,17'd21264,17'd21416,17'd21266,17'd21417,17'd21418,17'd21419,17'd21420,17'd20960,17'd21421,17'd21422,17'd21423,17'd19826,17'd20502,17'd20966,17'd21424,17'd21274,17'd21425,17'd20665,17'd20667,17'd21426,17'd21427,17'd20817,17'd20364,17'd20515,17'd21428,17'd20972,17'd21429,17'd20976,17'd21430,17'd21121,17'd21431,17'd21432,17'd21433,17'd21434,17'd21435,17'd21435,17'd21436,17'd21437,17'd21438,17'd21439,17'd21440,17'd21441,17'd21442,17'd21443,17'd20518,17'd21444,17'd21445,17'd20219,17'd20088,17'd21446,17'd21293,17'd21447,17'd21448,17'd21449,17'd21297,17'd21298,17'd21450,17'd21299,17'd21139,17'd21451,17'd21452,17'd12136,17'd10882,17'd8915,17'd14026,17'd20995,17'd21305,17'd20997,17'd20537,17'd21307,17'd20694,17'd21001,17'd21001,17'd16247,17'd16247,17'd16371,17'd17065,17'd15724,17'd17283,17'd17063,17'd16844,17'd16246,17'd16118,17'd15604,17'd15603,17'd15605,17'd16371,17'd21453,17'd19714,17'd19715,17'd21454,17'd21455,17'd21456,17'd11582,17'd21457,17'd21007,17'd19854,17'd20553,17'd21458,17'd19723,17'd21459,17'd21460,17'd21461,17'd21462,17'd21463,17'd21464,17'd21465,17'd21466,17'd21467,17'd21468,17'd963,17'd2588,17'd19493,17'd21469,17'd6578,17'd2759,17'd21470,17'd4563,17'd9116,17'd8490,17'd7688,17'd11189,17'd10248,17'd9406,17'd9255,17'd11873,17'd21471,17'd11330,17'd11192,17'd12640,17'd9948,17'd9794,17'd20567,17'd21472,17'd12023,17'd8956,17'd9111,17'd10249,17'd10249,17'd20716,17'd21163,17'd21163,17'd21163,17'd11053,17'd8647,17'd10390,17'd4568,17'd4566,17'd3724,17'd7350,17'd6876,17'd6877,17'd5187,17'd6411,17'd3417,17'd4417,17'd2771,17'd1822,17'd590,17'd17075,17'd17552
},
'{
17'd1127,17'd14,17'd0,17'd0,17'd12,17'd12,17'd2423,17'd806,17'd21,17'd4,17'd6,17'd6,17'd5205,17'd8190,17'd10795,17'd8340,17'd8340,17'd8340,17'd8040,17'd8040,17'd5205,17'd5205,17'd3753,17'd3594,17'd24,17'd24,17'd24,17'd24,17'd24,17'd24,17'd6,17'd7,17'd3753,17'd3753,17'd7383,17'd1690,17'd467,17'd286,17'd6744,17'd18037,17'd3255,17'd2942,17'd1972,17'd1134,17'd57,17'd61,17'd21473,17'd19610,17'd21474,17'd21475,17'd21476,17'd21332,17'd21477,17'd21478,17'd21479,17'd21480,17'd15249,17'd13310,17'd21481,17'd13077,17'd21482,17'd20419,17'd19120,17'd12941,17'd20581,17'd13449,17'd18404,17'd13827,17'd21181,17'd21483,17'd21484,17'd21036,17'd14622,17'd14764,17'd12361,17'd16765,17'd12361,17'd12530,17'd12955,17'd12679,17'd13209,17'd13092,17'd13092,17'd13092,17'd13209,17'd12528,17'd15137,17'd16286,17'd12530,17'd13840,17'd11913,17'd11913,17'd12531,17'd12531,17'd12532,17'd19006,17'd17689,17'd16986,17'd21185,17'd21185,17'd19256,17'd18658,17'd21345,17'd6299,17'd21485,17'd18415,17'd20294,17'd21486,17'd21487,17'd21487,17'd21488,17'd7580,17'd21489,17'd10119,17'd9705,17'd9845,17'd9706,17'd9580,17'd9579,17'd9845,17'd9988,17'd10698,17'd10948,17'd11092,17'd11483,17'd21347,17'd13854,17'd14779,17'd14636,17'd21490,17'd21193,17'd21491,17'd21492,17'd21493,17'd15790,17'd14784,17'd21494,17'd21495,17'd18433,17'd18674,17'd21496,17'd11939,17'd21497,17'd20898,17'd21498,17'd13359,17'd20901,17'd19774,17'd20900,17'd12094,17'd21499,17'd21500,17'd21501,17'd21502,17'd16797,17'd10854,17'd21503,17'd15295,17'd10335,17'd17601,17'd17599,17'd10478,17'd11132,17'd11399,17'd14673,17'd11964,17'd18917,17'd15184,17'd12414,17'd15434,17'd12860,17'd12416,17'd12416,17'd12415,17'd21504,17'd19407,17'd19408,17'd12582,17'd19643,17'd13516,17'd13762,17'd15185,17'd21361,17'd21362,17'd21363,17'd21505,17'd18917,17'd17604,17'd12115,17'd18560,17'd12262,17'd12420,17'd21506,17'd14809,17'd12575,17'd12414,17'd18450,17'd18450,17'd16203,17'd14807,17'd14003,17'd13515,17'd12417,17'd13364,17'd12862,17'd16070,17'd8874,17'd21507,17'd8728,17'd18919,17'd8254,17'd15692,17'd21508,17'd13377,17'd19536,17'd14141,17'd21509,17'd21510,17'd16805,17'd21511,17'd21512,17'd21513,17'd21514,17'd21515,17'd21516,17'd21517,17'd17025,17'd21518,17'd17363,17'd134,17'd132,17'd135,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd136,17'd136,17'd136,17'd130,17'd132,17'd132,17'd131,17'd11541,17'd20627,17'd21519,17'd21520,17'd21521,17'd21522,17'd21523,17'd21524,17'd21525,17'd21526,17'd21527,17'd21528,17'd21529,17'd21530,17'd21531,17'd21532,17'd21533,17'd21534,17'd21535,17'd21536,17'd21537,17'd21538,17'd21539,17'd21540,17'd21541,17'd21542,17'd21543,17'd21544,17'd21545,17'd21546,17'd21547,17'd21548,17'd21549,17'd21550,17'd21551,17'd21552,17'd21553,17'd21554,17'd21555,17'd21097,17'd21556,17'd21557,17'd21558,17'd21559,17'd21560,17'd21561,17'd21562,17'd21563,17'd21564,17'd21565,17'd20346,17'd21566,17'd21567,17'd21264,17'd18943,17'd21568,17'd21569,17'd21570,17'd21571,17'd21419,17'd21572,17'd21573,17'd21574,17'd21575,17'd21576,17'd20502,17'd20811,17'd21577,17'd20811,17'd20815,17'd21275,17'd20360,17'd21427,17'd20817,17'd20364,17'd21578,17'd21579,17'd21580,17'd21581,17'd21582,17'd21279,17'd21583,17'd21122,17'd21584,17'd21282,17'd21434,17'd21585,17'd21586,17'd21587,17'd21588,17'd21589,17'd21590,17'd21591,17'd21592,17'd21593,17'd21594,17'd21595,17'd21596,17'd20679,17'd21597,17'd21598,17'd21599,17'd21600,17'd21601,17'd21602,17'd21603,17'd21603,17'd21604,17'd21605,17'd21136,17'd21606,17'd21607,17'd21608,17'd21609,17'd21610,17'd21611,17'd20842,17'd21612,17'd21613,17'd21305,17'd21306,17'd20536,17'd21307,17'd20694,17'd21001,17'd21001,17'd16121,17'd16121,17'd16247,17'd16371,17'd15724,17'd17282,17'd17063,17'd16844,17'd16246,17'd16118,17'd15852,17'd15723,17'd15605,17'd15093,17'd21001,17'd18022,17'd21614,17'd21615,17'd20117,17'd20699,17'd11436,17'd21616,17'd21617,17'd19854,17'd20553,17'd18977,17'd19721,17'd21618,17'd21619,17'd21318,17'd21620,17'd21621,17'd21622,17'd21623,17'd21624,17'd927,17'd18514,17'd621,17'd967,17'd19603,17'd21625,17'd6252,17'd2759,17'd21470,17'd6249,17'd4871,17'd8490,17'd8318,17'd11189,17'd9252,17'd9535,17'd9255,17'd11724,17'd11874,17'd11192,17'd11192,17'd9948,17'd11192,17'd20715,17'd21626,17'd21627,17'd21627,17'd9406,17'd8956,17'd20716,17'd9794,17'd21628,17'd21163,17'd21163,17'd21163,17'd11053,17'd8647,17'd10390,17'd21327,17'd21629,17'd4411,17'd20717,17'd6876,17'd6877,17'd7040,17'd7201,17'd5048,17'd4417,17'd2110,17'd964,17'd15741,17'd17552,17'd21630
},
'{
17'd466,17'd2,17'd0,17'd0,17'd12,17'd12,17'd2423,17'd2423,17'd21,17'd4,17'd6,17'd7,17'd8190,17'd8190,17'd8340,17'd10795,17'd8340,17'd8340,17'd8040,17'd8040,17'd5205,17'd3753,17'd6,17'd5,17'd24,17'd24,17'd24,17'd24,17'd24,17'd284,17'd5,17'd7,17'd3753,17'd3753,17'd7554,17'd7383,17'd21631,17'd7061,17'd18037,17'd3907,17'd11208,17'd2430,17'd1838,17'd21632,17'd59,17'd14871,17'd21473,17'd21633,17'd21634,17'd21635,17'd21636,17'd21637,17'd21638,17'd21639,17'd21640,17'd2627,17'd5530,17'd21641,17'd21642,17'd21643,17'd21644,17'd21645,17'd12940,17'd10556,17'd20287,17'd20582,17'd21646,17'd21342,17'd21647,17'd21648,17'd20884,17'd20147,17'd14764,17'd12530,17'd12361,17'd12361,17'd12362,17'd13094,17'd12679,17'd19127,17'd13092,17'd13092,17'd12678,17'd13092,17'd12955,17'd15137,17'd15137,17'd12360,17'd12218,17'd12530,17'd12361,17'd12361,17'd12532,17'd12532,17'd19006,17'd19006,17'd19620,17'd21649,17'd21650,17'd17319,17'd18060,17'd18658,17'd21651,17'd21186,17'd20586,17'd18659,17'd21652,17'd21653,17'd21654,17'd21654,17'd8217,17'd12816,17'd8844,17'd9843,17'd9705,17'd9845,17'd9705,17'd9705,17'd9705,17'd9705,17'd10566,17'd11765,17'd11235,17'd11235,17'd11917,17'd21655,17'd21656,17'd21657,17'd21490,17'd21658,17'd21193,17'd18310,17'd21492,17'd21659,17'd16297,17'd13858,17'd21660,17'd21661,17'd21662,17'd13749,17'd11649,17'd21497,17'd20898,17'd21498,17'd13637,17'd21663,17'd21664,17'd20900,17'd13131,17'd21665,17'd21666,17'd21667,17'd21668,17'd12857,17'd10737,17'd17124,17'd9342,17'd16793,17'd16328,17'd21669,17'd15943,17'd10991,17'd10739,17'd10990,17'd13516,17'd16326,17'd13883,17'd12578,17'd12418,17'd12416,17'd12416,17'd12415,17'd18564,17'd12254,17'd19407,17'd17348,17'd17722,17'd16326,17'd13645,17'd11964,17'd15185,17'd16325,17'd21363,17'd21505,17'd21505,17'd21361,17'd16204,17'd17968,17'd21670,17'd18330,17'd12858,17'd12995,17'd14526,17'd14809,17'd12856,17'd12109,17'd13882,17'd15184,17'd21671,17'd17348,17'd14807,17'd12579,17'd12419,17'd16064,17'd10477,17'd9346,17'd8882,17'd8730,17'd9744,17'd17849,17'd15188,17'd14937,17'd14937,17'd15439,17'd9891,17'd10343,17'd21672,17'd21673,17'd21674,17'd7956,17'd21675,17'd9748,17'd21676,17'd21677,17'd21678,17'd16217,17'd7812,17'd21679,17'd17363,17'd133,17'd132,17'd132,17'd5593,17'd5593,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd5593,17'd131,17'd11541,17'd131,17'd134,17'd134,17'd130,17'd128,17'd133,17'd21680,17'd21681,17'd21682,17'd21683,17'd21684,17'd21685,17'd21686,17'd21687,17'd21688,17'd21689,17'd21690,17'd21691,17'd21692,17'd21693,17'd21694,17'd21694,17'd21695,17'd21696,17'd21697,17'd21698,17'd21699,17'd21700,17'd21701,17'd21702,17'd21703,17'd21704,17'd21705,17'd21706,17'd21707,17'd21708,17'd21709,17'd21710,17'd21711,17'd21712,17'd21713,17'd21714,17'd21715,17'd21716,17'd21717,17'd21718,17'd21719,17'd21720,17'd21721,17'd21722,17'd21723,17'd21724,17'd20205,17'd21725,17'd21726,17'd21727,17'd21728,17'd21729,17'd20207,17'd21730,17'd21731,17'd21732,17'd19055,17'd21569,17'd21733,17'd21734,17'd21735,17'd21736,17'd20802,17'd21574,17'd21737,17'd20661,17'd20502,17'd21738,17'd20811,17'd21739,17'd21740,17'd20667,17'd21426,17'd20816,17'd20228,17'd21741,17'd21578,17'd21742,17'd20825,17'd21278,17'd20977,17'd21279,17'd21743,17'd21744,17'd21434,17'd21434,17'd21437,17'd21592,17'd21591,17'd21745,17'd21746,17'd21747,17'd21748,17'd21747,17'd21749,17'd21590,17'd21750,17'd21751,17'd21752,17'd21753,17'd21754,17'd20519,17'd20519,17'd21755,17'd21756,17'd21757,17'd21758,17'd21759,17'd21760,17'd21761,17'd21762,17'd21763,17'd21764,17'd21765,17'd21608,17'd21452,17'd21766,17'd11159,17'd21767,17'd21768,17'd20995,17'd21769,17'd21770,17'd20998,17'd20539,17'd20694,17'd20540,17'd21309,17'd21453,17'd16247,17'd17065,17'd17065,17'd17065,17'd20542,17'd21771,17'd21772,17'd21772,17'd15852,17'd15604,17'd15724,17'd15093,17'd21001,17'd18260,17'd21773,17'd21774,17'd21775,17'd21776,17'd21777,17'd11437,17'd20701,17'd21778,17'd19352,17'd18750,17'd12314,17'd19723,17'd21779,17'd3692,17'd21780,17'd21781,17'd21782,17'd21783,17'd21784,17'd21785,17'd18514,17'd635,17'd594,17'd21161,17'd21786,17'd6578,17'd2403,17'd21787,17'd4563,17'd8318,17'd9116,17'd8318,17'd9116,17'd8794,17'd9535,17'd9255,17'd11329,17'd11874,17'd9256,17'd10249,17'd9948,17'd9948,17'd20715,17'd12024,17'd8490,17'd8955,17'd8798,17'd21788,17'd8799,17'd8956,17'd9406,17'd21472,17'd21472,17'd12321,17'd9950,17'd9797,17'd8490,17'd4718,17'd4721,17'd4412,17'd20717,17'd21789,17'd21790,17'd7040,17'd7201,17'd3417,17'd4417,17'd21791,17'd20271,17'd17422,17'd17075,17'd21630
},
'{
17'd466,17'd2,17'd0,17'd0,17'd12,17'd12,17'd2423,17'd2423,17'd25,17'd4,17'd6,17'd7,17'd8190,17'd8190,17'd8340,17'd10795,17'd8040,17'd8040,17'd8040,17'd8040,17'd3753,17'd3753,17'd5,17'd5,17'd24,17'd284,17'd284,17'd24,17'd5,17'd5,17'd5,17'd6,17'd3594,17'd5,17'd7383,17'd1691,17'd7385,17'd7060,17'd4431,17'd9816,17'd12036,17'd14446,17'd1134,17'd1555,17'd59,17'd14871,17'd21473,17'd21633,17'd21792,17'd21635,17'd21793,17'd21794,17'd21795,17'd21796,17'd21797,17'd21798,17'd21799,17'd21800,17'd21801,17'd21802,17'd21803,17'd19748,17'd21804,17'd21805,17'd20287,17'd20145,17'd13827,17'd21181,17'd21806,17'd21807,17'd21036,17'd14622,17'd12530,17'd12530,17'd12361,17'd12361,17'd12362,17'd13094,17'd12679,17'd19127,17'd13092,17'd13092,17'd13092,17'd13093,17'd14890,17'd15137,17'd12360,17'd12360,17'd12530,17'd12530,17'd13969,17'd12361,17'd12531,17'd20886,17'd19006,17'd18774,17'd17206,17'd21808,17'd16164,17'd16519,17'd18060,17'd18658,17'd21651,17'd6299,17'd21809,17'd20736,17'd8214,17'd21810,17'd8215,17'd8215,17'd13213,17'd7414,17'd10119,17'd9843,17'd9705,17'd9705,17'd9705,17'd9705,17'd9705,17'd10120,17'd11765,17'd11765,17'd11235,17'd11766,17'd11917,17'd21655,17'd21656,17'd20891,17'd21658,17'd20162,17'd21193,17'd18311,17'd20164,17'd21350,17'd15919,17'd10705,17'd21811,17'd21812,17'd21813,17'd12395,17'd12712,17'd21201,17'd21814,17'd20306,17'd13130,17'd21815,17'd21664,17'd13359,17'd18676,17'd21816,17'd21817,17'd21818,17'd21819,17'd11807,17'd10326,17'd21820,17'd21821,17'd9339,17'd18556,17'd11401,17'd12863,17'd11132,17'd10854,17'd11808,17'd18444,17'd15053,17'd12109,17'd15434,17'd12416,17'd12416,17'd12415,17'd12415,17'd18564,17'd12254,17'd19407,17'd20314,17'd18443,17'd18444,17'd18444,17'd19158,17'd16325,17'd21361,17'd21363,17'd21505,17'd21361,17'd18443,17'd12115,17'd18682,17'd21822,17'd18447,17'd11958,17'd13517,17'd21207,17'd14526,17'd12995,17'd12109,17'd13882,17'd18565,17'd14130,17'd21671,17'd16203,17'd13882,17'd18679,17'd17121,17'd10856,17'd15682,17'd8724,17'd9047,17'd21823,17'd21824,17'd15693,17'd14937,17'd15193,17'd7620,17'd14678,17'd21825,17'd21826,17'd21827,17'd15573,17'd21828,17'd21829,17'd19538,17'd21830,17'd21831,17'd21832,17'd21833,17'd7979,17'd7980,17'd17363,17'd133,17'd11541,17'd134,17'd131,17'd131,17'd132,17'd132,17'd134,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd5593,17'd20466,17'd131,17'd131,17'd11541,17'd132,17'd20623,17'd21834,17'd21835,17'd21836,17'd21522,17'd21837,17'd21838,17'd21535,17'd21839,17'd21690,17'd21840,17'd21841,17'd21842,17'd21843,17'd21844,17'd21845,17'd21845,17'd21846,17'd21845,17'd21847,17'd21844,17'd21848,17'd21849,17'd21850,17'd21851,17'd21852,17'd21853,17'd21854,17'd21855,17'd21856,17'd21857,17'd21858,17'd21859,17'd21860,17'd21861,17'd21862,17'd21863,17'd21864,17'd21865,17'd21866,17'd21867,17'd21868,17'd21408,17'd21869,17'd21870,17'd21871,17'd21872,17'd21873,17'd21874,17'd21875,17'd21876,17'd21877,17'd21878,17'd21879,17'd21880,17'd21881,17'd18592,17'd21882,17'd21883,17'd21884,17'd21885,17'd21886,17'd21735,17'd21887,17'd20960,17'd21888,17'd21889,17'd21890,17'd20812,17'd21274,17'd20811,17'd21275,17'd21740,17'd20360,17'd21426,17'd20816,17'd20228,17'd21741,17'd21891,17'd21892,17'd21893,17'd21582,17'd21894,17'd21124,17'd21895,17'd21896,17'd21897,17'd21898,17'd21899,17'd21900,17'd21901,17'd21902,17'd21903,17'd21904,17'd21905,17'd21906,17'd21907,17'd21908,17'd21909,17'd21910,17'd21911,17'd21912,17'd21596,17'd21754,17'd20519,17'd21913,17'd21914,17'd21756,17'd21915,17'd21916,17'd21917,17'd21918,17'd21919,17'd21920,17'd21606,17'd21921,17'd21922,17'd21923,17'd21924,17'd21925,17'd21926,17'd21927,17'd21928,17'd21929,17'd20535,17'd21770,17'd20999,17'd20846,17'd20694,17'd21309,17'd21309,17'd16121,17'd16371,17'd17065,17'd17065,17'd17903,17'd21930,17'd21772,17'd21772,17'd15852,17'd15604,17'd15724,17'd15093,17'd20695,17'd18620,17'd21931,17'd15478,17'd21932,17'd21933,17'd21934,17'd21935,17'd21936,17'd21778,17'd20855,17'd21937,17'd20553,17'd20120,17'd10243,17'd21938,17'd21939,17'd21940,17'd21941,17'd21942,17'd21943,17'd21159,17'd21944,17'd635,17'd404,17'd8483,17'd21945,17'd6252,17'd2402,17'd21470,17'd4563,17'd9116,17'd9116,17'd9116,17'd5034,17'd21946,17'd9535,17'd9254,17'd10078,17'd9256,17'd20566,17'd20716,17'd20714,17'd20716,17'd21947,17'd21948,17'd8318,17'd8796,17'd8955,17'd8798,17'd21019,17'd9536,17'd21947,17'd21472,17'd21472,17'd21472,17'd9797,17'd9797,17'd8490,17'd4718,17'd3233,17'd3578,17'd3723,17'd21789,17'd21790,17'd7040,17'd7526,17'd4079,17'd3737,17'd21791,17'd279,17'd15492,17'd179,17'd17552
},
'{
17'd2,17'd2,17'd2,17'd2,17'd2,17'd13,17'd2423,17'd16747,17'd23,17'd4,17'd6,17'd5205,17'd8340,17'd8340,17'd8190,17'd8190,17'd8040,17'd8040,17'd5205,17'd3753,17'd3753,17'd3594,17'd24,17'd24,17'd5,17'd284,17'd284,17'd24,17'd6,17'd6,17'd5,17'd5,17'd5,17'd5,17'd7384,17'd1691,17'd7385,17'd6744,17'd3907,17'd11208,17'd2264,17'd1972,17'd21949,17'd56,17'd20869,17'd14750,17'd21950,17'd21951,17'd1985,17'd21952,17'd21953,17'd21954,17'd21955,17'd21956,17'd3928,17'd13075,17'd21957,17'd12795,17'd21958,17'd21959,17'd21960,17'd13080,17'd12941,17'd17090,17'd21961,17'd13828,17'd17091,17'd21343,17'd21648,17'd21962,17'd21963,17'd14622,17'd12530,17'd12530,17'd12530,17'd12530,17'd14621,17'd12955,17'd12679,17'd12527,17'd14469,17'd13092,17'd12679,17'd12955,17'd14890,17'd12530,17'd12530,17'd12530,17'd12530,17'd13840,17'd13969,17'd12361,17'd20424,17'd20886,17'd17941,17'd19511,17'd21964,17'd19384,17'd17319,17'd16519,17'd16028,17'd21965,17'd21966,17'd17097,17'd7247,17'd21967,17'd21968,17'd21968,17'd21969,17'd21969,17'd8366,17'd7414,17'd10119,17'd9843,17'd9705,17'd9705,17'd9843,17'd9705,17'd10120,17'd10120,17'd12068,17'd12068,17'd21970,17'd21971,17'd21655,17'd21656,17'd20742,17'd20741,17'd21193,17'd21193,17'd20745,17'd18788,17'd18067,17'd16297,17'd21972,17'd21973,17'd21974,17'd21975,17'd16429,17'd12093,17'd21976,17'd21977,17'd20445,17'd21978,17'd12235,17'd21979,17'd15676,17'd21980,17'd21497,17'd21359,17'd20447,17'd21981,17'd21982,17'd10990,17'd9473,17'd21983,17'd21984,17'd15187,17'd12585,17'd15176,17'd19282,17'd11132,17'd10854,17'd11965,17'd16204,17'd13761,17'd12578,17'd12418,17'd12416,17'd21504,17'd12415,17'd12415,17'd15434,17'd12579,17'd19408,17'd17722,17'd18444,17'd21985,17'd16326,17'd16442,17'd20314,17'd20314,17'd20314,17'd19408,17'd16442,17'd16326,17'd11965,17'd18682,17'd18683,17'd12113,17'd13252,17'd13517,17'd13515,17'd15570,17'd12580,17'd12419,17'd13761,17'd13883,17'd11959,17'd15184,17'd15184,17'd19645,17'd21986,17'd10164,17'd21983,17'd15297,17'd8730,17'd21987,17'd17849,17'd16691,17'd21988,17'd16447,17'd14680,17'd15058,17'd12868,17'd18922,17'd21989,17'd21990,17'd21991,17'd21828,17'd21060,17'd21992,17'd21993,17'd21994,17'd11005,17'd15701,17'd21995,17'd11977,17'd14275,17'd11289,17'd889,17'd133,17'd133,17'd1197,17'd1197,17'd1197,17'd128,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd133,17'd15823,17'd21375,17'd20629,17'd21996,17'd21997,17'd21998,17'd21838,17'd21999,17'd22000,17'd22001,17'd22002,17'd22003,17'd22004,17'd22005,17'd21844,17'd22006,17'd22007,17'd22008,17'd22006,17'd21847,17'd22005,17'd22009,17'd22010,17'd22010,17'd22011,17'd22012,17'd22012,17'd21850,17'd22013,17'd22014,17'd22015,17'd22016,17'd22017,17'd22018,17'd22019,17'd22020,17'd22021,17'd22022,17'd22023,17'd22024,17'd22025,17'd22026,17'd22027,17'd21555,17'd22028,17'd22029,17'd22030,17'd22031,17'd22032,17'd22033,17'd20204,17'd22034,17'd22035,17'd22036,17'd22037,17'd22038,17'd22039,17'd22040,17'd18714,17'd22041,17'd22042,17'd22043,17'd22044,17'd22045,17'd22046,17'd22047,17'd22048,17'd22049,17'd22050,17'd21890,17'd20967,17'd22051,17'd20966,17'd21275,17'd21115,17'd20507,17'd21426,17'd20816,17'd20227,17'd20365,17'd22052,17'd22053,17'd21893,17'd22054,17'd21441,17'd22055,17'd21286,17'd22056,17'd22057,17'd22058,17'd22059,17'd22060,17'd22061,17'd22062,17'd22063,17'd22064,17'd22065,17'd22066,17'd22066,17'd22067,17'd22068,17'd22069,17'd22070,17'd22071,17'd21912,17'd21596,17'd22072,17'd22073,17'd22074,17'd22075,17'd22075,17'd22076,17'd22077,17'd21760,17'd21918,17'd21762,17'd22078,17'd22079,17'd22080,17'd22081,17'd22082,17'd22083,17'd11014,17'd22084,17'd22085,17'd21145,17'd22086,17'd20535,17'd20998,17'd22087,17'd20694,17'd21453,17'd21309,17'd15988,17'd16247,17'd16371,17'd17065,17'd17903,17'd20542,17'd22088,17'd18021,17'd16843,17'd17283,17'd17282,17'd15605,17'd16247,17'd18620,17'd22089,17'd21614,17'd15227,17'd22090,17'd22091,17'd9241,17'd10646,17'd22092,17'd20120,17'd19352,17'd18860,17'd20120,17'd19596,17'd22093,17'd22094,17'd22095,17'd22096,17'd22097,17'd22098,17'd22099,17'd1809,17'd621,17'd430,17'd22100,17'd22101,17'd21162,17'd22102,17'd21470,17'd3718,17'd5034,17'd4718,17'd4871,17'd4562,17'd8168,17'd8797,17'd11593,17'd10527,17'd9537,17'd9796,17'd9796,17'd20716,17'd20716,17'd9535,17'd22103,17'd9116,17'd8171,17'd8172,17'd22104,17'd8493,17'd10526,17'd21947,17'd21472,17'd21472,17'd21472,17'd9797,17'd8804,17'd8490,17'd4718,17'd3233,17'd3578,17'd3723,17'd21789,17'd21790,17'd7040,17'd7526,17'd4079,17'd4080,17'd22105,17'd22106,17'd180,17'd15355,17'd17075
},
'{
17'd2,17'd2,17'd2,17'd466,17'd466,17'd2,17'd12,17'd8814,17'd23,17'd5,17'd3753,17'd5205,17'd8340,17'd8340,17'd8190,17'd8190,17'd8340,17'd8040,17'd5205,17'd3753,17'd3594,17'd3594,17'd24,17'd24,17'd24,17'd284,17'd284,17'd5,17'd6,17'd5,17'd5,17'd5,17'd5,17'd23,17'd1691,17'd467,17'd7061,17'd6744,17'd3755,17'd3431,17'd2263,17'd1971,17'd989,17'd820,17'd21329,17'd14750,17'd21950,17'd22107,17'd1985,17'd22108,17'd22109,17'd22110,17'd22111,17'd22112,17'd22113,17'd12511,17'd22114,17'd12795,17'd22115,17'd21482,17'd20419,17'd12798,17'd12941,17'd13588,17'd22116,17'd18165,17'd20583,17'd21806,17'd21807,17'd22117,17'd16027,17'd14622,17'd12530,17'd12530,17'd12530,17'd12218,17'd12955,17'd13093,17'd12679,17'd12527,17'd12357,17'd13209,17'd12955,17'd14890,17'd12218,17'd12218,17'd12530,17'd12530,17'd12530,17'd12530,17'd13969,17'd16765,17'd20886,17'd17317,17'd17689,17'd17206,17'd20735,17'd18060,17'd17320,17'd16519,17'd15645,17'd22118,17'd21966,17'd17323,17'd6768,17'd22119,17'd22120,17'd21810,17'd9439,17'd9439,17'd8366,17'd7749,17'd10119,17'd9843,17'd9843,17'd9843,17'd9843,17'd9843,17'd10120,17'd10120,17'd11765,17'd12068,17'd21970,17'd11917,17'd13610,17'd21657,17'd20742,17'd20741,17'd21193,17'd20034,17'd19269,17'd22121,17'd22122,17'd15788,17'd10440,17'd22123,17'd22124,17'd22125,17'd12237,17'd22126,17'd22127,17'd22128,17'd22129,17'd20753,17'd12235,17'd17593,17'd13131,17'd22126,17'd11946,17'd20171,17'd22130,17'd16313,17'd17121,17'd10479,17'd9338,17'd17840,17'd9346,17'd22131,17'd11527,17'd21206,17'd11132,17'd11131,17'd11129,17'd13516,17'd13883,17'd12414,17'd12418,17'd14003,17'd21504,17'd19534,17'd12415,17'd18564,17'd12253,17'd14130,17'd17722,17'd16442,17'd19643,17'd21985,17'd18443,17'd21361,17'd20314,17'd20314,17'd19408,17'd11959,17'd15185,17'd11964,17'd11965,17'd10989,17'd11963,17'd12857,17'd13252,17'd15433,17'd13517,17'd17348,17'd12420,17'd12419,17'd11960,17'd13883,17'd11959,17'd13882,17'd18565,17'd22132,17'd14666,17'd10857,17'd16910,17'd8567,17'd8571,17'd9745,17'd17352,17'd17016,17'd22133,17'd22134,17'd22135,17'd8427,17'd13529,17'd22136,17'd22137,17'd22138,17'd20613,17'd22139,17'd22140,17'd22141,17'd22142,17'd22143,17'd22144,17'd13533,17'd22145,17'd22146,17'd15821,17'd22147,17'd8444,17'd17363,17'd8132,17'd542,17'd542,17'd133,17'd133,17'd128,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd134,17'd16090,17'd20623,17'd22148,17'd22149,17'd22150,17'd22151,17'd22152,17'd22153,17'd22154,17'd21697,17'd22004,17'd22155,17'd22156,17'd22157,17'd22158,17'd22159,17'd22160,17'd22160,17'd22161,17'd22162,17'd22156,17'd22163,17'd22164,17'd22165,17'd22005,17'd22009,17'd22166,17'd22167,17'd22168,17'd22167,17'd22011,17'd22169,17'd22170,17'd22171,17'd22172,17'd22173,17'd22174,17'd22175,17'd22176,17'd22177,17'd22178,17'd22179,17'd22180,17'd22181,17'd22182,17'd22183,17'd22184,17'd22030,17'd22185,17'd22186,17'd21722,17'd22187,17'd22188,17'd22189,17'd22190,17'd22191,17'd22192,17'd22193,17'd22194,17'd22195,17'd22196,17'd22197,17'd22198,17'd22199,17'd22200,17'd21886,17'd22201,17'd21110,17'd22202,17'd22203,17'd22204,17'd22205,17'd22206,17'd20966,17'd21275,17'd20225,17'd20507,17'd21426,17'd20816,17'd20229,17'd20516,17'd22207,17'd22208,17'd22209,17'd22210,17'd21287,17'd21286,17'd22211,17'd22212,17'd22213,17'd22214,17'd22215,17'd22216,17'd22217,17'd22218,17'd22219,17'd22220,17'd22221,17'd22222,17'd22222,17'd22223,17'd22067,17'd22224,17'd22225,17'd22226,17'd22227,17'd22228,17'd22229,17'd22230,17'd22231,17'd22232,17'd22233,17'd22234,17'd22235,17'd22236,17'd22237,17'd22238,17'd22239,17'd22079,17'd22240,17'd22241,17'd22242,17'd22243,17'd22244,17'd22245,17'd22246,17'd22247,17'd21145,17'd22248,17'd22249,17'd20537,17'd20846,17'd21453,17'd21309,17'd15607,17'd15988,17'd16371,17'd17065,17'd17779,17'd17903,17'd22250,17'd18021,17'd16843,17'd16843,17'd17282,17'd15724,17'd16371,17'd18741,17'd22251,17'd22252,17'd14852,17'd16489,17'd22253,17'd11858,17'd22254,17'd12170,17'd22255,17'd20553,17'd18748,17'd22256,17'd20121,17'd22257,17'd22258,17'd22259,17'd22260,17'd22261,17'd22262,17'd20263,17'd22263,17'd22264,17'd611,17'd187,17'd22101,17'd21326,17'd8487,17'd2571,17'd13291,17'd4562,17'd4719,17'd4562,17'd22265,17'd8167,17'd8796,17'd10077,17'd9255,17'd12919,17'd21163,17'd21163,17'd21628,17'd21628,17'd22266,17'd8167,17'd4872,17'd8018,17'd8171,17'd11592,17'd8955,17'd9946,17'd9535,17'd21472,17'd9535,17'd21472,17'd9797,17'd9251,17'd11189,17'd4871,17'd4568,17'd3578,17'd3723,17'd21789,17'd21790,17'd6882,17'd7202,17'd4417,17'd21791,17'd22105,17'd22267,17'd252,17'd20720,17'd21165
},
'{
17'd13,17'd13,17'd466,17'd466,17'd466,17'd13,17'd2423,17'd8814,17'd4,17'd5,17'd3753,17'd8040,17'd8340,17'd8340,17'd8190,17'd8190,17'd8340,17'd8340,17'd5205,17'd3753,17'd3753,17'd3594,17'd24,17'd24,17'd284,17'd284,17'd5,17'd6,17'd5,17'd24,17'd22268,17'd5,17'd5,17'd23,17'd1691,17'd285,17'd7061,17'd18037,17'd3754,17'd12036,17'd1973,17'd1837,17'd821,17'd58,17'd61,17'd64,17'd22269,17'd22270,17'd18636,17'd22271,17'd22272,17'd22273,17'd2959,17'd22274,17'd22275,17'd22276,17'd22277,17'd22278,17'd21643,17'd22279,17'd19748,17'd22280,17'd22281,17'd22282,17'd22116,17'd13827,17'd22283,17'd20733,17'd20734,17'd21036,17'd14622,17'd12361,17'd12530,17'd12530,17'd14890,17'd14890,17'd12528,17'd12679,17'd12527,17'd12527,17'd14469,17'd16284,17'd12528,17'd14890,17'd12218,17'd12956,17'd12680,17'd11913,17'd12530,17'd12218,17'd12362,17'd12361,17'd12532,17'd17204,17'd17689,17'd21649,17'd19384,17'd15899,17'd16034,17'd16769,17'd21965,17'd16522,17'd16770,17'd17323,17'd21186,17'd11088,17'd22284,17'd21968,17'd9439,17'd9439,17'd8684,17'd7749,17'd10119,17'd10119,17'd8844,17'd8844,17'd10119,17'd10119,17'd11916,17'd11916,17'd22285,17'd12961,17'd11766,17'd11917,17'd13610,17'd22286,17'd20742,17'd20299,17'd20034,17'd19268,17'd22121,17'd22287,17'd22288,17'd13615,17'd22289,17'd18315,17'd22290,17'd22291,17'd12406,17'd21201,17'd21048,17'd22292,17'd22293,17'd21663,17'd17593,17'd12087,17'd18676,17'd22294,17'd18801,17'd15044,17'd22295,17'd15186,17'd22296,17'd10742,17'd16793,17'd9339,17'd11809,17'd16070,17'd11132,17'd10854,17'd11131,17'd11131,17'd11129,17'd11807,17'd13761,17'd12414,17'd12417,17'd14003,17'd22297,17'd19534,17'd12415,17'd12254,17'd12579,17'd18198,17'd16442,17'd16326,17'd18444,17'd18681,17'd18197,17'd18559,17'd17474,17'd17474,17'd11959,17'd11960,17'd19158,17'd13516,17'd13645,17'd12262,17'd12113,17'd12419,17'd12995,17'd15685,17'd12580,17'd16321,17'd12420,17'd12857,17'd12857,17'd12113,17'd11960,17'd15054,17'd14669,17'd17838,17'd12116,17'd21984,17'd8567,17'd10607,17'd18808,17'd22298,17'd17850,17'd12265,17'd13376,17'd14681,17'd17018,17'd22299,17'd22300,17'd7625,17'd7956,17'd22301,17'd19647,17'd22302,17'd22303,17'd15310,17'd22304,17'd22305,17'd22306,17'd22307,17'd10037,17'd10189,17'd22308,17'd22309,17'd20463,17'd22146,17'd20621,17'd22310,17'd22311,17'd14276,17'd542,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd720,17'd4163,17'd11413,17'd22312,17'd22313,17'd22314,17'd22315,17'd22316,17'd22317,17'd22318,17'd22319,17'd22320,17'd22321,17'd22322,17'd22323,17'd22324,17'd22325,17'd22326,17'd22327,17'd22328,17'd22329,17'd22330,17'd22331,17'd22332,17'd22332,17'd22333,17'd22334,17'd22334,17'd22159,17'd22158,17'd22157,17'd22335,17'd22336,17'd21696,17'd22337,17'd22338,17'd22339,17'd22340,17'd22341,17'd22342,17'd22343,17'd22344,17'd22345,17'd22346,17'd22347,17'd22348,17'd22349,17'd22350,17'd22351,17'd22352,17'd22353,17'd22354,17'd22355,17'd22356,17'd22357,17'd22358,17'd22359,17'd22360,17'd22361,17'd22362,17'd22363,17'd22364,17'd22194,17'd22365,17'd22366,17'd22367,17'd22368,17'd22369,17'd22045,17'd22370,17'd22371,17'd22372,17'd22373,17'd22374,17'd22375,17'd22376,17'd20664,17'd21740,17'd22377,17'd22378,17'd20507,17'd20968,17'd20227,17'd22379,17'd22380,17'd21892,17'd22381,17'd20979,17'd22382,17'd22383,17'd22384,17'd22234,17'd22385,17'd22386,17'd22387,17'd22388,17'd22389,17'd22390,17'd22218,17'd22391,17'd22392,17'd22392,17'd22223,17'd22222,17'd22393,17'd22394,17'd22395,17'd22396,17'd22397,17'd22398,17'd22399,17'd22230,17'd22400,17'd22401,17'd22402,17'd22403,17'd22404,17'd22405,17'd22406,17'd22407,17'd22408,17'd22409,17'd22410,17'd22411,17'd22242,17'd22412,17'd22413,17'd10627,17'd22414,17'd22246,17'd22415,17'd22086,17'd21147,17'd22416,17'd22417,17'd22418,17'd22419,17'd22420,17'd18742,17'd16247,17'd17065,17'd17779,17'd17903,17'd20542,17'd21930,17'd16843,17'd16842,17'd17901,17'd22421,17'd18619,17'd22422,17'd22423,17'd20544,17'd13408,17'd15343,17'd22424,17'd22425,17'd21935,17'd22426,17'd21316,17'd20854,17'd18265,17'd18859,17'd22427,17'd22428,17'd22429,17'd22430,17'd22431,17'd22432,17'd22433,17'd22434,17'd22435,17'd933,17'd611,17'd20270,17'd22436,17'd9249,17'd3409,17'd2402,17'd13291,17'd4562,17'd4719,17'd4718,17'd19104,17'd5034,17'd8954,17'd10391,17'd9255,17'd12919,17'd21163,17'd21163,17'd22437,17'd21628,17'd22438,17'd5034,17'd4717,17'd14983,17'd9944,17'd22439,17'd7857,17'd11592,17'd8955,17'd8796,17'd9534,17'd8797,17'd11596,17'd7687,17'd7685,17'd6576,17'd7349,17'd3578,17'd3723,17'd22440,17'd22441,17'd22442,17'd22443,17'd22444,17'd22445,17'd22446,17'd22267,17'd252,17'd22447,17'd22448
},
'{
17'd3430,17'd3430,17'd466,17'd466,17'd466,17'd2,17'd12,17'd8814,17'd4,17'd5,17'd3753,17'd8040,17'd8340,17'd8340,17'd8190,17'd8190,17'd8340,17'd8340,17'd5205,17'd3753,17'd3594,17'd3594,17'd24,17'd24,17'd284,17'd24,17'd5,17'd6,17'd5,17'd24,17'd22268,17'd6,17'd4,17'd23,17'd467,17'd286,17'd6902,17'd4431,17'd3255,17'd2942,17'd2121,17'd1700,17'd821,17'd664,17'd14749,17'd14750,17'd21473,17'd22449,17'd18636,17'd22450,17'd22451,17'd22452,17'd14876,17'd22453,17'd22454,17'd22455,17'd22456,17'd22278,17'd22457,17'd20141,17'd12797,17'd22458,17'd13314,17'd18650,17'd18289,17'd13827,17'd22283,17'd22459,17'd22460,17'd18173,17'd14622,17'd12361,17'd12530,17'd12530,17'd14890,17'd12955,17'd12679,17'd12527,17'd12527,17'd12527,17'd16284,17'd13209,17'd12955,17'd12814,17'd12956,17'd11627,17'd12680,17'd12680,17'd12218,17'd12218,17'd12362,17'd12532,17'd17941,17'd18774,17'd21649,17'd20735,17'd16659,17'd16034,17'd15524,17'd17322,17'd21965,17'd22461,17'd22462,17'd6133,17'd20887,17'd20426,17'd22463,17'd22464,17'd13327,17'd9439,17'd8366,17'd7749,17'd10119,17'd8844,17'd8844,17'd8844,17'd10119,17'd10119,17'd11916,17'd11916,17'd22285,17'd12961,17'd11766,17'd11917,17'd22286,17'd21657,17'd20741,17'd20299,17'd19141,17'd19268,17'd20037,17'd22465,17'd22466,17'd9594,17'd19028,17'd10712,17'd22467,17'd16902,17'd22294,17'd22468,17'd20750,17'd21980,17'd20753,17'd22469,17'd12560,17'd18799,17'd18800,17'd22470,17'd22471,17'd14925,17'd21360,17'd14673,17'd12116,17'd9190,17'd15682,17'd14674,17'd14383,17'd11528,17'd10475,17'd10854,17'd11131,17'd11130,17'd13516,17'd11961,17'd12577,17'd12253,17'd12416,17'd12416,17'd22297,17'd19534,17'd18564,17'd12579,17'd11959,17'd16325,17'd18327,17'd21985,17'd18681,17'd22472,17'd18559,17'd20314,17'd17474,17'd16321,17'd13883,17'd13135,17'd13516,17'd13516,17'd18444,17'd15185,17'd11960,17'd12109,17'd12995,17'd13252,17'd11959,17'd11960,17'd12113,17'd12113,17'd12113,17'd12857,17'd11960,17'd15299,17'd13000,17'd12863,17'd9339,17'd8721,17'd22473,17'd9483,17'd22474,17'd8579,17'd17128,17'd7786,17'd16802,17'd22475,17'd22476,17'd22477,17'd22478,17'd22479,17'd22480,17'd22480,17'd22481,17'd19161,17'd22482,17'd22483,17'd22484,17'd22485,17'd22486,17'd11007,17'd11007,17'd22487,17'd22487,17'd15201,17'd22488,17'd13533,17'd22145,17'd17861,17'd22489,17'd15959,17'd14275,17'd17363,17'd133,17'd1045,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd134,17'd16090,17'd20624,17'd22490,17'd22491,17'd22492,17'd22493,17'd22000,17'd22494,17'd22495,17'd22496,17'd22322,17'd22497,17'd22498,17'd22499,17'd22325,17'd22500,17'd22329,17'd22328,17'd22501,17'd22501,17'd22501,17'd22502,17'd22503,17'd22326,17'd22504,17'd22505,17'd22505,17'd22505,17'd22506,17'd22507,17'd22508,17'd22509,17'd22510,17'd22511,17'd22512,17'd22513,17'd22514,17'd22515,17'd22516,17'd22517,17'd22518,17'd22519,17'd22520,17'd22521,17'd22522,17'd22523,17'd22524,17'd22525,17'd22526,17'd22353,17'd22527,17'd22528,17'd22529,17'd22530,17'd22531,17'd22532,17'd22533,17'd22534,17'd22535,17'd22536,17'd22537,17'd22364,17'd22538,17'd22539,17'd22540,17'd22541,17'd22542,17'd22543,17'd22544,17'd22545,17'd22546,17'd22547,17'd22548,17'd22549,17'd22550,17'd22551,17'd22552,17'd22377,17'd22553,17'd20506,17'd20094,17'd20095,17'd22554,17'd22555,17'd20677,17'd22556,17'd20979,17'd21595,17'd22557,17'd22558,17'd22559,17'd22560,17'd22560,17'd22561,17'd22562,17'd22563,17'd22408,17'd22390,17'd22564,17'd22565,17'd22391,17'd22566,17'd22567,17'd22221,17'd22567,17'd22568,17'd22569,17'd22570,17'd22571,17'd22070,17'd22572,17'd22573,17'd22574,17'd22575,17'd22576,17'd22577,17'd22578,17'd22579,17'd22580,17'd22581,17'd22582,17'd22583,17'd22411,17'd22584,17'd22585,17'd22586,17'd22587,17'd22588,17'd22589,17'd22590,17'd21145,17'd22086,17'd22591,17'd22592,17'd22593,17'd21148,17'd17904,17'd18022,17'd16121,17'd16371,17'd17065,17'd17779,17'd17903,17'd17283,17'd16842,17'd16842,17'd22594,17'd17062,17'd17065,17'd18498,17'd19087,17'd22595,17'd13926,17'd15857,17'd22596,17'd19851,17'd21777,17'd12011,17'd22597,17'd13567,17'd22598,17'd18749,17'd13288,17'd22599,17'd22600,17'd22601,17'd22602,17'd22603,17'd22604,17'd22605,17'd22606,17'd431,17'd611,17'd8950,17'd22436,17'd22607,17'd3728,17'd2402,17'd13291,17'd4406,17'd5033,17'd4406,17'd19242,17'd22608,17'd14591,17'd9946,17'd9536,17'd21019,17'd22609,17'd22609,17'd21163,17'd21947,17'd8954,17'd22265,17'd4873,17'd7344,17'd17294,17'd14984,17'd7857,17'd11592,17'd9534,17'd8796,17'd9534,17'd9534,17'd10248,17'd7687,17'd7685,17'd7343,17'd4718,17'd3578,17'd3723,17'd22610,17'd22611,17'd22612,17'd22443,17'd22444,17'd22446,17'd22613,17'd22106,17'd252,17'd22614,17'd22448
},
'{
17'd3430,17'd3430,17'd466,17'd466,17'd466,17'd13,17'd806,17'd2933,17'd4,17'd3753,17'd5793,17'd8040,17'd8340,17'd8340,17'd8190,17'd5205,17'd8040,17'd8040,17'd3753,17'd3753,17'd5,17'd24,17'd24,17'd24,17'd23,17'd23,17'd24,17'd5,17'd5,17'd24,17'd3594,17'd3594,17'd5,17'd23,17'd285,17'd285,17'd7060,17'd4431,17'd3254,17'd3253,17'd22615,17'd1970,17'd821,17'd58,17'd22616,17'd64,17'd22269,17'd22449,17'd18636,17'd1986,17'd16267,17'd22617,17'd3766,17'd22618,17'd22619,17'd22620,17'd22621,17'd22622,17'd22623,17'd20141,17'd12797,17'd12941,17'd22624,17'd22625,17'd13826,17'd17436,17'd22626,17'd22627,17'd22628,17'd18173,17'd14470,17'd12361,17'd12361,17'd12530,17'd14890,17'd12528,17'd19127,17'd12527,17'd12527,17'd15516,17'd22629,17'd16284,17'd12679,17'd12065,17'd12956,17'd11627,17'd12680,17'd12680,17'd12362,17'd12362,17'd12361,17'd22630,17'd19382,17'd18774,17'd16986,17'd16164,17'd16034,17'd16034,17'd22631,17'd22632,17'd15262,17'd5543,17'd16770,17'd16882,17'd20735,17'd22633,17'd22634,17'd12533,17'd9439,17'd9004,17'd7414,17'd7749,17'd8844,17'd8844,17'd22635,17'd8844,17'd10119,17'd10120,17'd11916,17'd11916,17'd22285,17'd12364,17'd11917,17'd21655,17'd21657,17'd21657,17'd20439,17'd20035,17'd22636,17'd18426,17'd20038,17'd22637,17'd21494,17'd22638,17'd22639,17'd22640,17'd12088,17'd12407,17'd22641,17'd21357,17'd22642,17'd15423,17'd18320,17'd12559,17'd12236,17'd12243,17'd13997,17'd15561,17'd22643,17'd22644,17'd11520,17'd13647,17'd13370,17'd22645,17'd17480,17'd22646,17'd21669,17'd11527,17'd10739,17'd20910,17'd22647,17'd11808,17'd11667,17'd13364,17'd12413,17'd12578,17'd12418,17'd14525,17'd22297,17'd22297,17'd12416,17'd14807,17'd18198,17'd18443,17'd21985,17'd21985,17'd14258,17'd21362,17'd20314,17'd19408,17'd14807,17'd12420,17'd12858,17'd12262,17'd11965,17'd13516,17'd19158,17'd18198,17'd16321,17'd12580,17'd13136,17'd13136,17'd13883,17'd13883,17'd12113,17'd12260,17'd14002,17'd12111,17'd11960,17'd13646,17'd11398,17'd10024,17'd9043,17'd8567,17'd8574,17'd14812,17'd10339,17'd8578,17'd22648,17'd7788,17'd19781,17'd22649,17'd22650,17'd22651,17'd14270,17'd22652,17'd22653,17'd22654,17'd22655,17'd22656,17'd22657,17'd22658,17'd13897,17'd17360,17'd22659,17'd22660,17'd17245,17'd22661,17'd22662,17'd22662,17'd10755,17'd17860,17'd11007,17'd10491,17'd10621,17'd12274,17'd22663,17'd22663,17'd22664,17'd15823,17'd11541,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd20762,17'd11413,17'd22665,17'd22666,17'd22667,17'd21382,17'd22668,17'd22669,17'd22670,17'd22671,17'd22335,17'd22672,17'd22673,17'd22674,17'd22675,17'd22676,17'd22505,17'd22333,17'd22677,17'd22332,17'd22678,17'd22679,17'd22679,17'd22680,17'd22327,17'd22325,17'd22681,17'd22334,17'd22682,17'd22682,17'd22683,17'd22156,17'd22684,17'd22685,17'd22686,17'd22687,17'd22688,17'd22689,17'd22690,17'd22691,17'd22692,17'd22693,17'd22694,17'd22695,17'd22696,17'd22697,17'd22698,17'd22699,17'd22700,17'd22701,17'd22526,17'd22353,17'd22527,17'd22702,17'd22703,17'd22704,17'd21723,17'd22705,17'd22706,17'd22707,17'd22708,17'd22709,17'd22710,17'd22711,17'd19671,17'd22539,17'd22712,17'd22713,17'd22714,17'd22715,17'd21734,17'd22716,17'd22717,17'd22718,17'd22719,17'd22720,17'd22721,17'd22722,17'd22552,17'd22377,17'd22553,17'd20667,17'd20094,17'd22723,17'd22724,17'd22555,17'd22725,17'd22726,17'd22727,17'd22728,17'd22729,17'd22730,17'd22731,17'd22732,17'd22732,17'd22733,17'd22734,17'd22735,17'd22736,17'd22737,17'd22738,17'd22739,17'd22218,17'd22740,17'd22220,17'd22567,17'd22741,17'd22221,17'd22742,17'd22742,17'd22740,17'd22743,17'd22744,17'd22212,17'd22745,17'd22746,17'd22747,17'd22748,17'd22749,17'd22750,17'd22751,17'd22752,17'd22753,17'd22754,17'd22755,17'd22756,17'd22757,17'd22758,17'd22759,17'd7824,17'd22760,17'd22761,17'd22415,17'd22762,17'd22763,17'd22764,17'd21148,17'd22765,17'd15340,17'd17904,17'd18742,17'd18620,17'd16371,17'd17779,17'd15724,17'd17282,17'd22594,17'd22766,17'd22594,17'd17062,17'd17065,17'd18498,17'd22767,17'd20543,17'd18971,17'd14425,17'd18744,17'd21776,17'd22768,17'd22769,17'd21617,17'd17540,17'd22770,17'd22771,17'd18750,17'd22772,17'd22773,17'd22774,17'd22775,17'd22776,17'd22777,17'd22778,17'd22435,17'd1822,17'd430,17'd8950,17'd22779,17'd22780,17'd3580,17'd22102,17'd13422,17'd4405,17'd19104,17'd4405,17'd19242,17'd22265,17'd21946,17'd8955,17'd9406,17'd8646,17'd20567,17'd22609,17'd12023,17'd9535,17'd14591,17'd22781,17'd22782,17'd7345,17'd17419,17'd14984,17'd7857,17'd11592,17'd9534,17'd14180,17'd13810,17'd8955,17'd11596,17'd7687,17'd7685,17'd6724,17'd7519,17'd7196,17'd3577,17'd22783,17'd22784,17'd22785,17'd22786,17'd22444,17'd22446,17'd22787,17'd279,17'd180,17'd22788,17'd22448
},
'{
17'd3430,17'd3430,17'd466,17'd466,17'd466,17'd2,17'd3,17'd2933,17'd8,17'd6,17'd3753,17'd8040,17'd8340,17'd8340,17'd8190,17'd5205,17'd8040,17'd5793,17'd3753,17'd3594,17'd5,17'd24,17'd24,17'd24,17'd4,17'd23,17'd284,17'd24,17'd6,17'd5,17'd3594,17'd5,17'd4,17'd23,17'd285,17'd27,17'd6744,17'd3755,17'd2940,17'd2262,17'd22615,17'd1970,17'd1555,17'd58,17'd22616,17'd14750,17'd21473,17'd22449,17'd18636,17'd22789,17'd22790,17'd22791,17'd22792,17'd6609,17'd11895,17'd22793,17'd22794,17'd22795,17'd21340,17'd22796,17'd22797,17'd13314,17'd22798,17'd14088,17'd18527,17'd22799,17'd16877,17'd22800,17'd22801,17'd18173,17'd14470,17'd12361,17'd12361,17'd12218,17'd14890,17'd12528,17'd19127,17'd22802,17'd12527,17'd15516,17'd12528,17'd12679,17'd13093,17'd12065,17'd12218,17'd11627,17'd12680,17'd12957,17'd12362,17'd12361,17'd22630,17'd12681,17'd17689,17'd21649,17'd16164,17'd16519,17'd16169,17'd15902,17'd15770,17'd15010,17'd15262,17'd22461,17'd16770,17'd18658,17'd20735,17'd7083,17'd21967,17'd22634,17'd21969,17'd7414,17'd7414,17'd12816,17'd7749,17'd7748,17'd22635,17'd8844,17'd10119,17'd10120,17'd11916,17'd11480,17'd11765,17'd11766,17'd11917,17'd14229,17'd21657,17'd22803,17'd19762,17'd19141,17'd22804,17'd17459,17'd15919,17'd10439,17'd22805,17'd22806,17'd22807,17'd11786,17'd12402,17'd22294,17'd22808,17'd22809,17'd13504,17'd12087,17'd16790,17'd16790,17'd12568,17'd19639,17'd22810,17'd13360,17'd22811,17'd12999,17'd10990,17'd16912,17'd22812,17'd22813,17'd22814,17'd22815,17'd19642,17'd15176,17'd10854,17'd20451,17'd22816,17'd11807,17'd13364,17'd12413,17'd12578,17'd12859,17'd14525,17'd21057,17'd22297,17'd12416,17'd12253,17'd14130,17'd16325,17'd16326,17'd11397,17'd22817,17'd14258,17'd21362,17'd22818,17'd22819,17'd12579,17'd12419,17'd12114,17'd18682,17'd18682,17'd11964,17'd16325,17'd11959,17'd19408,17'd12106,17'd13519,17'd12259,17'd15053,17'd13883,17'd13135,17'd18328,17'd12858,17'd13363,17'd13366,17'd16069,17'd22820,17'd10025,17'd8873,17'd8728,17'd17481,17'd9196,17'd21987,17'd12119,17'd11968,17'd10746,17'd12727,17'd22821,17'd22822,17'd22823,17'd20613,17'd22824,17'd22825,17'd22826,17'd22827,17'd22828,17'd22829,17'd22830,17'd22831,17'd22832,17'd22833,17'd11681,17'd22834,17'd22835,17'd22836,17'd22835,17'd22837,17'd17614,17'd10350,17'd15313,17'd22838,17'd22839,17'd19542,17'd22840,17'd22841,17'd22842,17'd13777,17'd20466,17'd134,17'd130,17'd130,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd22843,17'd22844,17'd22667,17'd22845,17'd22846,17'd22847,17'd22320,17'd22848,17'd22849,17'd22850,17'd22851,17'd22852,17'd22853,17'd22854,17'd22855,17'd22856,17'd22857,17'd22858,17'd22859,17'd22678,17'd22331,17'd22680,17'd22680,17'd22677,17'd22856,17'd22860,17'd22334,17'd22159,17'd22683,17'd22507,17'd22861,17'd22862,17'd22863,17'd22864,17'd22865,17'd22866,17'd22867,17'd22868,17'd22869,17'd22870,17'd22871,17'd22872,17'd22873,17'd22874,17'd22875,17'd22876,17'd22877,17'd22878,17'd22879,17'd22880,17'd22353,17'd22881,17'd22882,17'd22883,17'd22884,17'd22885,17'd22886,17'd22887,17'd22706,17'd22888,17'd22889,17'd22890,17'd22891,17'd21726,17'd22892,17'd22893,17'd22894,17'd22895,17'd22896,17'd22897,17'd22898,17'd22899,17'd22900,17'd22901,17'd22902,17'd22903,17'd22722,17'd22904,17'd22905,17'd22905,17'd20667,17'd20667,17'd20094,17'd22906,17'd22907,17'd20678,17'd22908,17'd22909,17'd22910,17'd22911,17'd22912,17'd22913,17'd22732,17'd22914,17'd22915,17'd22916,17'd22917,17'd22917,17'd22918,17'd22738,17'd22564,17'd22739,17'd22919,17'd22740,17'd22920,17'd22921,17'd22221,17'd22741,17'd22921,17'd22392,17'd22740,17'd22922,17'd22397,17'd22070,17'd22226,17'd22923,17'd22924,17'd22925,17'd22926,17'd22927,17'd22928,17'd22929,17'd22930,17'd22931,17'd22932,17'd22933,17'd22934,17'd22935,17'd10196,17'd22936,17'd22588,17'd22937,17'd22938,17'd22939,17'd20843,17'd22940,17'd22941,17'd17655,17'd15476,17'd18022,17'd18260,17'd16247,17'd17065,17'd15724,17'd16610,17'd22594,17'd22766,17'd22594,17'd17062,17'd17065,17'd18498,17'd22942,17'd22943,17'd19088,17'd22944,17'd19224,17'd21933,17'd22945,17'd11582,17'd22946,17'd22947,17'd22770,17'd22948,17'd18860,17'd22949,17'd22950,17'd22951,17'd22952,17'd22953,17'd22954,17'd22955,17'd22956,17'd621,17'd442,17'd20270,17'd22957,17'd22958,17'd12638,17'd8487,17'd2248,17'd19104,17'd3878,17'd22781,17'd19242,17'd22265,17'd21946,17'd8796,17'd9535,17'd12023,17'd22959,17'd21626,17'd12024,17'd9535,17'd14590,17'd22960,17'd5503,17'd6723,17'd17073,17'd14984,17'd9405,17'd10076,17'd14062,17'd14180,17'd13810,17'd9534,17'd10248,17'd8490,17'd7685,17'd7343,17'd4718,17'd7519,17'd3577,17'd22610,17'd22961,17'd22785,17'd22786,17'd22962,17'd22613,17'd22963,17'd20271,17'd15626,17'd15355,17'd22964
},
'{
17'd8971,17'd3430,17'd466,17'd466,17'd22965,17'd4089,17'd1128,17'd21,17'd4,17'd3594,17'd5793,17'd8040,17'd8340,17'd8340,17'd5205,17'd5205,17'd8040,17'd8040,17'd3753,17'd3594,17'd24,17'd24,17'd23,17'd4,17'd24,17'd24,17'd3594,17'd3594,17'd5,17'd5,17'd5,17'd24,17'd23,17'd23,17'd467,17'd28,17'd4091,17'd3255,17'd2602,17'd2600,17'd22966,17'd21949,17'd22967,17'd666,17'd482,17'd14603,17'd22968,17'd486,17'd22789,17'd22969,17'd22970,17'd3446,17'd22971,17'd22972,17'd22973,17'd22455,17'd22974,17'd21339,17'd13700,17'd12939,17'd13313,17'd13447,17'd22625,17'd22975,17'd22799,17'd22976,17'd22977,17'd22978,17'd22979,17'd14470,17'd13969,17'd12362,17'd14764,17'd14890,17'd21184,17'd13092,17'd15763,17'd19127,17'd19127,17'd12527,17'd12955,17'd13093,17'd17096,17'd14621,17'd14764,17'd12218,17'd13094,17'd12815,17'd11913,17'd20424,17'd18884,17'd18774,17'd19007,17'd21808,17'd16289,17'd22980,17'd16290,17'd14765,17'd16165,17'd15644,17'd22118,17'd22981,17'd18658,17'd19384,17'd22119,17'd13472,17'd22634,17'd12533,17'd9701,17'd7413,17'd7580,17'd7414,17'd9004,17'd8366,17'd7414,17'd7749,17'd7749,17'd9570,17'd10120,17'd9844,17'd11092,17'd22982,17'd11917,17'd21656,17'd21348,17'd22803,17'd20161,17'd17821,17'd17334,17'd22983,17'd14906,17'd22984,17'd22985,17'd16674,17'd22986,17'd22987,17'd21499,17'd22988,17'd22989,17'd21980,17'd15674,17'd17593,17'd12088,17'd12089,17'd13876,17'd18800,17'd18677,17'd22990,17'd15563,17'd10737,17'd9618,17'd12117,17'd9189,17'd15569,17'd12116,17'd10166,17'd10477,17'd13886,17'd11669,17'd22991,17'd18327,17'd19920,17'd12413,17'd12855,17'd13512,17'd13643,17'd14525,17'd14525,17'd12415,17'd12108,17'd21671,17'd22992,17'd18443,17'd22817,17'd11397,17'd14264,17'd22472,17'd21362,17'd22818,17'd22819,17'd21671,17'd18198,17'd16204,17'd17968,17'd18560,17'd13362,17'd11960,17'd14130,17'd11959,17'd13883,17'd12858,17'd11957,17'd12858,17'd13135,17'd18806,17'd13883,17'd15299,17'd11667,17'd16069,17'd15176,17'd14804,17'd17716,17'd16067,17'd14675,17'd8574,17'd8887,17'd11405,17'd22993,17'd22994,17'd14390,17'd22995,17'd15572,17'd10610,17'd7620,17'd22996,17'd13653,17'd22997,17'd22998,17'd22999,17'd23000,17'd23001,17'd23002,17'd23003,17'd23004,17'd23005,17'd14397,17'd13774,17'd23006,17'd23007,17'd23008,17'd23009,17'd23010,17'd23011,17'd9754,17'd23012,17'd10618,17'd23013,17'd23014,17'd14399,17'd23015,17'd23016,17'd14016,17'd541,17'd20762,17'd20762,17'd1481,17'd11541,17'd131,17'd11541,17'd131,17'd131,17'd11541,17'd132,17'd132,17'd20466,17'd20622,17'd23017,17'd23018,17'd23019,17'd23020,17'd23021,17'd23022,17'd23023,17'd23024,17'd23025,17'd23026,17'd23027,17'd23028,17'd23028,17'd23029,17'd23030,17'd23031,17'd23032,17'd23033,17'd23034,17'd23035,17'd23036,17'd23037,17'd22678,17'd22680,17'd23038,17'd22332,17'd22332,17'd22506,17'd22161,17'd22507,17'd22507,17'd22683,17'd23039,17'd23040,17'd23041,17'd23042,17'd23043,17'd22510,17'd23044,17'd23045,17'd23046,17'd23047,17'd23048,17'd23049,17'd23050,17'd23051,17'd23052,17'd23053,17'd23054,17'd23055,17'd23056,17'd23057,17'd23058,17'd23059,17'd23060,17'd23061,17'd23062,17'd23063,17'd23064,17'd23065,17'd23066,17'd23067,17'd23068,17'd22536,17'd23069,17'd23070,17'd23071,17'd23072,17'd23073,17'd23074,17'd23075,17'd23076,17'd23077,17'd22717,17'd23078,17'd23079,17'd22903,17'd22376,17'd23080,17'd23081,17'd23082,17'd23083,17'd20506,17'd20224,17'd19967,17'd23084,17'd23085,17'd23086,17'd23087,17'd23088,17'd23089,17'd23090,17'd23091,17'd22733,17'd23092,17'd23093,17'd23094,17'd22918,17'd22407,17'd23095,17'd22564,17'd22752,17'd22391,17'd22928,17'd22567,17'd22392,17'd22392,17'd22392,17'd23096,17'd23096,17'd23097,17'd23097,17'd22220,17'd23098,17'd22225,17'd22069,17'd23099,17'd23100,17'd23101,17'd22224,17'd23102,17'd23103,17'd23104,17'd23105,17'd23106,17'd23107,17'd23108,17'd23109,17'd23110,17'd22759,17'd7989,17'd22588,17'd23111,17'd23112,17'd23113,17'd23114,17'd23115,17'd23116,17'd15094,17'd14971,17'd18742,17'd18742,17'd16121,17'd17065,17'd15724,17'd17282,17'd17283,17'd20542,17'd20542,17'd20542,17'd17903,17'd17065,17'd19221,17'd16121,17'd18260,17'd20849,17'd23117,17'd23118,17'd19851,17'd21777,17'd23119,17'd23120,17'd16490,17'd14731,17'd18029,17'd23121,17'd23122,17'd23123,17'd23124,17'd23125,17'd23126,17'd23127,17'd23128,17'd2738,17'd430,17'd187,17'd9662,17'd23129,17'd3582,17'd3729,17'd2105,17'd19104,17'd4232,17'd3573,17'd4870,17'd3397,17'd7513,17'd8795,17'd8796,17'd11189,17'd23130,17'd23131,17'd10248,17'd8796,17'd7513,17'd23132,17'd23133,17'd23134,17'd23135,17'd23136,17'd9405,17'd8019,17'd8491,17'd8795,17'd14062,17'd8796,17'd7858,17'd7686,17'd7685,17'd4872,17'd9116,17'd7349,17'd7861,17'd7522,17'd22961,17'd23137,17'd22443,17'd23138,17'd2415,17'd23139,17'd648,17'd20720,17'd15492,17'd17185
},
'{
17'd8971,17'd3430,17'd466,17'd466,17'd1416,17'd3905,17'd11,17'd21,17'd4,17'd3594,17'd5793,17'd8040,17'd8040,17'd8040,17'd5205,17'd5205,17'd8040,17'd5205,17'd3753,17'd5,17'd24,17'd24,17'd23,17'd4,17'd24,17'd24,17'd3594,17'd3594,17'd5,17'd5,17'd5,17'd5,17'd23,17'd25,17'd286,17'd28,17'd3755,17'd3431,17'd2263,17'd2121,17'd22966,17'd989,17'd825,17'd666,17'd482,17'd14603,17'd22968,17'd14604,17'd23140,17'd23141,17'd23142,17'd3607,17'd23143,17'd23144,17'd22973,17'd23145,17'd12663,17'd23146,17'd23147,17'd13701,17'd16647,17'd23148,17'd23149,17'd18527,17'd22626,17'd23150,17'd23151,17'd23152,17'd23153,17'd16287,17'd12361,17'd12530,17'd14890,17'd14890,17'd21184,17'd13092,17'd22802,17'd19127,17'd19127,17'd12527,17'd11626,17'd23154,17'd17096,17'd14621,17'd14764,17'd14621,17'd12218,17'd12362,17'd12531,17'd20886,17'd23155,17'd21649,17'd21650,17'd19256,17'd17320,17'd16411,17'd14765,17'd15260,17'd15768,17'd15523,17'd22981,17'd18297,17'd19384,17'd23156,17'd20426,17'd22633,17'd22634,17'd12533,17'd9701,17'd6931,17'd7412,17'd7413,17'd9004,17'd9004,17'd7414,17'd7414,17'd7749,17'd9570,17'd9844,17'd9844,17'd10949,17'd11918,17'd13610,17'd21044,17'd20891,17'd23157,17'd19522,17'd17107,17'd16183,17'd14784,17'd12827,17'd23158,17'd23159,17'd23160,17'd23161,17'd12570,17'd11946,17'd22988,17'd21814,17'd22293,17'd12559,17'd12843,17'd12089,17'd12401,17'd23162,17'd19776,17'd18913,17'd23163,17'd23164,17'd10475,17'd23165,17'd8721,17'd8874,17'd16549,17'd10166,17'd10474,17'd16320,17'd11399,17'd11525,17'd23166,17'd23167,17'd11959,17'd12578,17'd12256,17'd13643,17'd13643,17'd14525,17'd12416,17'd18564,17'd23168,17'd21505,17'd21361,17'd23169,17'd21985,17'd18327,17'd23167,17'd21363,17'd23170,17'd22819,17'd22819,17'd19408,17'd18917,17'd17604,17'd19922,17'd12262,17'd11963,17'd11960,17'd14130,17'd11959,17'd15053,17'd12996,17'd11963,17'd12858,17'd12996,17'd13135,17'd13646,17'd23171,17'd23172,17'd12584,17'd16912,17'd9344,17'd17123,17'd8726,17'd8572,17'd8576,17'd9196,17'd23173,17'd23174,17'd23175,17'd16448,17'd12727,17'd23176,17'd23177,17'd15441,17'd23178,17'd16076,17'd21058,17'd23179,17'd23180,17'd16080,17'd23181,17'd8267,17'd23182,17'd23183,17'd23184,17'd23185,17'd23185,17'd23186,17'd23187,17'd23188,17'd19164,17'd23189,17'd23190,17'd23191,17'd23192,17'd23193,17'd17136,17'd17615,17'd14274,17'd13533,17'd23015,17'd13899,17'd23194,17'd541,17'd1481,17'd133,17'd131,17'd131,17'd11541,17'd11541,17'd131,17'd132,17'd134,17'd20466,17'd20624,17'd20629,17'd23195,17'd23196,17'd23197,17'd23198,17'd23199,17'd23200,17'd23201,17'd23202,17'd23027,17'd23203,17'd23204,17'd23205,17'd23206,17'd23207,17'd23208,17'd23208,17'd23209,17'd23210,17'd23211,17'd23212,17'd23213,17'd23214,17'd23215,17'd23216,17'd23217,17'd23218,17'd23218,17'd22329,17'd22330,17'd22856,17'd22506,17'd22333,17'd23219,17'd22333,17'd23220,17'd23221,17'd21845,17'd21845,17'd23222,17'd22864,17'd22514,17'd23223,17'd23224,17'd23225,17'd23226,17'd23227,17'd23228,17'd23229,17'd23230,17'd23231,17'd22185,17'd23232,17'd23233,17'd23234,17'd23060,17'd23235,17'd23236,17'd23237,17'd23238,17'd23239,17'd23066,17'd21874,17'd23240,17'd22535,17'd23241,17'd19184,17'd23242,17'd23243,17'd23244,17'd23245,17'd23246,17'd23247,17'd23248,17'd23249,17'd23250,17'd23251,17'd23252,17'd23253,17'd23254,17'd23255,17'd23256,17'd23257,17'd23258,17'd20093,17'd23259,17'd20830,17'd23260,17'd23261,17'd23262,17'd23263,17'd20497,17'd22732,17'd22733,17'd23264,17'd21298,17'd23265,17'd23266,17'd22407,17'd23095,17'd23095,17'd22752,17'd23267,17'd23268,17'd22928,17'd22567,17'd22567,17'd22392,17'd23096,17'd23096,17'd23096,17'd23269,17'd23270,17'd22223,17'd22067,17'd23271,17'd23272,17'd21908,17'd23272,17'd23271,17'd22067,17'd23273,17'd23274,17'd23275,17'd23276,17'd23107,17'd23107,17'd23277,17'd23278,17'd23279,17'd22935,17'd7824,17'd23280,17'd23281,17'd23282,17'd23283,17'd23284,17'd23285,17'd23286,17'd14046,17'd13406,17'd15340,17'd17904,17'd15988,17'd16247,17'd15605,17'd15724,17'd17903,17'd17903,17'd18373,17'd18373,17'd17903,17'd17065,17'd15336,17'd15337,17'd15988,17'd23287,17'd15479,17'd18622,17'd23288,17'd23289,17'd23290,17'd23120,17'd23291,17'd14731,17'd23292,17'd18860,17'd23293,17'd23294,17'd23295,17'd23296,17'd23297,17'd23298,17'd23299,17'd23300,17'd430,17'd187,17'd23301,17'd10389,17'd3411,17'd3728,17'd2105,17'd3718,17'd3397,17'd3396,17'd3876,17'd3573,17'd5184,17'd23302,17'd14436,17'd8168,17'd23303,17'd23304,17'd8794,17'd8954,17'd23305,17'd23306,17'd23307,17'd23308,17'd23309,17'd23136,17'd8795,17'd8019,17'd8491,17'd8491,17'd14062,17'd14180,17'd7856,17'd7685,17'd7684,17'd7343,17'd9116,17'd4719,17'd4567,17'd7522,17'd5640,17'd23310,17'd7872,17'd23311,17'd23312,17'd23313,17'd648,17'd648,17'd15626,17'd15492
},
'{
17'd2595,17'd2595,17'd466,17'd466,17'd1416,17'd3905,17'd11,17'd23,17'd5,17'd3753,17'd5793,17'd8040,17'd8040,17'd8040,17'd5205,17'd5205,17'd5205,17'd3753,17'd3753,17'd5,17'd24,17'd23,17'd23,17'd23,17'd24,17'd24,17'd5,17'd5,17'd5,17'd5,17'd5,17'd5,17'd1691,17'd467,17'd286,17'd29,17'd3255,17'd2942,17'd2263,17'd22615,17'd22966,17'd21949,17'd19609,17'd666,17'd482,17'd14603,17'd22968,17'd14604,17'd2128,17'd22790,17'd23314,17'd23315,17'd23316,17'd23317,17'd23318,17'd23145,17'd23319,17'd23320,17'd23147,17'd23321,17'd19374,17'd23322,17'd23149,17'd18527,17'd22626,17'd23323,17'd23151,17'd22117,17'd23324,17'd16027,17'd12361,17'd12530,17'd14890,17'd14890,17'd13209,17'd13092,17'd14469,17'd14469,17'd19127,17'd12527,17'd12813,17'd23325,17'd13211,17'd14621,17'd12218,17'd12218,17'd12218,17'd12530,17'd11913,17'd12681,17'd17941,17'd21964,17'd21650,17'd17320,17'd17690,17'd16411,17'd16032,17'd15009,17'd15645,17'd22118,17'd16170,17'd18658,17'd20735,17'd20426,17'd11088,17'd22633,17'd9573,17'd9701,17'd7086,17'd7413,17'd7414,17'd8218,17'd23326,17'd9004,17'd8218,17'd7579,17'd7748,17'd8065,17'd9844,17'd10947,17'd23327,17'd10289,17'd21657,17'd21657,17'd23328,17'd20161,17'd17458,17'd23329,17'd14907,17'd19908,17'd23330,17'd23331,17'd10712,17'd16429,17'd23332,17'd18800,17'd23333,17'd21049,17'd20305,17'd13506,17'd23334,17'd23334,17'd13506,17'd20305,17'd23335,17'd11658,17'd19153,17'd15678,17'd23336,17'd10328,17'd9339,17'd8720,17'd9345,17'd11277,17'd11670,17'd11669,17'd10854,17'd11131,17'd21206,17'd23337,17'd19920,17'd15184,17'd12578,17'd12576,17'd18684,17'd13643,17'd22297,17'd21504,17'd12255,17'd23168,17'd22992,17'd18681,17'd21985,17'd18327,17'd16442,17'd21361,17'd22818,17'd22819,17'd23168,17'd21671,17'd15053,17'd12422,17'd12115,17'd17968,17'd11963,17'd13135,17'd11959,17'd11959,17'd18198,17'd12996,17'd11963,17'd11963,17'd16204,17'd16204,17'd11806,17'd11667,17'd23338,17'd12720,17'd23339,17'd23340,17'd15569,17'd9044,17'd11403,17'd23341,17'd23342,17'd8578,17'd23343,17'd8420,17'd15692,17'd14531,17'd10029,17'd16073,17'd17238,17'd23344,17'd23345,17'd13653,17'd10610,17'd23346,17'd23347,17'd15308,17'd23348,17'd19927,17'd23349,17'd23349,17'd23350,17'd23351,17'd20324,17'd23352,17'd23353,17'd23354,17'd23185,17'd23187,17'd23355,17'd17613,17'd14537,17'd23356,17'd15819,17'd23357,17'd23358,17'd23359,17'd15958,17'd17616,17'd22310,17'd16219,17'd13900,17'd15823,17'd132,17'd134,17'd131,17'd131,17'd132,17'd132,17'd356,17'd15823,17'd23360,17'd22844,17'd23196,17'd23361,17'd23362,17'd23363,17'd23364,17'd23365,17'd23366,17'd23367,17'd23368,17'd23369,17'd23370,17'd23371,17'd23372,17'd23373,17'd23374,17'd23375,17'd23376,17'd23377,17'd23378,17'd23379,17'd23380,17'd23381,17'd23382,17'd23383,17'd23384,17'd23385,17'd23386,17'd23387,17'd23388,17'd23215,17'd23389,17'd23218,17'd23390,17'd22326,17'd23391,17'd23392,17'd23393,17'd23394,17'd23395,17'd23396,17'd23397,17'd23398,17'd23399,17'd23400,17'd23401,17'd23402,17'd23403,17'd23404,17'd23405,17'd23233,17'd23406,17'd23407,17'd23408,17'd23409,17'd23410,17'd23411,17'd23412,17'd23413,17'd23414,17'd23415,17'd23416,17'd22188,17'd23417,17'd23418,17'd23419,17'd20205,17'd23420,17'd23421,17'd23422,17'd23423,17'd23424,17'd23425,17'd22200,17'd22046,17'd23426,17'd23427,17'd23428,17'd23429,17'd23430,17'd23431,17'd23432,17'd23433,17'd20666,17'd20223,17'd23434,17'd23435,17'd23436,17'd23437,17'd23438,17'd21756,17'd23439,17'd23440,17'd23441,17'd23442,17'd23443,17'd23265,17'd23444,17'd22563,17'd22390,17'd22390,17'd22565,17'd23268,17'd22392,17'd23097,17'd23097,17'd23097,17'd22222,17'd22222,17'd22222,17'd23445,17'd23445,17'd23445,17'd23446,17'd23447,17'd23448,17'd23449,17'd21904,17'd21904,17'd22064,17'd22221,17'd23450,17'd23451,17'd23452,17'd23453,17'd23454,17'd23455,17'd23456,17'd23457,17'd23279,17'd22935,17'd9503,17'd23458,17'd23459,17'd23460,17'd23461,17'd23462,17'd22763,17'd23285,17'd14045,17'd12306,17'd14971,17'd15340,17'd19590,17'd16247,17'd15093,17'd15605,17'd17779,17'd17903,17'd23463,17'd18373,17'd17779,17'd17065,17'd16119,17'd16121,17'd18260,17'd23464,17'd23465,17'd21775,17'd19989,17'd23466,17'd23467,17'd21617,17'd23468,17'd14731,17'd23292,17'd18860,17'd19595,17'd23469,17'd23470,17'd23471,17'd23472,17'd23473,17'd23474,17'd23475,17'd933,17'd267,17'd8485,17'd20564,17'd20401,17'd12638,17'd1954,17'd3404,17'd3402,17'd4870,17'd3226,17'd6240,17'd23476,17'd7854,17'd23477,17'd8017,17'd21946,17'd14590,17'd11189,17'd14590,17'd23478,17'd23479,17'd23480,17'd23481,17'd23482,17'd23483,17'd8491,17'd8491,17'd8170,17'd8491,17'd14062,17'd8796,17'd7858,17'd7029,17'd7685,17'd4872,17'd9116,17'd7519,17'd7861,17'd4071,17'd23484,17'd23137,17'd23485,17'd23486,17'd23487,17'd23488,17'd23489,17'd648,17'd180,17'd15626
},
'{
17'd2595,17'd2595,17'd466,17'd466,17'd17,17'd18,17'd10,17'd4,17'd6,17'd3753,17'd5793,17'd8040,17'd8040,17'd8040,17'd5205,17'd3753,17'd3753,17'd3753,17'd6,17'd5,17'd23,17'd22,17'd22,17'd23,17'd24,17'd24,17'd5,17'd5,17'd5,17'd5,17'd5,17'd4,17'd1832,17'd285,17'd28,17'd289,17'd3254,17'd2943,17'd2785,17'd22615,17'd23490,17'd989,17'd825,17'd666,17'd482,17'd14603,17'd668,17'd2614,17'd23491,17'd22970,17'd2799,17'd23492,17'd23493,17'd23494,17'd23318,17'd23495,17'd23496,17'd13312,17'd22796,17'd19619,17'd23497,17'd23498,17'd18649,17'd17678,17'd23499,17'd23500,17'd23152,17'd23153,17'd16163,17'd15764,17'd12218,17'd12530,17'd14890,17'd12955,17'd13209,17'd13092,17'd14469,17'd14469,17'd22802,17'd12527,17'd12813,17'd17096,17'd14621,17'd14621,17'd12218,17'd13094,17'd12218,17'd11913,17'd12531,17'd17941,17'd17205,17'd15765,17'd19256,17'd16033,17'd16411,17'd16987,17'd16032,17'd15261,17'd21965,17'd22118,17'd23501,17'd15898,17'd15765,17'd20426,17'd11088,17'd11088,17'd9573,17'd9701,17'd7086,17'd7413,17'd8218,17'd23326,17'd9004,17'd9004,17'd7414,17'd7579,17'd8065,17'd9570,17'd10566,17'd10949,17'd11919,17'd10433,17'd23328,17'd23328,17'd23502,17'd19522,17'd23503,17'd15026,17'd23504,17'd23505,17'd23506,17'd19148,17'd23507,17'd12241,17'd12989,17'd13997,17'd21049,17'd23508,17'd19914,17'd16901,17'd20601,17'd15676,17'd13131,17'd23509,17'd11795,17'd12852,17'd12249,17'd16906,17'd23510,17'd18441,17'd9191,17'd9346,17'd16549,17'd11135,17'd15176,17'd11399,17'd10854,17'd11131,17'd10990,17'd17125,17'd15184,17'd12253,17'd12256,17'd12257,17'd13760,17'd12418,17'd19534,17'd23511,17'd23512,17'd22819,17'd16325,17'd18444,17'd22817,17'd23513,17'd22992,17'd23170,17'd23514,17'd23515,17'd21671,17'd18198,17'd16204,17'd12115,17'd12115,17'd12262,17'd11806,17'd13883,17'd11959,17'd18198,17'd15053,17'd16204,17'd13362,17'd19157,17'd12115,17'd11807,17'd11667,17'd13000,17'd21986,17'd19532,17'd23516,17'd10743,17'd9345,17'd16681,17'd9046,17'd23517,17'd8574,17'd8732,17'd12426,17'd16691,17'd15440,17'd23518,17'd13768,17'd8734,17'd23519,17'd23520,17'd23521,17'd7619,17'd23522,17'd14683,17'd23523,17'd8429,17'd8588,17'd23524,17'd23525,17'd17487,17'd15309,17'd14395,17'd23526,17'd15577,17'd13009,17'd23527,17'd23528,17'd23529,17'd23530,17'd13010,17'd14820,17'd10614,17'd12125,17'd11819,17'd11681,17'd23358,17'd23531,17'd23532,17'd23533,17'd23534,17'd23535,17'd23536,17'd131,17'd132,17'd132,17'd132,17'd132,17'd1197,17'd133,17'd23537,17'd23538,17'd23539,17'd23540,17'd23362,17'd23541,17'd23542,17'd23543,17'd23544,17'd23205,17'd23545,17'd23370,17'd23546,17'd23547,17'd23548,17'd23549,17'd23550,17'd23551,17'd23552,17'd23553,17'd23554,17'd23555,17'd23556,17'd23557,17'd23558,17'd23559,17'd23560,17'd23561,17'd23562,17'd23563,17'd23564,17'd23565,17'd23566,17'd23387,17'd23567,17'd23568,17'd23569,17'd23570,17'd23571,17'd23572,17'd23573,17'd23574,17'd23575,17'd23576,17'd23577,17'd23578,17'd23579,17'd23580,17'd23581,17'd23582,17'd23583,17'd23584,17'd23585,17'd23586,17'd23587,17'd23588,17'd23589,17'd23410,17'd23590,17'd23235,17'd23591,17'd23592,17'd23593,17'd23594,17'd22888,17'd23595,17'd23417,17'd22188,17'd23596,17'd23597,17'd23598,17'd23599,17'd23600,17'd23601,17'd23602,17'd23603,17'd23604,17'd23605,17'd22901,17'd23606,17'd23607,17'd23608,17'd23608,17'd23429,17'd23609,17'd23080,17'd23610,17'd23611,17'd20831,17'd21598,17'd23612,17'd21914,17'd21756,17'd21602,17'd21603,17'd21448,17'd21297,17'd21762,17'd23613,17'd23614,17'd23615,17'd23616,17'd23617,17'd23618,17'd23619,17'd23620,17'd23621,17'd23620,17'd23620,17'd23622,17'd23623,17'd23624,17'd23624,17'd23624,17'd23623,17'd23625,17'd23626,17'd23446,17'd23448,17'd22067,17'd22067,17'd22221,17'd22222,17'd23106,17'd23275,17'd23452,17'd23455,17'd23454,17'd23455,17'd23627,17'd23457,17'd23279,17'd23628,17'd8608,17'd7824,17'd8144,17'd23629,17'd23630,17'd23631,17'd23632,17'd23633,17'd14045,17'd12904,17'd13558,17'd17655,17'd16955,17'd16121,17'd14570,17'd15605,17'd17779,17'd17779,17'd23463,17'd18373,17'd17903,17'd17065,17'd15475,17'd15337,17'd15988,17'd20384,17'd23634,17'd16127,17'd23118,17'd20699,17'd23635,17'd22946,17'd23636,17'd22948,17'd15100,17'd21937,17'd19353,17'd23637,17'd23638,17'd23639,17'd23640,17'd23641,17'd2553,17'd23642,17'd23643,17'd2588,17'd3415,17'd23644,17'd23645,17'd3235,17'd18986,17'd2406,17'd4870,17'd5633,17'd2912,17'd5633,17'd23646,17'd23647,17'd23648,17'd22608,17'd7853,17'd21946,17'd8168,17'd23649,17'd23650,17'd23651,17'd23652,17'd23653,17'd23134,17'd23654,17'd23302,17'd8491,17'd8491,17'd8491,17'd14062,17'd14062,17'd8171,17'd7685,17'd7684,17'd4872,17'd9116,17'd4718,17'd4567,17'd6875,17'd5640,17'd23655,17'd7870,17'd23656,17'd23657,17'd23313,17'd23489,17'd648,17'd180,17'd15492
},
'{
17'd2595,17'd2595,17'd466,17'd466,17'd13,17'd3,17'd808,17'd4,17'd6,17'd3753,17'd5793,17'd8040,17'd8040,17'd8040,17'd3753,17'd3753,17'd3753,17'd3753,17'd5,17'd24,17'd22,17'd22,17'd22,17'd22,17'd24,17'd24,17'd5,17'd5,17'd5,17'd5,17'd4,17'd23,17'd1832,17'd285,17'd6744,17'd3595,17'd3254,17'd2943,17'd2785,17'd23658,17'd23490,17'd1134,17'd991,17'd667,17'd14450,17'd483,17'd832,17'd23659,17'd23660,17'd23661,17'd23662,17'd6448,17'd23663,17'd23664,17'd22793,17'd23665,17'd21643,17'd13195,17'd20580,17'd13959,17'd23666,17'd23667,17'd14201,17'd15755,17'd23668,17'd23669,17'd22117,17'd23153,17'd16163,17'd13969,17'd12218,17'd12530,17'd12955,17'd12679,17'd14469,17'd14469,17'd14469,17'd14469,17'd22802,17'd12527,17'd12813,17'd13211,17'd14764,17'd14621,17'd13094,17'd13094,17'd12680,17'd11913,17'd12532,17'd19753,17'd16986,17'd19384,17'd17694,17'd16768,17'd17811,17'd15260,17'd16032,17'd15770,17'd23670,17'd23670,17'd15766,17'd15766,17'd10429,17'd13471,17'd9574,17'd9158,17'd8687,17'd7086,17'd8366,17'd9004,17'd9004,17'd23326,17'd9004,17'd8366,17'd7749,17'd8685,17'd10119,17'd20435,17'd10698,17'd11092,17'd10289,17'd23671,17'd10290,17'd23502,17'd20033,17'd22122,17'd21351,17'd23672,17'd10705,17'd23673,17'd23674,17'd18673,17'd13237,17'd18800,17'd12097,17'd23675,17'd22128,17'd23676,17'd17833,17'd23677,17'd15172,17'd12243,17'd18189,17'd13997,17'd17007,17'd16062,17'd23678,17'd10324,17'd20174,17'd14804,17'd23679,17'd11809,17'd14928,17'd12863,17'd21206,17'd11668,17'd11275,17'd11130,17'd10736,17'd18679,17'd23680,17'd15434,17'd12256,17'd12257,17'd12856,17'd12418,17'd19534,17'd23681,17'd23515,17'd21505,17'd19158,17'd13645,17'd18444,17'd16325,17'd22818,17'd23515,17'd23682,17'd23515,17'd19408,17'd15053,17'd12262,17'd18560,17'd15810,17'd13362,17'd11960,17'd11959,17'd19408,17'd17722,17'd18917,17'd12422,17'd12262,17'd15810,17'd11964,17'd13253,17'd11666,17'd15182,17'd16320,17'd23683,17'd21056,17'd9478,17'd17840,17'd16910,17'd23684,17'd12424,17'd8574,17'd8414,17'd23685,17'd8252,17'd7952,17'd23686,17'd7949,17'd11278,17'd11278,17'd23687,17'd23688,17'd23689,17'd14141,17'd23690,17'd7626,17'd19038,17'd19289,17'd17973,17'd17973,17'd18690,17'd13379,17'd8265,17'd9625,17'd8741,17'd7305,17'd7965,17'd7965,17'd8267,17'd8117,17'd23691,17'd20460,17'd23692,17'd23693,17'd23694,17'd23695,17'd23696,17'd11005,17'd18210,17'd23697,17'd23698,17'd23699,17'd23700,17'd1045,17'd130,17'd720,17'd130,17'd356,17'd1045,17'd22312,17'd23701,17'd23702,17'd23703,17'd23704,17'd23705,17'd23706,17'd23707,17'd23708,17'd23709,17'd23710,17'd23711,17'd23712,17'd23713,17'd23714,17'd23715,17'd23716,17'd23717,17'd23718,17'd23719,17'd23720,17'd23719,17'd23721,17'd23722,17'd23723,17'd23724,17'd23725,17'd23726,17'd23727,17'd23728,17'd23729,17'd23730,17'd23731,17'd23732,17'd23733,17'd23734,17'd23735,17'd23736,17'd23737,17'd23738,17'd23739,17'd23740,17'd23741,17'd23742,17'd23743,17'd23744,17'd23745,17'd23746,17'd23747,17'd23748,17'd23749,17'd23750,17'd23751,17'd23752,17'd22702,17'd23753,17'd23754,17'd23588,17'd23755,17'd23756,17'd23757,17'd23758,17'd23759,17'd23760,17'd23761,17'd23594,17'd23762,17'd23763,17'd23764,17'd23239,17'd22889,17'd23765,17'd23598,17'd23766,17'd23767,17'd23768,17'd23245,17'd23769,17'd23770,17'd23771,17'd23772,17'd23773,17'd23774,17'd23775,17'd23428,17'd23776,17'd23777,17'd20814,17'd23778,17'd20985,17'd23779,17'd23780,17'd23781,17'd21757,17'd23782,17'd23783,17'd23784,17'd21760,17'd23785,17'd23786,17'd22408,17'd22409,17'd23787,17'd23788,17'd23789,17'd22755,17'd23790,17'd22931,17'd23791,17'd23791,17'd23791,17'd23791,17'd23791,17'd23792,17'd23792,17'd23106,17'd23793,17'd23794,17'd23625,17'd23446,17'd22066,17'd22066,17'd22066,17'd23795,17'd23796,17'd23107,17'd23797,17'd23627,17'd23457,17'd23627,17'd23457,17'd23798,17'd8911,17'd8289,17'd7659,17'd7326,17'd23799,17'd6382,17'd5914,17'd23800,17'd23801,17'd23802,17'd13165,17'd11314,17'd13407,17'd13925,17'd22420,17'd18742,17'd16121,17'd15093,17'd17779,17'd17779,17'd23463,17'd18373,17'd17903,17'd17779,17'd15475,17'd17533,17'd19590,17'd20250,17'd23803,17'd20546,17'd19850,17'd23804,17'd23805,17'd20549,17'd23806,17'd14056,17'd14307,17'd18379,17'd21937,17'd23807,17'd23808,17'd23809,17'd23810,17'd23811,17'd23812,17'd23813,17'd23814,17'd1242,17'd9790,17'd23815,17'd19494,17'd3410,17'd19495,17'd1816,17'd3395,17'd3226,17'd2748,17'd2910,17'd5638,17'd23135,17'd23816,17'd23476,17'd23816,17'd7194,17'd7513,17'd7194,17'd5782,17'd23817,17'd23818,17'd23819,17'd5781,17'd23820,17'd23483,17'd11444,17'd8491,17'd8491,17'd14062,17'd9534,17'd8020,17'd7686,17'd7346,17'd4872,17'd6576,17'd7519,17'd7861,17'd3576,17'd23484,17'd23821,17'd23485,17'd23822,17'd23823,17'd23313,17'd23489,17'd23489,17'd15626,17'd17422
},
'{
17'd2595,17'd2595,17'd2595,17'd466,17'd13,17'd806,17'd25,17'd4,17'd6,17'd3753,17'd5793,17'd8040,17'd8040,17'd8040,17'd3753,17'd3753,17'd3753,17'd3753,17'd5,17'd24,17'd22,17'd5518,17'd22,17'd22,17'd24,17'd24,17'd5,17'd5,17'd5,17'd5,17'd23,17'd23,17'd285,17'd286,17'd4431,17'd3595,17'd2940,17'd3253,17'd23824,17'd22615,17'd22966,17'd990,17'd824,17'd667,17'd14450,17'd831,17'd996,17'd23825,17'd23826,17'd23827,17'd4101,17'd23828,17'd23663,17'd6914,17'd22621,17'd23829,17'd21802,17'd20141,17'd23830,17'd23831,17'd23666,17'd23832,17'd18049,17'd23833,17'd23834,17'd23835,17'd23836,17'd16287,17'd12361,17'd13969,17'd12530,17'd12814,17'd12528,17'd12527,17'd14469,17'd14469,17'd14469,17'd14469,17'd22802,17'd12527,17'd13093,17'd14621,17'd14764,17'd14621,17'd13094,17'd12218,17'd12680,17'd10815,17'd17204,17'd16766,17'd16164,17'd15899,17'd16290,17'd14892,17'd15520,17'd15260,17'd16032,17'd15770,17'd23837,17'd23837,17'd16880,17'd16880,17'd10429,17'd9574,17'd11232,17'd9158,17'd8536,17'd7413,17'd9004,17'd23326,17'd23326,17'd9004,17'd8366,17'd7749,17'd10287,17'd21489,17'd20435,17'd10698,17'd11092,17'd10289,17'd23671,17'd23838,17'd23502,17'd20298,17'd23839,17'd23840,17'd13858,17'd23841,17'd23842,17'd10000,17'd23843,17'd14119,17'd11937,17'd12246,17'd23844,17'd23845,17'd23846,17'd21051,17'd23847,17'd23848,17'd12710,17'd19639,17'd20305,17'd18912,17'd23849,17'd23850,17'd23851,17'd23852,17'd10744,17'd23853,17'd9480,17'd14928,17'd11528,17'd15176,17'd21206,17'd11668,17'd11275,17'd10989,17'd16797,17'd23854,17'd12578,17'd15434,17'd12575,17'd12575,17'd12575,17'd15434,17'd23855,17'd23512,17'd23170,17'd21361,17'd16326,17'd13516,17'd19158,17'd22992,17'd23515,17'd23682,17'd23856,17'd23168,17'd11959,17'd16204,17'd18560,17'd18682,17'd12262,17'd12996,17'd11960,17'd11959,17'd18198,17'd18197,17'd12422,17'd12262,17'd12262,17'd14262,17'd11807,17'd13137,17'd15432,17'd13001,17'd23683,17'd18323,17'd23857,17'd12117,17'd23858,17'd23859,17'd23860,17'd23861,17'd8572,17'd12725,17'd13004,17'd8102,17'd23862,17'd23863,17'd23864,17'd23865,17'd23866,17'd16690,17'd10180,17'd23867,17'd23868,17'd10030,17'd16449,17'd23869,17'd19038,17'd23870,17'd23870,17'd18091,17'd23871,17'd23872,17'd8740,17'd8116,17'd23873,17'd23874,17'd8741,17'd8266,17'd23875,17'd13530,17'd16452,17'd23876,17'd23877,17'd23878,17'd23879,17'd23880,17'd17736,17'd18576,17'd23881,17'd23882,17'd23883,17'd23884,17'd23885,17'd134,17'd128,17'd136,17'd1481,17'd17363,17'd23886,17'd23887,17'd23888,17'd23889,17'd23890,17'd23891,17'd23892,17'd23893,17'd23894,17'd23895,17'd23896,17'd23897,17'd23898,17'd23899,17'd23900,17'd23901,17'd23902,17'd23903,17'd23904,17'd23905,17'd23905,17'd23906,17'd23907,17'd23718,17'd23908,17'd23909,17'd23910,17'd23911,17'd23912,17'd23913,17'd23914,17'd23915,17'd23916,17'd23917,17'd23732,17'd23918,17'd23919,17'd23920,17'd23921,17'd23922,17'd23384,17'd23923,17'd23924,17'd23925,17'd23926,17'd23927,17'd23928,17'd23929,17'd23930,17'd23931,17'd23932,17'd23933,17'd23934,17'd23935,17'd23936,17'd22884,17'd23937,17'd23938,17'd23939,17'd23940,17'd23941,17'd23412,17'd23942,17'd23943,17'd23944,17'd23945,17'd23415,17'd23946,17'd23947,17'd23948,17'd22888,17'd23949,17'd23950,17'd23951,17'd23952,17'd23953,17'd23954,17'd23074,17'd23955,17'd23956,17'd23957,17'd23958,17'd23959,17'd22902,17'd22374,17'd23960,17'd22550,17'd20967,17'd23961,17'd19695,17'd20102,17'd21599,17'd23962,17'd21757,17'd21915,17'd23963,17'd23964,17'd23965,17'd23966,17'd23967,17'd22239,17'd22409,17'd22410,17'd23968,17'd23968,17'd23969,17'd23969,17'd23970,17'd23970,17'd23971,17'd23791,17'd23792,17'd23792,17'd23792,17'd23792,17'd23792,17'd23796,17'd23793,17'd23972,17'd23625,17'd23625,17'd23625,17'd23973,17'd23973,17'd23108,17'd23278,17'd23798,17'd6840,17'd23974,17'd6840,17'd6840,17'd8911,17'd8911,17'd8289,17'd7659,17'd7163,17'd23975,17'd8144,17'd6382,17'd23461,17'd23976,17'd23977,17'd23978,17'd11314,17'd13166,17'd13406,17'd15476,17'd18022,17'd15988,17'd14570,17'd17065,17'd17779,17'd23463,17'd23463,17'd17903,17'd17779,17'd15603,17'd15336,17'd16121,17'd19479,17'd23979,17'd23980,17'd19224,17'd23981,17'd23982,17'd11582,17'd23983,17'd17908,17'd15100,17'd18379,17'd18029,17'd19721,17'd23984,17'd2880,17'd23985,17'd23986,17'd23987,17'd23988,17'd1665,17'd210,17'd19493,17'd2577,17'd8165,17'd4061,17'd4231,17'd2914,17'd2912,17'd2912,17'd2744,17'd2746,17'd23989,17'd23482,17'd23990,17'd23646,17'd23305,17'd23816,17'd23305,17'd23991,17'd23481,17'd23992,17'd23993,17'd23994,17'd23995,17'd23996,17'd23483,17'd11444,17'd8491,17'd8491,17'd14062,17'd13934,17'd8019,17'd7685,17'd7516,17'd4717,17'd6576,17'd7193,17'd7518,17'd3405,17'd23484,17'd23997,17'd7870,17'd23998,17'd23999,17'd23313,17'd24000,17'd23489,17'd15626,17'd17185
},
'{
17'd4247,17'd4247,17'd2595,17'd466,17'd13,17'd806,17'd25,17'd4,17'd6,17'd3753,17'd5793,17'd5793,17'd8040,17'd5793,17'd5793,17'd5793,17'd3753,17'd3594,17'd5,17'd24,17'd22,17'd5518,17'd5518,17'd22,17'd24,17'd24,17'd5,17'd5,17'd4,17'd23,17'd23,17'd22,17'd285,17'd27,17'd4431,17'd3433,17'd2940,17'd3253,17'd23824,17'd22615,17'd22966,17'd1281,17'd1137,17'd667,17'd16637,17'd994,17'd1710,17'd2952,17'd24001,17'd23315,17'd24002,17'd6607,17'd24003,17'd6914,17'd24004,17'd24005,17'd24006,17'd23147,17'd24007,17'd24008,17'd16399,17'd24009,17'd16153,17'd24010,17'd24011,17'd22117,17'd21963,17'd16287,17'd12362,17'd11764,17'd12530,17'd12065,17'd12679,17'd12527,17'd12357,17'd14469,17'd14469,17'd14469,17'd15516,17'd12527,17'd12955,17'd14621,17'd12218,17'd13094,17'd13094,17'd12218,17'd11764,17'd11629,17'd17941,17'd19754,17'd16164,17'd16169,17'd24012,17'd15008,17'd24013,17'd15642,17'd16032,17'd15645,17'd23501,17'd16028,17'd16880,17'd16880,17'd10429,17'd9574,17'd11232,17'd9573,17'd7086,17'd7413,17'd9004,17'd24014,17'd23326,17'd8366,17'd7414,17'd7749,17'd21489,17'd24015,17'd20436,17'd10567,17'd10122,17'd10289,17'd23502,17'd24016,17'd24017,17'd17822,17'd19766,17'd20039,17'd10821,17'd20894,17'd24018,17'd24019,17'd24020,17'd12239,17'd12570,17'd11946,17'd24021,17'd24022,17'd24023,17'd24024,17'd24025,17'd24026,17'd21355,17'd21665,17'd12407,17'd18438,17'd24027,17'd16791,17'd24028,17'd18332,17'd9191,17'd9344,17'd15566,17'd11276,17'd11527,17'd11132,17'd21206,17'd11668,17'd24029,17'd11807,17'd21204,17'd15686,17'd12256,17'd12859,17'd12418,17'd12418,17'd12253,17'd18564,17'd24030,17'd24031,17'd21363,17'd14258,17'd18444,17'd19158,17'd15053,17'd21671,17'd24032,17'd24033,17'd23856,17'd22819,17'd15053,17'd12262,17'd18682,17'd18560,17'd11963,17'd11806,17'd11960,17'd18198,17'd18917,17'd16204,17'd13516,17'd13516,17'd11964,17'd13762,17'd17125,17'd24034,17'd24035,17'd10326,17'd24036,17'd9471,17'd24037,17'd24038,17'd24039,17'd24040,17'd15684,17'd9195,17'd8572,17'd24041,17'd12867,17'd14384,17'd24042,17'd24043,17'd8887,17'd9048,17'd24044,17'd13649,17'd12727,17'd24045,17'd24046,17'd7462,17'd13529,17'd17020,17'd10863,17'd18922,17'd18922,17'd24047,17'd8587,17'd24048,17'd19650,17'd24049,17'd15445,17'd16337,17'd15697,17'd23000,17'd24050,17'd14535,17'd24051,17'd24052,17'd14272,17'd23876,17'd12732,17'd24053,17'd22832,17'd11682,17'd17736,17'd15068,17'd24054,17'd24055,17'd23700,17'd13777,17'd1481,17'd20762,17'd1480,17'd24056,17'd24057,17'd24058,17'd24059,17'd24060,17'd24061,17'd24062,17'd24063,17'd24064,17'd23897,17'd24065,17'd23898,17'd24066,17'd24067,17'd24068,17'd23903,17'd24069,17'd24070,17'd24071,17'd24071,17'd24072,17'd23906,17'd24073,17'd24074,17'd24075,17'd24076,17'd24077,17'd24078,17'd23724,17'd24079,17'd24080,17'd24081,17'd24082,17'd23381,17'd24083,17'd24084,17'd24085,17'd24086,17'd24087,17'd24088,17'd24089,17'd24090,17'd24091,17'd24092,17'd24093,17'd24094,17'd24095,17'd24096,17'd24097,17'd24098,17'd23931,17'd24099,17'd24100,17'd24101,17'd24102,17'd24103,17'd23412,17'd24104,17'd24105,17'd24106,17'd24107,17'd24108,17'd24109,17'd23412,17'd24110,17'd24111,17'd24112,17'd24113,17'd23946,17'd24114,17'd24114,17'd23763,17'd23417,17'd24115,17'd24116,17'd24117,17'd24118,17'd24119,17'd24120,17'd24121,17'd24122,17'd24123,17'd24124,17'd23959,17'd24125,17'd24126,17'd24127,17'd24128,17'd20812,17'd24129,17'd24130,17'd19696,17'd24131,17'd24132,17'd24133,17'd24134,17'd21758,17'd24135,17'd24136,17'd24137,17'd22734,17'd24138,17'd24139,17'd24140,17'd23968,17'd22411,17'd22584,17'd22584,17'd22757,17'd24141,17'd24141,17'd24142,17'd24142,17'd22932,17'd22933,17'd24143,17'd24143,17'd23108,17'd9637,17'd9637,17'd24144,17'd24145,17'd24146,17'd24147,17'd23797,17'd23457,17'd10881,17'd7656,17'd8142,17'd4678,17'd4679,17'd4679,17'd24148,17'd7006,17'd24149,17'd8143,17'd8143,17'd7326,17'd23799,17'd6212,17'd24150,17'd23800,17'd23801,17'd23802,17'd24151,17'd12904,17'd12306,17'd17655,17'd22420,17'd15725,17'd16121,17'd18498,17'd18619,17'd24152,17'd23463,17'd17903,17'd17779,17'd15724,17'd14570,17'd16121,17'd18260,17'd20251,17'd20545,17'd21615,17'd24153,17'd24154,17'd24155,17'd24156,17'd13567,17'd15100,17'd24157,17'd23292,17'd19486,17'd24158,17'd24159,17'd24160,17'd24161,17'd24162,17'd24163,17'd24164,17'd20008,17'd10073,17'd24165,17'd8316,17'd13057,17'd13421,17'd1252,17'd1387,17'd2748,17'd14738,17'd24166,17'd24167,17'd5781,17'd24168,17'd5638,17'd24168,17'd5779,17'd5779,17'd24169,17'd24170,17'd24171,17'd24172,17'd24173,17'd24174,17'd24175,17'd24176,17'd9945,17'd8170,17'd8170,17'd8491,17'd9405,17'd8020,17'd7029,17'd6871,17'd5635,17'd4872,17'd7193,17'd7689,17'd3405,17'd23484,17'd22611,17'd24177,17'd24178,17'd24179,17'd24180,17'd24000,17'd23489,17'd180,17'd15492
},
'{
17'd1688,17'd4247,17'd4247,17'd466,17'd13,17'd8814,17'd23,17'd5,17'd3753,17'd3753,17'd5793,17'd5793,17'd8040,17'd5793,17'd5793,17'd5793,17'd3753,17'd5,17'd5,17'd24,17'd5518,17'd5518,17'd5518,17'd5518,17'd24,17'd5,17'd5,17'd5,17'd4,17'd23,17'd22,17'd21,17'd286,17'd28,17'd4431,17'd3254,17'd2940,17'd2262,17'd1973,17'd22615,17'd22966,17'd1281,17'd1137,17'd1140,17'd1142,17'd1143,17'd997,17'd24181,17'd24182,17'd24183,17'd5391,17'd6607,17'd24003,17'd12042,17'd24184,17'd23496,17'd13195,17'd22796,17'd24185,17'd24186,17'd16399,17'd24187,17'd24188,17'd24189,17'd24190,17'd23836,17'd16287,17'd20885,17'd12680,17'd11627,17'd24191,17'd11626,17'd12679,17'd15516,17'd12357,17'd14469,17'd14469,17'd12357,17'd15516,17'd12813,17'd13211,17'd14621,17'd12218,17'd13094,17'd13094,17'd11913,17'd11361,17'd10427,17'd17205,17'd15765,17'd16028,17'd24192,17'd24193,17'd24194,17'd24195,17'd24013,17'd15769,17'd15645,17'd23501,17'd16028,17'd16880,17'd15766,17'd10429,17'd9574,17'd9574,17'd9573,17'd6931,17'd7580,17'd7086,17'd24196,17'd24197,17'd7414,17'd7414,17'd8685,17'd24198,17'd9845,17'd9989,17'd10567,17'd10122,17'd11484,17'd24016,17'd24199,17'd17948,17'd19766,17'd19767,17'd13735,17'd24200,17'd24201,17'd24202,17'd24203,17'd11109,17'd12989,17'd23335,17'd11946,17'd24204,17'd22468,17'd24205,17'd21050,17'd24206,17'd12096,17'd18800,17'd17960,17'd19275,17'd12852,17'd23850,17'd10604,17'd16319,17'd21984,17'd9189,17'd16549,17'd11135,17'd11670,17'd14518,17'd14518,17'd10476,17'd11130,17'd18444,17'd13883,17'd12576,17'd12256,17'd12256,17'd12859,17'd12416,17'd12254,17'd18564,17'd24207,17'd24208,17'd24209,17'd21361,17'd18681,17'd18444,17'd16442,17'd11959,17'd22819,17'd24033,17'd24033,17'd23515,17'd20314,17'd12996,17'd12115,17'd18682,17'd15810,17'd11806,17'd13882,17'd11960,17'd13883,17'd12996,17'd12262,17'd10989,17'd10989,17'd11964,17'd11522,17'd23172,17'd24210,17'd11524,17'd20754,17'd9472,17'd24037,17'd19415,17'd21984,17'd24211,17'd17472,17'd24212,17'd8885,17'd8412,17'd8247,17'd24213,17'd8578,17'd8413,17'd24214,17'd8577,17'd24215,17'd16333,17'd24216,17'd14269,17'd14012,17'd8586,17'd19783,17'd15695,17'd13771,17'd13771,17'd23523,17'd16570,17'd22136,17'd16570,17'd16570,17'd24217,17'd24218,17'd7465,17'd9893,17'd19650,17'd19650,17'd19650,17'd18088,17'd8588,17'd18336,17'd17487,17'd23351,17'd14144,17'd13896,17'd23189,17'd13012,17'd24219,17'd24220,17'd24221,17'd24222,17'd22840,17'd24223,17'd6198,17'd719,17'd17363,17'd24224,17'd24225,17'd23889,17'd24226,17'd24227,17'd24228,17'd24229,17'd24230,17'd24231,17'd23714,17'd23715,17'd24067,17'd24232,17'd24069,17'd24233,17'd24234,17'd24072,17'd24235,17'd24235,17'd24236,17'd24072,17'd24237,17'd24238,17'd23906,17'd24239,17'd24240,17'd24241,17'd24242,17'd24243,17'd24244,17'd23556,17'd23557,17'd24245,17'd24246,17'd24247,17'd23381,17'd24248,17'd23731,17'd24249,17'd24250,17'd24251,17'd24252,17'd23917,17'd24253,17'd24254,17'd23567,17'd24255,17'd24256,17'd24257,17'd24258,17'd24259,17'd24260,17'd24261,17'd24262,17'd24263,17'd24264,17'd24265,17'd24266,17'd24267,17'd24268,17'd24269,17'd24270,17'd24271,17'd24272,17'd24273,17'd24274,17'd24275,17'd24276,17'd24277,17'd24278,17'd24279,17'd23593,17'd24280,17'd24281,17'd19556,17'd24282,17'd24283,17'd24284,17'd24285,17'd24286,17'd24287,17'd24288,17'd24289,17'd23959,17'd24290,17'd24291,17'd22050,17'd24292,17'd24293,17'd24294,17'd19826,17'd20683,17'd20089,17'd21130,17'd20657,17'd24295,17'd23091,17'd22914,17'd21135,17'd24296,17'd24297,17'd21606,17'd24298,17'd22240,17'd24299,17'd24300,17'd24301,17'd24302,17'd24303,17'd22585,17'd22757,17'd24304,17'd24304,17'd24305,17'd24305,17'd22933,17'd24306,17'd23278,17'd8607,17'd10881,17'd8607,17'd23627,17'd24307,17'd24307,17'd23974,17'd6839,17'd7493,17'd24308,17'd4680,17'd4679,17'd4680,17'd4680,17'd24148,17'd24309,17'd7006,17'd7658,17'd6544,17'd7008,17'd23975,17'd6211,17'd23460,17'd24310,17'd23800,17'd24311,17'd11036,17'd11180,17'd11314,17'd14970,17'd17904,17'd15607,17'd15988,17'd18498,17'd18619,17'd18619,17'd24152,17'd17779,17'd17779,17'd15605,17'd14570,17'd16121,17'd19590,17'd21931,17'd24312,17'd20253,17'd24313,17'd24314,17'd24315,17'd24316,17'd22947,17'd18265,17'd15481,17'd14431,17'd19352,17'd24317,17'd24318,17'd24319,17'd24320,17'd24321,17'd24322,17'd18631,17'd430,17'd1678,17'd411,17'd24323,17'd7851,17'd1676,17'd5778,17'd14589,17'd2744,17'd2562,17'd24324,17'd24325,17'd24174,17'd23481,17'd23989,17'd5782,17'd24168,17'd24168,17'd23482,17'd23819,17'd24326,17'd24327,17'd24328,17'd24329,17'd24330,17'd7683,17'd9945,17'd8170,17'd8018,17'd8491,17'd8795,17'd8171,17'd7346,17'd7028,17'd5635,17'd4717,17'd4717,17'd9116,17'd3405,17'd7198,17'd22611,17'd24331,17'd24178,17'd24179,17'd24180,17'd24332,17'd23489,17'd24333,17'd15626
},
'{
17'd1688,17'd1831,17'd4247,17'd466,17'd13,17'd8814,17'd23,17'd6,17'd3753,17'd5205,17'd8040,17'd8040,17'd5793,17'd5793,17'd5793,17'd8040,17'd3594,17'd5,17'd24,17'd22,17'd5518,17'd5518,17'd22,17'd22,17'd5,17'd5,17'd5,17'd5,17'd1690,17'd1691,17'd285,17'd26,17'd27,17'd652,17'd4091,17'd3254,17'd2940,17'd3253,17'd23824,17'd22615,17'd1282,17'd1135,17'd16967,17'd17079,17'd1141,17'd1287,17'd1146,17'd24334,17'd3445,17'd12041,17'd6447,17'd6607,17'd24335,17'd24336,17'd12342,17'd24337,17'd24338,17'd24339,17'd24340,17'd17088,17'd18880,17'd18049,17'd24341,17'd24342,17'd24343,17'd24344,17'd16027,17'd16765,17'd11764,17'd11627,17'd12065,17'd24345,17'd22802,17'd14469,17'd12357,17'd12357,17'd12678,17'd13092,17'd12528,17'd24346,17'd12955,17'd14621,17'd24347,17'd12815,17'd11764,17'd11764,17'd10815,17'd18533,17'd19754,17'd11231,17'd24348,17'd24349,17'd24193,17'd14892,17'd15900,17'd24013,17'd24350,17'd18534,17'd16519,17'd17320,17'd17319,17'd19384,17'd15517,17'd10428,17'd6143,17'd6769,17'd6769,17'd7087,17'd8368,17'd8536,17'd7413,17'd24351,17'd8685,17'd10118,17'd9579,17'd9706,17'd9847,17'd9991,17'd10433,17'd10125,17'd24352,17'd17821,17'd17107,17'd16181,17'd14783,17'd9855,17'd23673,17'd24353,17'd24354,17'd24355,17'd23677,17'd24356,17'd19776,17'd24357,17'd21053,17'd12572,17'd24358,17'd23847,17'd24359,17'd21976,17'd12407,17'd12099,17'd11510,17'd16062,17'd24360,17'd11133,17'd20175,17'd9044,17'd24361,17'd19279,17'd12585,17'd15176,17'd10991,17'd10740,17'd10603,17'd14931,17'd13520,17'd12109,17'd14523,17'd16799,17'd14523,17'd12418,17'd12416,17'd12255,17'd23855,17'd24030,17'd24362,17'd24363,17'd19921,17'd18443,17'd16442,17'd21361,17'd19408,17'd23512,17'd12255,17'd20452,17'd21671,17'd18917,17'd18082,17'd17968,17'd12262,17'd11962,17'd11961,17'd11960,17'd11960,17'd16204,17'd11965,17'd10853,17'd20910,17'd11965,17'd18327,17'd14379,17'd17343,17'd24364,17'd17842,17'd24365,17'd16319,17'd9478,17'd9337,17'd15180,17'd24366,17'd10174,17'd9042,17'd24367,17'd24368,17'd8572,17'd9887,17'd9047,17'd8730,17'd8572,17'd8733,17'd17482,17'd11534,17'd13893,17'd12728,17'd24369,17'd13894,17'd14684,17'd24370,17'd24370,17'd24371,17'd24372,17'd24373,17'd15061,17'd10030,17'd16079,17'd14532,17'd14532,17'd20617,17'd14817,17'd13529,17'd24374,17'd16694,17'd15951,17'd24375,17'd24376,17'd16212,17'd24377,17'd24378,17'd24379,17'd23187,17'd23189,17'd10348,17'd11540,17'd24380,17'd24381,17'd23532,17'd24382,17'd14275,17'd889,17'd24383,17'd24384,17'd24385,17'd24386,17'd24387,17'd24388,17'd24389,17'd24390,17'd24391,17'd24392,17'd24393,17'd24394,17'd24395,17'd24069,17'd24396,17'd24397,17'd24398,17'd24399,17'd24400,17'd24401,17'd24400,17'd24402,17'd24403,17'd24403,17'd24403,17'd24237,17'd24404,17'd24405,17'd24406,17'd24407,17'd24408,17'd24409,17'd24410,17'd24079,17'd23913,17'd24411,17'd24412,17'd24413,17'd23730,17'd24414,17'd24415,17'd24416,17'd24417,17'd24418,17'd24419,17'd24420,17'd24421,17'd24422,17'd24423,17'd24424,17'd24425,17'd24426,17'd24427,17'd24428,17'd24429,17'd24430,17'd24431,17'd24432,17'd24433,17'd24434,17'd24435,17'd24436,17'd23411,17'd24437,17'd24438,17'd24439,17'd24440,17'd24111,17'd24441,17'd24441,17'd24442,17'd24443,17'd24444,17'd24445,17'd24446,17'd24447,17'd24448,17'd24449,17'd24450,17'd24451,17'd24452,17'd24453,17'd24454,17'd24455,17'd24456,17'd22374,17'd24457,17'd24458,17'd24459,17'd24460,17'd24461,17'd19688,17'd24462,17'd24463,17'd20355,17'd24464,17'd24465,17'd24466,17'd24467,17'd19452,17'd24468,17'd24469,17'd21138,17'd21299,17'd24470,17'd24471,17'd24472,17'd22242,17'd24473,17'd22412,17'd24474,17'd24474,17'd24474,17'd22585,17'd24305,17'd24305,17'd24306,17'd23278,17'd23457,17'd7493,17'd7493,17'd8607,17'd8607,17'd23974,17'd24475,17'd23974,17'd4678,17'd4679,17'd24476,17'd24477,17'd24478,17'd5912,17'd6381,17'd5322,17'd24479,17'd6702,17'd7324,17'd6702,17'd7008,17'd24480,17'd6211,17'd6382,17'd23630,17'd24481,17'd24482,17'd24482,17'd10237,17'd24483,17'd24484,17'd17655,17'd15606,17'd15606,17'd18620,17'd18499,17'd18259,17'd18499,17'd17903,17'd17903,17'd15605,17'd15093,17'd16247,17'd18260,17'd19985,17'd24485,17'd24486,17'd24487,17'd19989,17'd22425,17'd24488,17'd12313,17'd18028,17'd15481,17'd23292,17'd18137,17'd24489,17'd24490,17'd24491,17'd24492,17'd24493,17'd24494,17'd24495,17'd24496,17'd8483,17'd190,17'd24497,17'd1393,17'd18272,17'd24498,17'd14589,17'd14738,17'd24499,17'd24500,17'd23818,17'd23994,17'd24501,17'd24502,17'd24329,17'd23995,17'd24174,17'd24174,17'd24328,17'd24503,17'd24503,17'd24504,17'd23819,17'd5781,17'd7683,17'd23483,17'd7854,17'd7854,17'd8491,17'd8795,17'd8171,17'd8169,17'd5365,17'd5635,17'd5501,17'd7193,17'd7689,17'd3405,17'd24505,17'd22441,17'd22442,17'd24178,17'd24506,17'd24507,17'd24332,17'd24332,17'd180,17'd24333
},
'{
17'd3250,17'd2422,17'd1688,17'd466,17'd12,17'd8814,17'd23,17'd6,17'd5205,17'd5205,17'd8040,17'd8040,17'd5793,17'd5793,17'd5793,17'd5205,17'd5,17'd5,17'd23,17'd22,17'd5518,17'd5518,17'd5518,17'd22,17'd5,17'd24,17'd24,17'd5,17'd1690,17'd1691,17'd285,17'd286,17'd28,17'd29,17'd3755,17'd3254,17'd2940,17'd3253,17'd23824,17'd24508,17'd16966,17'd1282,17'd1135,17'd1139,17'd1426,17'd24509,17'd24510,17'd12791,17'd4903,17'd24511,17'd6447,17'd6607,17'd24512,17'd22455,17'd24513,17'd24514,17'd20020,17'd24515,17'd19509,17'd14200,17'd18880,17'd24188,17'd24516,17'd24517,17'd24518,17'd24519,17'd16765,17'd16658,17'd11764,17'd11627,17'd12065,17'd24345,17'd15763,17'd12357,17'd12357,17'd12678,17'd13092,17'd12679,17'd12217,17'd12814,17'd12218,17'd13094,17'd12815,17'd11913,17'd11913,17'd11629,17'd11087,17'd16766,17'd15765,17'd17319,17'd24520,17'd24521,17'd15385,17'd14892,17'd15900,17'd16520,17'd19009,17'd19129,17'd16519,17'd17320,17'd17319,17'd16164,17'd15517,17'd9300,17'd7418,17'd7418,17'd6141,17'd6141,17'd7417,17'd7417,17'd7411,17'd10117,17'd24522,17'd24523,17'd9163,17'd24524,17'd9707,17'd9849,17'd10291,17'd10126,17'd24525,17'd16668,17'd16048,17'd13858,17'd9996,17'd24526,17'd24527,17'd24528,17'd24529,17'd11251,17'd11940,17'd11944,17'd24530,17'd24357,17'd21499,17'd24531,17'd24532,17'd24358,17'd24533,17'd21976,17'd13248,17'd24534,17'd24535,17'd24536,17'd19156,17'd9884,17'd9192,17'd8720,17'd14674,17'd14383,17'd19919,17'd21206,17'd10475,17'd10740,17'd10603,17'd11519,17'd11960,17'd12253,17'd15811,17'd14930,17'd14809,17'd12417,17'd12255,17'd23681,17'd24537,17'd24538,17'd24539,17'd14259,17'd19158,17'd16442,17'd21361,17'd21505,17'd23512,17'd24030,17'd23855,17'd12253,17'd13883,17'd16204,17'd17968,17'd17968,17'd13362,17'd11806,17'd11960,17'd13883,17'd13135,17'd12262,17'd20910,17'd10738,17'd10853,17'd10989,17'd17478,17'd24540,17'd24541,17'd17966,17'd24542,17'd17719,17'd10742,17'd18332,17'd16793,17'd24543,17'd24361,17'd10336,17'd24544,17'd8884,17'd16562,17'd8412,17'd24545,17'd24546,17'd24547,17'd11811,17'd16691,17'd10860,17'd24548,17'd15058,17'd14141,17'd18568,17'd16693,17'd24549,17'd24550,17'd10030,17'd16079,17'd12729,17'd8428,17'd24551,17'd13770,17'd14678,17'd14678,17'd14678,17'd24552,17'd24553,17'd16692,17'd13894,17'd12729,17'd7462,17'd24554,17'd7794,17'd15696,17'd15815,17'd24555,17'd23000,17'd24556,17'd24557,17'd24558,17'd24559,17'd24560,17'd10188,17'd16699,17'd24561,17'd19292,17'd24562,17'd24563,17'd24564,17'd24565,17'd24387,17'd24566,17'd24567,17'd24568,17'd24569,17'd24570,17'd24571,17'd24572,17'd24573,17'd24234,17'd24574,17'd24398,17'd24575,17'd24576,17'd24398,17'd24399,17'd24402,17'd24402,17'd24577,17'd24578,17'd24578,17'd24403,17'd24237,17'd24404,17'd24579,17'd24580,17'd24581,17'd24582,17'd24583,17'd24584,17'd24078,17'd24585,17'd24586,17'd24587,17'd24588,17'd24589,17'd24590,17'd24415,17'd24252,17'd24417,17'd24417,17'd24248,17'd24591,17'd23209,17'd24592,17'd24593,17'd24594,17'd24595,17'd24596,17'd24597,17'd24598,17'd24599,17'd24600,17'd24601,17'd24602,17'd24603,17'd24604,17'd22704,17'd24605,17'd24606,17'd24432,17'd24437,17'd24607,17'd24608,17'd24609,17'd24610,17'd24611,17'd24442,17'd24612,17'd24613,17'd24614,17'd24615,17'd24616,17'd24617,17'd24618,17'd24619,17'd24620,17'd24621,17'd24622,17'd24623,17'd24624,17'd24625,17'd24626,17'd24627,17'd24628,17'd24629,17'd24630,17'd24631,17'd19687,17'd19578,17'd19822,17'd20087,17'd20218,17'd24632,17'd24633,17'd18962,17'd18487,17'd24634,17'd24635,17'd19817,17'd24636,17'd24637,17'd20991,17'd21922,17'd24638,17'd24639,17'd24640,17'd24641,17'd24474,17'd24474,17'd22585,17'd24642,17'd24305,17'd24643,17'd24306,17'd24644,17'd8911,17'd8289,17'd24645,17'd7493,17'd7006,17'd24309,17'd24646,17'd24148,17'd4679,17'd24477,17'd24647,17'd24648,17'd4992,17'd5323,17'd24649,17'd24650,17'd6702,17'd7324,17'd7324,17'd6545,17'd24480,17'd6547,17'd6382,17'd6384,17'd23461,17'd24651,17'd6706,17'd6852,17'd24652,17'd24653,17'd24654,17'd17904,17'd15726,17'd18742,17'd24655,17'd18259,17'd18499,17'd17903,17'd17779,17'd15605,17'd15093,17'd16247,17'd19590,17'd19847,17'd23464,17'd24656,17'd16372,17'd24153,17'd24657,17'd24658,17'd24659,17'd16958,17'd15732,17'd24660,17'd13929,17'd19486,17'd4385,17'd24661,17'd24662,17'd24663,17'd24664,17'd24665,17'd24666,17'd1957,17'd1823,17'd24323,17'd7027,17'd5942,17'd24498,17'd14589,17'd24667,17'd24499,17'd24668,17'd24669,17'd24501,17'd24670,17'd24670,17'd24170,17'd23995,17'd24329,17'd24170,17'd24671,17'd24672,17'd24672,17'd24504,17'd23819,17'd5781,17'd7515,17'd23483,17'd7854,17'd7854,17'd8491,17'd8795,17'd8171,17'd8169,17'd5365,17'd5635,17'd5501,17'd4717,17'd9116,17'd3405,17'd24505,17'd22441,17'd22612,17'd6880,17'd21791,17'd24507,17'd24332,17'd24332,17'd180,17'd24333
},
'{
17'd2592,17'd2422,17'd1831,17'd466,17'd2423,17'd8814,17'd23,17'd6,17'd5205,17'd5205,17'd5205,17'd3753,17'd3753,17'd3753,17'd3753,17'd3753,17'd5,17'd5,17'd23,17'd22,17'd20,17'd20,17'd5518,17'd22,17'd23,17'd23,17'd1691,17'd1691,17'd1691,17'd1691,17'd285,17'd26,17'd7060,17'd4430,17'd3908,17'd3254,17'd2940,17'd3253,17'd23824,17'd24508,17'd1839,17'd1283,17'd1424,17'd1139,17'd24673,17'd24509,17'd24674,17'd24675,17'd24676,17'd24677,17'd24678,17'd23663,17'd7073,17'd23145,17'd23319,17'd24006,17'd24679,17'd24515,17'd24680,17'd17674,17'd24681,17'd15254,17'd24682,17'd24683,17'd24684,17'd24519,17'd16765,17'd13969,17'd13840,17'd12814,17'd12217,17'd12527,17'd12357,17'd12357,17'd12678,17'd12678,17'd12527,17'd12955,17'd12814,17'd12360,17'd12218,17'd24347,17'd12362,17'd11764,17'd12531,17'd17204,17'd17205,17'd21964,17'd16164,17'd16169,17'd18059,17'd24685,17'd14768,17'd14892,17'd15386,17'd24686,17'd24687,17'd24688,17'd16519,17'd16519,17'd16289,17'd16164,17'd10429,17'd9440,17'd7418,17'd5409,17'd6626,17'd6626,17'd6305,17'd10695,17'd9305,17'd9012,17'd8695,17'd9163,17'd9015,17'd9165,17'd9445,17'd9584,17'd19901,17'd18787,17'd16668,17'd16182,17'd21972,17'd24689,17'd21973,17'd24690,17'd24691,17'd24692,17'd24693,17'd24694,17'd12098,17'd24695,17'd24696,17'd24697,17'd24531,17'd24698,17'd24532,17'd24699,17'd24700,17'd21976,17'd16903,17'd11509,17'd24701,17'd24702,17'd9883,17'd23679,17'd9043,17'd10174,17'd11809,17'd11135,17'd12423,17'd11399,17'd16555,17'd24703,17'd10852,17'd11666,17'd15184,17'd18564,17'd15811,17'd22297,17'd14526,17'd12417,17'd23681,17'd24704,17'd24537,17'd24705,17'd24706,17'd17478,17'd19158,17'd16325,17'd19408,17'd23515,17'd24030,17'd24707,17'd16324,17'd15184,17'd12996,17'd12262,17'd17968,17'd12262,17'd13135,17'd11960,17'd11960,17'd13135,17'd13762,17'd10989,17'd24708,17'd24703,17'd10604,17'd12720,17'd11521,17'd23337,17'd12423,17'd24709,17'd10024,17'd11136,17'd10742,17'd18324,17'd16065,17'd15298,17'd8874,17'd8874,17'd9621,17'd8885,17'd16562,17'd9744,17'd24710,17'd24711,17'd24712,17'd24713,17'd17241,17'd11534,17'd24714,17'd7294,17'd7791,17'd24552,17'd10862,17'd13378,17'd24369,17'd24715,17'd8111,17'd8111,17'd7624,17'd14678,17'd14141,17'd11141,17'd12728,17'd14391,17'd24716,17'd16210,17'd17018,17'd17018,17'd14012,17'd18568,17'd15950,17'd24370,17'd18087,17'd13771,17'd20052,17'd24717,17'd24718,17'd24719,17'd23184,17'd24720,17'd10348,17'd10349,17'd10350,17'd16699,17'd24721,17'd24722,17'd24723,17'd24724,17'd24725,17'd24726,17'd24727,17'd24728,17'd24729,17'd24730,17'd24731,17'd24573,17'd24732,17'd24732,17'd24071,17'd24236,17'd24574,17'd24398,17'd24398,17'd24398,17'd24398,17'd24399,17'd24733,17'd24733,17'd24578,17'd24403,17'd24237,17'd24237,17'd24734,17'd24579,17'd23907,17'd23719,17'd24735,17'd24736,17'd24736,17'd24737,17'd24078,17'd23911,17'd24738,17'd24739,17'd24740,17'd24741,17'd24742,17'd24743,17'd24744,17'd24745,17'd24590,17'd24083,17'd24084,17'd23918,17'd24746,17'd24747,17'd24748,17'd24749,17'd24750,17'd24751,17'd24752,17'd24753,17'd24754,17'd24755,17'd24756,17'd24757,17'd24758,17'd24759,17'd24760,17'd24432,17'd24437,17'd24761,17'd24762,17'd24763,17'd24764,17'd24765,17'd24766,17'd24767,17'd24768,17'd24769,17'd24770,17'd24771,17'd24772,17'd24773,17'd24774,17'd24775,17'd24776,17'd24777,17'd24778,17'd24779,17'd22901,17'd24780,17'd24781,17'd24782,17'd24782,17'd24783,17'd24784,17'd19459,17'd19469,17'd19957,17'd20238,17'd24785,17'd19683,17'd24786,17'd17771,17'd16830,17'd17396,17'd17767,17'd19328,17'd24787,17'd18727,17'd24788,17'd24789,17'd21608,17'd21923,17'd24790,17'd24790,17'd24791,17'd24641,17'd24474,17'd24642,17'd24642,17'd24792,17'd24643,17'd23109,17'd24793,17'd24794,17'd11294,17'd8143,17'd6702,17'd6381,17'd24795,17'd24795,17'd24796,17'd5912,17'd24648,17'd24797,17'd5608,17'd4993,17'd5325,17'd5323,17'd5323,17'd24649,17'd24798,17'd5323,17'd5607,17'd24480,17'd6212,17'd5610,17'd24799,17'd24800,17'd6388,17'd6707,17'd10237,17'd24801,17'd24802,17'd15340,17'd24803,17'd22420,17'd18620,17'd20541,17'd22421,17'd17779,17'd17065,17'd17065,17'd16371,17'd16247,17'd19590,17'd19847,17'd23464,17'd20849,17'd24804,17'd24313,17'd24805,17'd11859,17'd24316,17'd24806,17'd16378,17'd15732,17'd22771,17'd24807,17'd24808,17'd24809,17'd24810,17'd24811,17'd24812,17'd24813,17'd927,17'd8639,17'd190,17'd2577,17'd8165,17'd24814,17'd14179,17'd14859,17'd14978,17'd24499,17'd24668,17'd24815,17'd24816,17'd24171,17'd23993,17'd24817,17'd24818,17'd24819,17'd24820,17'd24821,17'd24822,17'd24822,17'd24823,17'd24173,17'd24824,17'd23135,17'd24176,17'd7854,17'd7854,17'd23302,17'd8491,17'd9944,17'd24825,17'd24826,17'd16624,17'd5635,17'd6575,17'd7030,17'd3720,17'd24827,17'd22441,17'd23310,17'd24828,17'd24829,17'd2253,17'd24332,17'd24332,17'd180,17'd24333
},
'{
17'd2784,17'd2935,17'd1831,17'd466,17'd2423,17'd15494,17'd24,17'd6,17'd3753,17'd3753,17'd3753,17'd3753,17'd3753,17'd3753,17'd3753,17'd3753,17'd24,17'd24,17'd23,17'd22,17'd20,17'd2598,17'd5518,17'd22,17'd23,17'd23,17'd1691,17'd1691,17'd1691,17'd467,17'd285,17'd27,17'd4430,17'd4091,17'd3595,17'd3254,17'd2940,17'd3253,17'd2785,17'd2600,17'd1702,17'd1423,17'd1704,17'd1705,17'd24830,17'd24831,17'd24832,17'd24833,17'd24834,17'd24835,17'd6755,17'd23663,17'd12042,17'd24004,17'd23496,17'd20284,17'd24836,17'd14199,17'd24837,17'd24838,17'd18162,17'd15505,17'd24839,17'd24840,17'd24684,17'd24519,17'd16658,17'd13969,17'd12530,17'd12814,17'd24345,17'd12527,17'd12357,17'd12357,17'd12678,17'd13092,17'd13093,17'd12065,17'd13464,17'd11627,17'd12957,17'd12957,17'd11913,17'd11629,17'd17317,17'd16766,17'd16986,17'd20735,17'd16659,17'd16411,17'd18059,17'd17321,17'd14346,17'd15386,17'd15260,17'd15768,17'd19256,17'd16519,17'd16519,17'd19256,17'd16164,17'd15766,17'd9703,17'd7582,17'd6624,17'd5689,17'd6305,17'd9008,17'd24841,17'd8382,17'd8383,17'd8383,17'd24842,17'd24843,17'd12685,17'd11920,17'd9446,17'd9708,17'd17702,17'd17945,17'd24844,17'd24845,17'd24846,17'd24847,17'd24848,17'd21197,17'd23159,17'd24849,17'd14657,17'd12570,17'd20904,17'd24850,17'd24696,17'd23844,17'd24851,17'd24852,17'd14923,17'd12402,17'd22126,17'd21202,17'd11655,17'd24853,17'd24854,17'd10476,17'd11136,17'd20757,17'd9043,17'd15187,17'd19531,17'd12585,17'd12423,17'd21206,17'd16555,17'd10738,17'd10736,17'd11961,17'd15434,17'd16913,17'd19534,17'd24855,17'd13517,17'd14003,17'd23511,17'd24856,17'd24857,17'd23170,17'd24858,17'd21985,17'd16442,17'd22992,17'd22819,17'd23856,17'd24859,17'd24030,17'd21671,17'd13883,17'd12262,17'd18560,17'd12115,17'd16204,17'd13883,17'd13761,17'd13883,17'd12996,17'd11965,17'd20910,17'd24708,17'd10739,17'd24860,17'd15182,17'd16068,17'd11668,17'd13522,17'd9884,17'd11277,17'd23340,17'd10857,17'd10744,17'd24861,17'd9346,17'd8874,17'd10175,17'd17607,17'd9195,17'd8412,17'd8247,17'd8576,17'd24862,17'd24863,17'd11812,17'd12265,17'd15192,17'd15191,17'd13769,17'd11141,17'd14009,17'd16210,17'd24864,17'd24865,17'd24866,17'd24867,17'd24868,17'd18086,17'd7458,17'd14269,17'd17018,17'd24869,17'd24870,17'd20318,17'd24871,17'd16448,17'd24716,17'd24872,17'd8891,17'd24369,17'd13894,17'd19648,17'd15306,17'd24873,17'd24874,17'd19540,17'd17243,17'd18456,17'd8433,17'd24875,17'd11819,17'd24876,17'd13260,17'd24877,17'd24878,17'd24879,17'd24880,17'd24881,17'd24882,17'd24883,17'd24884,17'd24885,17'd24886,17'd24887,17'd24888,17'd24732,17'd24732,17'd24071,17'd24236,17'd24889,17'd24399,17'd24399,17'd24399,17'd24399,17'd24399,17'd24733,17'd24733,17'd24403,17'd24403,17'd24237,17'd24890,17'd24734,17'd24579,17'd23907,17'd24239,17'd24735,17'd24735,17'd24736,17'd24891,17'd24892,17'd23910,17'd24585,17'd24586,17'd24893,17'd24894,17'd24895,17'd24896,17'd24897,17'd24898,17'd24899,17'd24900,17'd24901,17'd24902,17'd24903,17'd24904,17'd24905,17'd24906,17'd24907,17'd21248,17'd23229,17'd24908,17'd24909,17'd24910,17'd24911,17'd24912,17'd23591,17'd24913,17'd24760,17'd24914,17'd24915,17'd24916,17'd24912,17'd24917,17'd24918,17'd24919,17'd24920,17'd24921,17'd24922,17'd24923,17'd24924,17'd24925,17'd21256,17'd24926,17'd24927,17'd24774,17'd24928,17'd24284,17'd24929,17'd24930,17'd24931,17'd24932,17'd24933,17'd24934,17'd24934,17'd19455,17'd19685,17'd19206,17'd24935,17'd24936,17'd24785,17'd24937,17'd19473,17'd19567,17'd17518,17'd17519,17'd17388,17'd17388,17'd24938,17'd19078,17'd19078,17'd18954,17'd24939,17'd24789,17'd24940,17'd24941,17'd21923,17'd24790,17'd24640,17'd24641,17'd24942,17'd24642,17'd24943,17'd24943,17'd24306,17'd23454,17'd24794,17'd7823,17'd7163,17'd6544,17'd5912,17'd6381,17'd24795,17'd24796,17'd5912,17'd5607,17'd24944,17'd5326,17'd5150,17'd5480,17'd5325,17'd4992,17'd24649,17'd24649,17'd24649,17'd4992,17'd24480,17'd23799,17'd5479,17'd5759,17'd5760,17'd5760,17'd6387,17'd6852,17'd24483,17'd24945,17'd17655,17'd16956,17'd15476,17'd18742,17'd20541,17'd22421,17'd17779,17'd17065,17'd17065,17'd17065,17'd16371,17'd18134,17'd20384,17'd19847,17'd21773,17'd22944,17'd17409,17'd23981,17'd20548,17'd24946,17'd24947,17'd19351,17'd16254,17'd23292,17'd18748,17'd22772,17'd24948,17'd24949,17'd24950,17'd24951,17'd24952,17'd24953,17'd1961,17'd190,17'd2922,17'd8165,17'd1392,17'd3223,17'd24954,17'd2561,17'd24955,17'd24668,17'd24956,17'd24171,17'd24956,17'd23993,17'd24957,17'd24958,17'd24959,17'd24173,17'd24960,17'd24822,17'd24961,17'd24823,17'd24173,17'd24962,17'd24963,17'd7683,17'd7854,17'd7514,17'd7855,17'd23302,17'd17294,17'd17073,17'd24964,17'd16740,17'd5635,17'd5635,17'd6576,17'd4564,17'd24827,17'd22441,17'd23655,17'd24965,17'd24966,17'd2253,17'd24332,17'd24332,17'd180,17'd180
},
'{
17'd4733,17'd14743,17'd1831,17'd1127,17'd2423,17'd15494,17'd24,17'd3753,17'd3753,17'd3753,17'd3753,17'd3753,17'd3753,17'd3753,17'd3753,17'd3753,17'd24,17'd23,17'd23,17'd22,17'd20,17'd2598,17'd5518,17'd22,17'd23,17'd23,17'd1691,17'd1691,17'd467,17'd285,17'd285,17'd27,17'd4430,17'd4248,17'd3908,17'd3433,17'd3256,17'd3253,17'd2785,17'd2785,17'd19874,17'd1422,17'd2267,17'd24967,17'd24830,17'd24968,17'd24969,17'd3444,17'd11894,17'd11613,17'd6755,17'd6756,17'd11895,17'd22974,17'd13194,17'd20878,17'd24836,17'd24970,17'd24971,17'd14996,17'd24972,17'd24973,17'd24974,17'd23153,17'd24344,17'd24344,17'd16163,17'd15764,17'd12530,17'd12065,17'd12679,17'd12527,17'd14469,17'd12357,17'd12678,17'd13092,17'd12955,17'd12814,17'd12956,17'd12956,17'd24975,17'd11913,17'd12531,17'd11629,17'd17689,17'd16986,17'd21808,17'd19256,17'd24348,17'd16033,17'd24192,17'd16768,17'd16290,17'd16769,17'd16769,17'd16769,17'd15899,17'd20585,17'd16880,17'd15898,17'd15517,17'd10429,17'd9159,17'd5409,17'd10946,17'd10695,17'd24976,17'd24977,17'd24978,17'd7760,17'd24979,17'd24980,17'd13612,17'd14640,17'd8703,17'd9314,17'd17583,17'd16997,17'd16668,17'd24844,17'd16046,17'd12963,17'd24981,17'd24982,17'd9858,17'd24983,17'd24984,17'd15667,17'd24985,17'd23335,17'd24530,17'd24986,17'd24987,17'd11943,17'd24988,17'd17833,17'd12406,17'd12244,17'd13997,17'd11795,17'd24989,17'd24990,17'd17009,17'd9883,17'd9191,17'd15682,17'd9346,17'd15048,17'd10479,17'd11400,17'd21206,17'd21206,17'd10475,17'd10737,17'd11962,17'd12110,17'd16685,17'd16913,17'd21504,17'd13515,17'd14003,17'd19534,17'd24991,17'd24856,17'd24992,17'd24993,17'd23513,17'd24994,17'd21361,17'd19408,17'd20452,17'd23681,17'd24859,17'd23168,17'd24995,17'd15185,17'd12115,17'd18560,17'd12262,17'd13135,17'd11960,17'd11960,17'd15185,17'd11964,17'd20451,17'd20910,17'd10854,17'd10990,17'd12720,17'd24035,17'd11524,17'd24996,17'd9741,17'd11809,17'd9340,17'd11809,17'd24997,17'd24998,17'd24998,17'd9344,17'd10174,17'd8720,17'd24999,17'd8724,17'd9744,17'd17481,17'd21987,17'd24862,17'd23343,17'd17352,17'd8255,17'd16801,17'd25000,17'd25001,17'd14938,17'd14140,17'd13377,17'd25002,17'd25003,17'd25004,17'd25005,17'd25005,17'd13377,17'd15439,17'd13893,17'd16567,17'd10747,17'd10747,17'd16567,17'd18921,17'd18921,17'd19536,17'd14269,17'd15194,17'd7956,17'd14678,17'd19648,17'd25006,17'd15306,17'd22136,17'd15062,17'd15063,17'd14819,17'd25007,17'd25008,17'd25009,17'd8438,17'd25010,17'd25011,17'd25012,17'd25013,17'd25014,17'd25015,17'd25016,17'd25017,17'd25018,17'd24571,17'd25019,17'd24888,17'd24888,17'd24234,17'd25020,17'd24071,17'd24236,17'd24890,17'd24403,17'd24403,17'd25021,17'd24237,17'd24237,17'd25022,17'd25022,17'd25023,17'd24237,17'd25024,17'd24404,17'd25025,17'd24405,17'd24580,17'd23719,17'd24582,17'd24582,17'd23908,17'd24891,17'd24892,17'd23910,17'd23911,17'd23725,17'd25026,17'd25027,17'd25028,17'd24893,17'd25029,17'd25030,17'd25031,17'd25032,17'd24246,17'd24743,17'd25033,17'd25034,17'd25035,17'd25036,17'd25037,17'd25038,17'd25039,17'd25040,17'd25041,17'd25042,17'd25043,17'd25044,17'd25045,17'd25046,17'd25047,17'd25048,17'd24915,17'd25049,17'd24916,17'd25050,17'd25051,17'd25052,17'd25053,17'd25054,17'd25055,17'd25056,17'd25057,17'd25058,17'd25059,17'd25060,17'd25061,17'd25062,17'd25062,17'd25063,17'd25064,17'd25065,17'd25066,17'd25067,17'd25068,17'd25069,17'd25069,17'd25070,17'd25070,17'd19571,17'd25071,17'd19570,17'd20527,17'd20373,17'd19069,17'd18127,17'd17649,17'd25072,17'd17388,17'd25073,17'd25074,17'd25075,17'd25076,17'd18613,17'd17167,17'd16356,17'd25077,17'd25078,17'd25079,17'd25080,17'd24790,17'd22243,17'd24942,17'd24942,17'd25081,17'd22758,17'd23278,17'd23109,17'd23279,17'd11158,17'd25082,17'd7326,17'd7007,17'd6545,17'd24796,17'd5322,17'd24649,17'd5607,17'd25083,17'd5479,17'd5478,17'd5150,17'd4993,17'd5325,17'd5324,17'd5324,17'd24649,17'd4992,17'd5608,17'd25083,17'd5479,17'd5759,17'd5760,17'd5760,17'd6388,17'd6706,17'd25084,17'd25085,17'd14970,17'd14971,17'd17655,17'd22420,17'd20695,17'd25086,17'd17779,17'd17065,17'd17065,17'd16371,17'd18498,17'd18134,17'd20384,17'd19847,17'd19714,17'd25087,17'd25088,17'd21933,17'd25089,17'd12311,17'd12312,17'd17071,17'd25090,17'd14431,17'd25091,17'd25092,17'd25093,17'd25094,17'd25095,17'd25096,17'd25097,17'd25098,17'd1379,17'd8812,17'd2922,17'd2576,17'd1677,17'd24498,17'd1385,17'd12645,17'd24499,17'd24668,17'd25099,17'd25100,17'd25099,17'd25101,17'd24173,17'd24820,17'd24328,17'd24671,17'd24823,17'd24961,17'd25102,17'd25103,17'd24328,17'd25104,17'd25105,17'd23820,17'd25106,17'd25106,17'd25107,17'd23483,17'd25108,17'd25109,17'd24964,17'd16740,17'd4065,17'd5635,17'd6724,17'd4564,17'd24827,17'd25110,17'd25111,17'd25112,17'd25113,17'd2415,17'd24000,17'd24332,17'd15355,17'd15355
},
'{
17'd6420,17'd15746,17'd3252,17'd1127,17'd2423,17'd10260,17'd24,17'd3753,17'd3753,17'd3594,17'd3594,17'd3753,17'd3753,17'd3753,17'd3753,17'd6,17'd23,17'd23,17'd23,17'd22,17'd20,17'd2598,17'd5518,17'd22,17'd23,17'd23,17'd1832,17'd1832,17'd285,17'd285,17'd27,17'd27,17'd4248,17'd3908,17'd3433,17'd3254,17'd2940,17'd2940,17'd2602,17'd2263,17'd19874,17'd1976,17'd3107,17'd4583,17'd4257,17'd25114,17'd3269,17'd25115,17'd25116,17'd6606,17'd7565,17'd24335,17'd22455,17'd23829,17'd22623,17'd25117,17'd25118,17'd19886,17'd25119,17'd25120,17'd15372,17'd25121,17'd25122,17'd25123,17'd24344,17'd24344,17'd16027,17'd14622,17'd12218,17'd11626,17'd12527,17'd12527,17'd14469,17'd14469,17'd13092,17'd12679,17'd12065,17'd12956,17'd11229,17'd25124,17'd24975,17'd11913,17'd11629,17'd17204,17'd18174,17'd21650,17'd18658,17'd18776,17'd15902,17'd15902,17'd16987,17'd16987,17'd15524,17'd15645,17'd15645,17'd24348,17'd20585,17'd20585,17'd15766,17'd15898,17'd15517,17'd9440,17'd7750,17'd5255,17'd10695,17'd9842,17'd24977,17'd25125,17'd7920,17'd25126,17'd25127,17'd25128,17'd10293,17'd10293,17'd25129,17'd16891,17'd16667,17'd16782,17'd25130,17'd25131,17'd25132,17'd11367,17'd25133,17'd25134,17'd25135,17'd25136,17'd17958,17'd13871,17'd24851,17'd18912,17'd22810,17'd25137,17'd11945,17'd11941,17'd25138,17'd16902,17'd22126,17'd12097,17'd18912,17'd25139,17'd25140,17'd25141,17'd25142,17'd10743,17'd9189,17'd8874,17'd9479,17'd10479,17'd19282,17'd21206,17'd21206,17'd21206,17'd10990,17'd11395,17'd11960,17'd15434,17'd12415,17'd19534,17'd14003,17'd14003,17'd19534,17'd24991,17'd24856,17'd24538,17'd24539,17'd24858,17'd25143,17'd14258,17'd19408,17'd23168,17'd23511,17'd23511,17'd24707,17'd23168,17'd19920,17'd11964,17'd17968,17'd12262,17'd12996,17'd11806,17'd13883,17'd13135,17'd11964,17'd11965,17'd25144,17'd20910,17'd11808,17'd14673,17'd17838,17'd17236,17'd19282,17'd16796,17'd15048,17'd9346,17'd9346,17'd9340,17'd25145,17'd25146,17'd9479,17'd22814,17'd8874,17'd9045,17'd23861,17'd8409,17'd9349,17'd8573,17'd25147,17'd25148,17'd17352,17'd11968,17'd25149,17'd25150,17'd25151,17'd12590,17'd21508,17'd14681,17'd22134,17'd25152,17'd15693,17'd12265,17'd12265,17'd13649,17'd25152,17'd15948,17'd16804,17'd10341,17'd19781,17'd19781,17'd15439,17'd13377,17'd8890,17'd25153,17'd25154,17'd25153,17'd14268,17'd25155,17'd14815,17'd18568,17'd12267,17'd12729,17'd14142,17'd18333,17'd19540,17'd18206,17'd25156,17'd25157,17'd25158,17'd12873,17'd25159,17'd25160,17'd25161,17'd25162,17'd25163,17'd25164,17'd25165,17'd25166,17'd25167,17'd24888,17'd25168,17'd25168,17'd24072,17'd24072,17'd24236,17'd24400,17'd25169,17'd25169,17'd25170,17'd25021,17'd25171,17'd24237,17'd24399,17'd24399,17'd25023,17'd24890,17'd24237,17'd24404,17'd24734,17'd24579,17'd23904,17'd24580,17'd25172,17'd24582,17'd24736,17'd24891,17'd23909,17'd24078,17'd23724,17'd25173,17'd25174,17'd25175,17'd25176,17'd25176,17'd25177,17'd25178,17'd25179,17'd25180,17'd24893,17'd23914,17'd24415,17'd25181,17'd25182,17'd25183,17'd25184,17'd24099,17'd25185,17'd25186,17'd25187,17'd25188,17'd25189,17'd25190,17'd24757,17'd23758,17'd25047,17'd24271,17'd25191,17'd25192,17'd25191,17'd25193,17'd25194,17'd25195,17'd25196,17'd25054,17'd25197,17'd25198,17'd25199,17'd25200,17'd25201,17'd25202,17'd25203,17'd25204,17'd25205,17'd25206,17'd23954,17'd25207,17'd25208,17'd25209,17'd25210,17'd25211,17'd25212,17'd25212,17'd25213,17'd19075,17'd19705,17'd19841,17'd20373,17'd19818,17'd19077,17'd18735,17'd25214,17'd17270,17'd17388,17'd19323,17'd25215,17'd25216,17'd25217,17'd25076,17'd18613,17'd16832,17'd25218,17'd24789,17'd25078,17'd25219,17'd24790,17'd24790,17'd22243,17'd25220,17'd25221,17'd25221,17'd22758,17'd25222,17'd24793,17'd25223,17'd25082,17'd25224,17'd7008,17'd6545,17'd5912,17'd6381,17'd24649,17'd5607,17'd5326,17'd5610,17'd5611,17'd4844,17'd5478,17'd4993,17'd4993,17'd5325,17'd5323,17'd4992,17'd5608,17'd24944,17'd5326,17'd25225,17'd5759,17'd5482,17'd5332,17'd6387,17'd6392,17'd25226,17'd13406,17'd14970,17'd15094,17'd15476,17'd21453,17'd20541,17'd17065,17'd17065,17'd17065,17'd16371,17'd18498,17'd18741,17'd20384,17'd19847,17'd19714,17'd20849,17'd20116,17'd25227,17'd25228,17'd19852,17'd25229,17'd25230,17'd25231,17'd15100,17'd25232,17'd18506,17'd25233,17'd22260,17'd25234,17'd25235,17'd25236,17'd25237,17'd792,17'd1380,17'd2764,17'd6888,17'd7027,17'd5498,17'd25238,17'd2243,17'd24955,17'd24668,17'd25099,17'd25099,17'd25239,17'd25101,17'd24328,17'd24328,17'd25240,17'd24504,17'd24823,17'd24961,17'd25102,17'd25241,17'd25240,17'd25104,17'd25105,17'd23996,17'd7515,17'd7515,17'd23654,17'd25107,17'd25242,17'd25243,17'd24964,17'd3717,17'd4233,17'd5635,17'd6724,17'd4564,17'd4565,17'd20267,17'd23655,17'd25244,17'd25245,17'd25246,17'd24000,17'd24332,17'd21165,17'd21165
},
'{
17'd4892,17'd6420,17'd14070,17'd1127,17'd2423,17'd10260,17'd24,17'd3753,17'd3753,17'd3753,17'd6,17'd6,17'd6,17'd6,17'd3753,17'd3594,17'd284,17'd22,17'd21,17'd21,17'd20,17'd20,17'd22,17'd23,17'd23,17'd23,17'd1832,17'd1832,17'd285,17'd285,17'd27,17'd980,17'd4248,17'd4090,17'd3909,17'd3433,17'd3256,17'd2940,17'd2601,17'd2263,17'd19874,17'd2431,17'd3107,17'd4583,17'd25247,17'd25114,17'd12790,17'd25248,17'd25116,17'd11613,17'd24678,17'd23494,17'd22621,17'd25249,17'd25250,17'd25251,17'd25252,17'd25253,17'd25254,17'd25255,17'd25256,17'd25257,17'd24684,17'd14622,17'd23324,17'd24344,17'd16027,17'd14470,17'd13211,17'd13093,17'd12527,17'd12527,17'd14469,17'd13462,17'd13092,17'd13209,17'd14890,17'd12530,17'd12956,17'd10690,17'd12680,17'd11913,17'd11362,17'd25258,17'd18174,17'd21808,17'd18060,17'd17810,17'd16033,17'd16987,17'd16290,17'd16290,17'd18534,17'd19256,17'd19256,17'd20585,17'd16880,17'd10113,17'd9703,17'd9703,17'd10694,17'd8537,17'd6468,17'd6140,17'd9576,17'd25259,17'd25260,17'd24979,17'd25261,17'd7267,17'd10702,17'd9316,17'd25262,17'd25263,17'd25264,17'd25265,17'd16781,17'd16781,17'd25131,17'd15405,17'd13107,17'd23505,17'd25266,17'd9716,17'd25267,17'd25268,17'd16677,17'd25269,17'd25270,17'd25271,17'd24986,17'd22470,17'd11790,17'd25272,17'd24024,17'd25273,17'd25274,17'd25275,17'd13998,17'd25276,17'd25277,17'd25278,17'd18196,17'd9193,17'd9194,17'd16795,17'd11277,17'd11670,17'd11131,17'd10854,17'd21206,17'd21206,17'd14810,17'd13253,17'd12414,17'd12415,17'd15811,17'd25279,17'd12417,17'd12579,17'd23855,17'd24991,17'd24707,17'd24209,17'd24706,17'd25143,17'd22472,17'd22992,17'd23168,17'd24030,17'd24991,17'd23511,17'd24030,17'd21671,17'd15185,17'd13645,17'd12115,17'd13362,17'd11806,17'd11961,17'd13520,17'd19158,17'd11965,17'd25144,17'd11131,17'd11275,17'd11397,17'd11396,17'd25280,17'd21206,17'd10329,17'd16319,17'd25281,17'd16318,17'd9345,17'd25282,17'd19531,17'd21669,17'd17473,17'd10173,17'd9189,17'd16067,17'd8728,17'd19535,17'd17481,17'd8414,17'd19923,17'd8249,17'd20612,17'd25283,17'd25284,17'd25285,17'd25286,17'd16334,17'd19034,17'd16919,17'd25287,17'd25288,17'd24044,17'd17353,17'd11674,17'd23866,17'd17127,17'd25289,17'd25290,17'd18203,17'd15056,17'd9197,17'd25291,17'd16332,17'd10179,17'd10860,17'd8255,17'd8254,17'd15693,17'd18920,17'd25154,17'd25292,17'd9891,17'd25293,17'd25294,17'd25295,17'd17611,17'd25296,17'd16213,17'd19651,17'd25297,17'd25298,17'd25299,17'd25300,17'd25301,17'd25302,17'd25303,17'd25304,17'd25305,17'd25306,17'd25167,17'd24888,17'd25168,17'd25307,17'd24399,17'd24399,17'd24403,17'd25308,17'd25309,17'd25309,17'd25310,17'd25169,17'd24237,17'd24404,17'd24890,17'd24403,17'd25023,17'd25023,17'd25023,17'd24890,17'd24238,17'd24579,17'd25311,17'd25312,17'd25313,17'd25172,17'd24582,17'd24583,17'd24584,17'd23723,17'd25176,17'd25176,17'd25314,17'd25315,17'd24892,17'd25316,17'd25317,17'd25318,17'd25319,17'd25320,17'd23912,17'd24739,17'd25032,17'd25321,17'd25322,17'd25323,17'd25324,17'd24099,17'd25325,17'd25326,17'd25327,17'd25328,17'd25189,17'd25329,17'd25330,17'd25331,17'd25332,17'd25333,17'd25191,17'd25334,17'd25335,17'd25336,17'd25337,17'd25338,17'd24609,17'd25339,17'd25340,17'd25341,17'd25342,17'd25343,17'd25344,17'd21872,17'd25345,17'd25346,17'd25347,17'd25348,17'd25349,17'd25350,17'd21735,17'd25351,17'd25210,17'd25212,17'd25352,17'd25352,17'd25353,17'd25354,17'd25355,17'd19331,17'd19069,17'd19709,17'd19816,17'd18014,17'd25214,17'd25356,17'd18486,17'd25357,17'd25072,17'd25074,17'd25358,17'd17394,17'd17773,17'd19451,17'd24788,17'd25359,17'd21608,17'd25219,17'd24790,17'd24790,17'd22243,17'd22243,17'd25220,17'd25360,17'd12135,17'd22758,17'd24644,17'd24644,17'd22759,17'd7824,17'd23975,17'd7008,17'd5607,17'd4992,17'd5323,17'd4992,17'd5326,17'd5758,17'd5481,17'd5611,17'd5609,17'd5478,17'd5326,17'd4994,17'd5324,17'd5324,17'd4993,17'd4993,17'd5326,17'd25225,17'd5759,17'd5482,17'd5332,17'd6388,17'd5919,17'd25361,17'd24653,17'd13925,17'd14971,17'd17655,17'd15224,17'd21001,17'd16247,17'd17065,17'd17065,17'd16371,17'd18619,17'd18741,17'd20384,17'd19847,17'd19714,17'd21614,17'd25362,17'd20117,17'd25363,17'd19592,17'd25364,17'd25365,17'd25366,17'd15616,17'd25367,17'd14172,17'd25368,17'd25369,17'd25234,17'd25370,17'd25371,17'd25372,17'd25373,17'd954,17'd4084,17'd2576,17'd780,17'd25374,17'd1105,17'd2100,17'd2396,17'd24955,17'd25099,17'd25099,17'd25375,17'd25376,17'd24504,17'd24504,17'd24172,17'd24327,17'd25377,17'd25378,17'd25379,17'd25377,17'd25240,17'd25380,17'd5781,17'd24175,17'd23135,17'd23135,17'd23654,17'd23483,17'd25381,17'd25109,17'd24964,17'd3717,17'd5032,17'd4065,17'd6724,17'd3082,17'd4565,17'd25382,17'd25111,17'd25112,17'd25383,17'd25246,17'd23489,17'd24332,17'd179,17'd17075
},
'{
17'd4892,17'd25384,17'd14070,17'd4247,17'd2423,17'd10260,17'd24,17'd3753,17'd5205,17'd3753,17'd3753,17'd6,17'd6,17'd6,17'd5,17'd24,17'd22,17'd22,17'd21,17'd20,17'd20,17'd20,17'd21,17'd23,17'd23,17'd23,17'd1832,17'd1832,17'd285,17'd27,17'd27,17'd652,17'd653,17'd3908,17'd3433,17'd3433,17'd3256,17'd2940,17'd2601,17'd2264,17'd19874,17'd2431,17'd2607,17'd25385,17'd25386,17'd3919,17'd25387,17'd25388,17'd11894,17'd6606,17'd24678,17'd23494,17'd22621,17'd22795,17'd21176,17'd25389,17'd25390,17'd25391,17'd18766,17'd25392,17'd25393,17'd25394,17'd23836,17'd15764,17'd23324,17'd24344,17'd16027,17'd14470,17'd17096,17'd12813,17'd12527,17'd13092,17'd14469,17'd13092,17'd13092,17'd12955,17'd12218,17'd12530,17'd12680,17'd12957,17'd11764,17'd14472,17'd17941,17'd25395,17'd17206,17'd19384,17'd18776,17'd18777,17'd16768,17'd16768,17'd15902,17'd15524,17'd18060,17'd18060,17'd16289,17'd16880,17'd10565,17'd9703,17'd9703,17'd10113,17'd15006,17'd7750,17'd6140,17'd9009,17'd25396,17'd24978,17'd24979,17'd25397,17'd7925,17'd9316,17'd25398,17'd25399,17'd9993,17'd16180,17'd16045,17'd15915,17'd16295,17'd16418,17'd15787,17'd25400,17'd11367,17'd19769,17'd23158,17'd25401,17'd17957,17'd17115,17'd14917,17'd11938,17'd21202,17'd24695,17'd24986,17'd11945,17'd25402,17'd24532,17'd25403,17'd24023,17'd25404,17'd25405,17'd11510,17'd25406,17'd11664,17'd10476,17'd25407,17'd8872,17'd8873,17'd25408,17'd11135,17'd19532,17'd10854,17'd10990,17'd11131,17'd10854,17'd11522,17'd14261,17'd15434,17'd16913,17'd21504,17'd13515,17'd13517,17'd12579,17'd23855,17'd24537,17'd24208,17'd21505,17'd25143,17'd25143,17'd21362,17'd24209,17'd23512,17'd24859,17'd23511,17'd23855,17'd23168,17'd18198,17'd16326,17'd14671,17'd12115,17'd12996,17'd11961,17'd11961,17'd13520,17'd13516,17'd20910,17'd25144,17'd11131,17'd10854,17'd11397,17'd11396,17'd11398,17'd19280,17'd17719,17'd24037,17'd9343,17'd25281,17'd18324,17'd11809,17'd25409,17'd15566,17'd17232,17'd9743,17'd9194,17'd23860,17'd12264,17'd12865,17'd8414,17'd19923,17'd8248,17'd8103,17'd10480,17'd25410,17'd8254,17'd12427,17'd25289,17'd25411,17'd17127,17'd13648,17'd25412,17'd23864,17'd9196,17'd24862,17'd24545,17'd9887,17'd24713,17'd23173,17'd11405,17'd11405,17'd25148,17'd25412,17'd25413,17'd23519,17'd17482,17'd17609,17'd17609,17'd15435,17'd12265,17'd15693,17'd15193,17'd25414,17'd25415,17'd11969,17'd7958,17'd15307,17'd14818,17'd19540,17'd15064,17'd14941,17'd25416,17'd25417,17'd25418,17'd25419,17'd25420,17'd25421,17'd25422,17'd25423,17'd25306,17'd24573,17'd24573,17'd24888,17'd25168,17'd25424,17'd25022,17'd25022,17'd25425,17'd25426,17'd25427,17'd25427,17'd25426,17'd24578,17'd24890,17'd24238,17'd24890,17'd24403,17'd25023,17'd25023,17'd25428,17'd25023,17'd25023,17'd24238,17'd25429,17'd25311,17'd25313,17'd25430,17'd25172,17'd25431,17'd24583,17'd23909,17'd24892,17'd23723,17'd25432,17'd25433,17'd25434,17'd24737,17'd25435,17'd25436,17'd25437,17'd25438,17'd24079,17'd23912,17'd25320,17'd25439,17'd25440,17'd25441,17'd25442,17'd25443,17'd25444,17'd25445,17'd25446,17'd25447,17'd25448,17'd25449,17'd25450,17'd25451,17'd23061,17'd23235,17'd25191,17'd25042,17'd25452,17'd25453,17'd25447,17'd25454,17'd24763,17'd25455,17'd25456,17'd25457,17'd25458,17'd25454,17'd25459,17'd25460,17'd25461,17'd25462,17'd25463,17'd25464,17'd25465,17'd25466,17'd25467,17'd25468,17'd20961,17'd20653,17'd25469,17'd20495,17'd25354,17'd18610,17'd24633,17'd19452,17'd19709,17'd19817,17'd19710,17'd25470,17'd25471,17'd25472,17'd25357,17'd17392,17'd25473,17'd25474,17'd25475,17'd17771,17'd18734,17'd25476,17'd25477,17'd25478,17'd25479,17'd25480,17'd21451,17'd25481,17'd24640,17'd24640,17'd22243,17'd25482,17'd25360,17'd25483,17'd22758,17'd23279,17'd25484,17'd10196,17'd23458,17'd23799,17'd24944,17'd5607,17'd5323,17'd5325,17'd5478,17'd5481,17'd5331,17'd5158,17'd5611,17'd5609,17'd5610,17'd5478,17'd5151,17'd5324,17'd5325,17'd5325,17'd5326,17'd25225,17'd5759,17'd5758,17'd5482,17'd5332,17'd5919,17'd24652,17'd14048,17'd13558,17'd14970,17'd15094,17'd15225,17'd21453,17'd16121,17'd16371,17'd16371,17'd16371,17'd18619,17'd18498,17'd18742,17'd19847,17'd19714,17'd20849,17'd23465,17'd16251,17'd25485,17'd21456,17'd11713,17'd25486,17'd19351,17'd25487,17'd25488,17'd25489,17'd25490,17'd2881,17'd25491,17'd25492,17'd25493,17'd25494,17'd25495,17'd3100,17'd2775,17'd2576,17'd1383,17'd25374,17'd1105,17'd2100,17'd2396,17'd24955,17'd25239,17'd25239,17'd25496,17'd25376,17'd24327,17'd24327,17'd25101,17'd24503,17'd25377,17'd25378,17'd25379,17'd25241,17'd24172,17'd25497,17'd5781,17'd24175,17'd23135,17'd23135,17'd25106,17'd23654,17'd25242,17'd25498,17'd24964,17'd15486,17'd3398,17'd4065,17'd6724,17'd3082,17'd2755,17'd25382,17'd25111,17'd25244,17'd23138,17'd25499,17'd612,17'd280,17'd179,17'd17075
},
'{
17'd4243,17'd6420,17'd7214,17'd12647,17'd8814,17'd4242,17'd5,17'd6,17'd3753,17'd3753,17'd3753,17'd3753,17'd3753,17'd5,17'd23,17'd23,17'd22,17'd22,17'd21,17'd20,17'd1128,17'd20,17'd21,17'd23,17'd23,17'd284,17'd22,17'd22,17'd20,17'd11,17'd19,17'd288,17'd468,17'd468,17'd3595,17'd3595,17'd4249,17'd3104,17'd2604,17'd2604,17'd2605,17'd2948,17'd3261,17'd25500,17'd25501,17'd25502,17'd4902,17'd6446,17'd7232,17'd24678,17'd25503,17'd23317,17'd22276,17'd25504,17'd25505,17'd25506,17'd25507,17'd25508,17'd25509,17'd18646,17'd25510,17'd24683,17'd25511,17'd16027,17'd24344,17'd24344,17'd23324,17'd15383,17'd13599,17'd13092,17'd12357,17'd12357,17'd13209,17'd12678,17'd13209,17'd15137,17'd12218,17'd12815,17'd12361,17'd11913,17'd12681,17'd17204,17'd25512,17'd19008,17'd19256,17'd16769,17'd16033,17'd16768,17'd16033,17'd16033,17'd17320,17'd16519,17'd16164,17'd16164,17'd16028,17'd16880,17'd10429,17'd10565,17'd10565,17'd9300,17'd7750,17'd5255,17'd9009,17'd25513,17'd7760,17'd25514,17'd8224,17'd7925,17'd7430,17'd7593,17'd9852,17'd25515,17'd15785,17'd25516,17'd9994,17'd9853,17'd25517,17'd25518,17'd25519,17'd25520,17'd25521,17'd25522,17'd9858,17'd10303,17'd18073,17'd17117,17'd13350,17'd16678,17'd22470,17'd24850,17'd24021,17'd24356,17'd11938,17'd15172,17'd12094,17'd21052,17'd13997,17'd11506,17'd11389,17'd25523,17'd24702,17'd17124,17'd9337,17'd25524,17'd25525,17'd15048,17'd12863,17'd12423,17'd11399,17'd10854,17'd10990,17'd13645,17'd14261,17'd16324,17'd16685,17'd12416,17'd13517,17'd13517,17'd12416,17'd16913,17'd18200,17'd18200,17'd16203,17'd22472,17'd23169,17'd24706,17'd24209,17'd25526,17'd25527,17'd25528,17'd16558,17'd12253,17'd11960,17'd12422,17'd13645,17'd11964,17'd12260,17'd12113,17'd11961,17'd11806,17'd19158,17'd11275,17'd10475,17'd16555,17'd24860,17'd10854,17'd14673,17'd16068,17'd19532,17'd9883,17'd9619,17'd18332,17'd9474,17'd25529,17'd19918,17'd25530,17'd15681,17'd15566,17'd17232,17'd15682,17'd25531,17'd23517,17'd25532,17'd24042,17'd11138,17'd25412,17'd17483,17'd25533,17'd17609,17'd17128,17'd13648,17'd10028,17'd12588,17'd9887,17'd24545,17'd8571,17'd8730,17'd8728,17'd8725,17'd8725,17'd8724,17'd8569,17'd16205,17'd16205,17'd16205,17'd8571,17'd8573,17'd8578,17'd8580,17'd17483,17'd17850,17'd14676,17'd16333,17'd13765,17'd23688,17'd12266,17'd20455,17'd19646,17'd25534,17'd25535,17'd15443,17'd25536,17'd8429,17'd25537,17'd15446,17'd25538,17'd25539,17'd25540,17'd25541,17'd25542,17'd25543,17'd25544,17'd25545,17'd25546,17'd24887,17'd25547,17'd25548,17'd24574,17'd24399,17'd25022,17'd24577,17'd25549,17'd25549,17'd25550,17'd25310,17'd25551,17'd25169,17'd25023,17'd25552,17'd25023,17'd24403,17'd24237,17'd25553,17'd25554,17'd25555,17'd25556,17'd25557,17'd25558,17'd25559,17'd25312,17'd25560,17'd25312,17'd25313,17'd25561,17'd25562,17'd24582,17'd24736,17'd23908,17'd24077,17'd25563,17'd25564,17'd23908,17'd25565,17'd25566,17'd25567,17'd24586,17'd24079,17'd25028,17'd25568,17'd25569,17'd25570,17'd25571,17'd25572,17'd25573,17'd25574,17'd21866,17'd25575,17'd25576,17'd25577,17'd25578,17'd25579,17'd25580,17'd24266,17'd25581,17'd25582,17'd25583,17'd25584,17'd25585,17'd25586,17'd25587,17'd25588,17'd25589,17'd25589,17'd25590,17'd25591,17'd25592,17'd25593,17'd25594,17'd25595,17'd25596,17'd25597,17'd25598,17'd25599,17'd25466,17'd22201,17'd21270,17'd25600,17'd25601,17'd25602,17'd25603,17'd25604,17'd25605,17'd24467,17'd19213,17'd25606,17'd19451,17'd25607,17'd25608,17'd25609,17'd25610,17'd25611,17'd25612,17'd25613,17'd20652,17'd21422,17'd19456,17'd25614,17'd25615,17'd25616,17'd19474,17'd25617,17'd25618,17'd25619,17'd25620,17'd25621,17'd24639,17'd25622,17'd25623,17'd22243,17'd25624,17'd25624,17'd22758,17'd25625,17'd23628,17'd8608,17'd25626,17'd5608,17'd5326,17'd5326,17'd5480,17'd5151,17'd5481,17'd5762,17'd25627,17'd5331,17'd5481,17'd5611,17'd5481,17'd5481,17'd5480,17'd5146,17'd4994,17'd24944,17'd25628,17'd25629,17'd5759,17'd5482,17'd5332,17'd6553,17'd6852,17'd25226,17'd24653,17'd13558,17'd14970,17'd14969,17'd15224,17'd16247,17'd16371,17'd16247,17'd16371,17'd16371,17'd18741,17'd18620,17'd18742,17'd19480,17'd20849,17'd24486,17'd25630,17'd25631,17'd25089,17'd25632,17'd25633,17'd15099,17'd16254,17'd18379,17'd25634,17'd25635,17'd25636,17'd25637,17'd25638,17'd25639,17'd25640,17'd25641,17'd1088,17'd2585,17'd598,17'd941,17'd1105,17'd945,17'd2100,17'd2396,17'd24668,17'd25642,17'd25642,17'd25643,17'd25644,17'd24503,17'd25645,17'd24503,17'd25376,17'd25241,17'd25103,17'd25103,17'd25241,17'd25240,17'd24819,17'd25646,17'd24169,17'd23135,17'd23135,17'd7515,17'd25106,17'd23996,17'd25647,17'd5636,17'd6242,17'd3399,17'd5501,17'd6576,17'd4564,17'd6578,17'd25110,17'd5641,17'd25648,17'd20866,17'd22445,17'd964,17'd638,17'd589,17'd280
},
'{
17'd4243,17'd6420,17'd7214,17'd12647,17'd16747,17'd10260,17'd5,17'd6,17'd6,17'd3753,17'd5793,17'd5793,17'd3753,17'd5,17'd23,17'd25,17'd22,17'd21,17'd20,17'd20,17'd1128,17'd11,17'd21,17'd25,17'd23,17'd284,17'd22,17'd21,17'd11,17'd19,17'd1277,17'd1277,17'd468,17'd468,17'd3595,17'd3595,17'd4249,17'd3104,17'd4739,17'd4739,17'd2605,17'd2948,17'd3261,17'd25649,17'd25501,17'd25650,17'd4902,17'd25651,17'd6755,17'd11742,17'd11742,17'd23494,17'd25652,17'd25653,17'd25654,17'd25507,17'd25655,17'd19885,17'd18047,17'd18769,17'd25656,17'd25657,17'd25658,17'd24519,17'd24344,17'd23324,17'd18173,17'd19005,17'd13599,17'd13092,17'd14469,17'd14469,17'd13209,17'd12527,17'd12955,17'd14764,17'd12362,17'd12362,17'd12361,17'd12531,17'd17317,17'd17205,17'd18656,17'd18060,17'd15645,17'd15524,17'd16768,17'd16987,17'd16033,17'd16034,17'd17207,17'd16289,17'd16164,17'd16164,17'd16028,17'd15766,17'd15765,17'd16410,17'd10429,17'd9440,17'd5255,17'd5253,17'd25659,17'd7918,17'd25514,17'd25127,17'd9021,17'd10435,17'd9852,17'd25515,17'd25660,17'd15539,17'd10437,17'd25661,17'd10572,17'd10436,17'd25662,17'd25663,17'd10297,17'd25664,17'd25665,17'd25666,17'd25667,17'd20748,17'd17115,17'd25668,17'd25669,17'd11948,17'd11796,17'd24986,17'd23844,17'd11941,17'd15172,17'd12093,17'd12406,17'd12403,17'd18912,17'd11655,17'd25406,17'd25277,17'd10602,17'd9473,17'd9347,17'd9193,17'd9478,17'd11277,17'd11400,17'd12584,17'd11399,17'd11131,17'd11965,17'd19158,17'd14130,17'd25670,17'd18564,17'd12108,17'd13517,17'd12417,17'd21504,17'd24991,17'd18200,17'd25671,17'd24995,17'd16442,17'd23167,17'd24993,17'd24705,17'd25526,17'd25672,17'd25528,17'd12860,17'd12580,17'd13135,17'd12262,17'd13516,17'd13762,17'd12858,17'd12113,17'd11806,17'd15185,17'd11397,17'd11130,17'd10475,17'd10740,17'd16320,17'd10604,17'd14810,17'd11524,17'd19280,17'd17719,17'd9619,17'd9478,17'd25673,17'd25674,17'd25675,17'd25676,17'd25530,17'd19279,17'd9743,17'd10336,17'd25677,17'd12264,17'd12865,17'd25678,17'd25679,17'd8419,17'd15301,17'd25680,17'd23864,17'd8733,17'd23343,17'd21987,17'd8571,17'd8724,17'd8886,17'd9045,17'd9041,17'd9041,17'd9194,17'd15684,17'd23859,17'd23859,17'd23859,17'd24212,17'd24212,17'd9195,17'd8724,17'd8572,17'd8248,17'd8580,17'd8250,17'd17128,17'd8255,17'd13006,17'd15694,17'd10180,17'd25681,17'd19646,17'd14392,17'd17130,17'd25682,17'd25683,17'd9893,17'd25684,17'd15446,17'd25685,17'd25686,17'd25687,17'd25688,17'd25689,17'd25690,17'd25691,17'd25692,17'd25693,17'd25694,17'd25695,17'd24398,17'd24399,17'd25022,17'd24577,17'd25549,17'd25549,17'd25550,17'd25550,17'd25551,17'd25170,17'd25021,17'd25023,17'd25552,17'd25023,17'd24403,17'd24403,17'd25553,17'd25696,17'd25555,17'd25697,17'd25698,17'd25429,17'd25699,17'd25700,17'd25701,17'd25699,17'd25311,17'd25702,17'd25703,17'd25562,17'd25704,17'd25705,17'd23722,17'd25706,17'd25434,17'd23908,17'd25707,17'd25708,17'd23723,17'd23911,17'd25175,17'd25173,17'd25709,17'd25710,17'd25711,17'd25712,17'd25713,17'd25714,17'd25715,17'd25716,17'd25717,17'd25718,17'd25719,17'd25720,17'd25721,17'd25722,17'd25723,17'd25724,17'd25725,17'd25726,17'd25727,17'd25728,17'd25729,17'd25730,17'd25731,17'd25732,17'd25733,17'd25734,17'd25735,17'd25736,17'd25737,17'd25580,17'd25738,17'd25739,17'd25740,17'd25741,17'd25742,17'd25743,17'd25744,17'd25745,17'd25746,17'd25747,17'd18611,17'd19210,17'd25748,17'd25749,17'd19976,17'd19213,17'd25750,17'd19568,17'd19709,17'd25751,17'd25752,17'd25753,17'd25754,17'd25755,17'd25756,17'd24291,17'd25757,17'd21737,17'd25758,17'd25749,17'd25759,17'd20530,17'd25760,17'd25761,17'd25762,17'd25763,17'd25764,17'd25765,17'd21609,17'd25766,17'd25623,17'd25623,17'd25624,17'd25081,17'd25767,17'd25768,17'd10196,17'd7327,17'd6212,17'd5479,17'd5609,17'd5150,17'd25769,17'd4844,17'd5336,17'd5336,17'd5331,17'd5331,17'd5158,17'd5158,17'd5481,17'd25770,17'd5151,17'd4993,17'd5326,17'd25628,17'd25629,17'd5759,17'd5482,17'd5760,17'd6387,17'd6852,17'd25226,17'd25085,17'd13406,17'd14970,17'd14724,17'd15225,17'd15988,17'd16247,17'd16247,17'd16371,17'd16371,17'd16247,17'd18620,17'd18742,17'd19480,17'd19223,17'd25771,17'd21932,17'd21933,17'd22091,17'd25772,17'd25773,17'd25774,17'd25775,17'd25776,17'd25634,17'd25777,17'd23123,17'd25778,17'd25779,17'd25780,17'd25781,17'd25782,17'd25783,17'd2930,17'd2589,17'd198,17'd1947,17'd944,17'd12645,17'd2396,17'd24668,17'd25642,17'd25643,17'd25784,17'd25785,17'd25376,17'd25645,17'd24503,17'd25376,17'd25241,17'd25103,17'd25103,17'd25241,17'd24504,17'd24817,17'd25786,17'd25787,17'd23309,17'd23135,17'd7515,17'd25106,17'd23996,17'd25647,17'd5780,17'd5945,17'd3227,17'd4407,17'd4718,17'd4564,17'd6578,17'd5369,17'd25788,17'd25789,17'd2926,17'd2416,17'd964,17'd963,17'd590,17'd770
},
'{
17'd4243,17'd6420,17'd7214,17'd12647,17'd16747,17'd10260,17'd23,17'd5,17'd6,17'd3753,17'd5793,17'd5793,17'd3753,17'd5,17'd23,17'd21,17'd20,17'd20,17'd20,17'd11,17'd11,17'd11,17'd21,17'd25,17'd23,17'd22,17'd22,17'd22,17'd20,17'd11,17'd19,17'd16,17'd289,17'd289,17'd3595,17'd3595,17'd4249,17'd4249,17'd4250,17'd25790,17'd2605,17'd4253,17'd3912,17'd25791,17'd25792,17'd5064,17'd11893,17'd7395,17'd6606,17'd11742,17'd11742,17'd25793,17'd22114,17'd25794,17'd25795,17'd25796,17'd25797,17'd19885,17'd25798,17'd25799,17'd25800,17'd25801,17'd24684,17'd24519,17'd23836,17'd21963,17'd25802,17'd19005,17'd13599,17'd13092,17'd14469,17'd16284,17'd12679,17'd12679,17'd14890,17'd12530,17'd12362,17'd12361,17'd12532,17'd12531,17'd17204,17'd19891,17'd18656,17'd16164,17'd16659,17'd16033,17'd16768,17'd16987,17'd17810,17'd17320,17'd17319,17'd16289,17'd16164,17'd16164,17'd15766,17'd15766,17'd15765,17'd11231,17'd10429,17'd13846,17'd5255,17'd5252,17'd25803,17'd25804,17'd25397,17'd7925,17'd9317,17'd25515,17'd15539,17'd25805,17'd25400,17'd13735,17'd10438,17'd10438,17'd10437,17'd14783,17'd25518,17'd25400,17'd25806,17'd21973,17'd22805,17'd25807,17'd25267,17'd17002,17'd16900,17'd13240,17'd25808,17'd11799,17'd25809,17'd25137,17'd25405,17'd11792,17'd24699,17'd13638,17'd12407,17'd18912,17'd11794,17'd16679,17'd25810,17'd10732,17'd25811,17'd11136,17'd9347,17'd12117,17'd15048,17'd11134,17'd10991,17'd13886,17'd10854,17'd11131,17'd10989,17'd11961,17'd12578,17'd15434,17'd12254,17'd12108,17'd13515,17'd12416,17'd23855,17'd18200,17'd16685,17'd22819,17'd22472,17'd22472,17'd22992,17'd24362,17'd24031,17'd24859,17'd24991,17'd18200,17'd12253,17'd11958,17'd16204,17'd12115,17'd11964,17'd11807,17'd12999,17'd12999,17'd11963,17'd13516,17'd22816,17'd22647,17'd10475,17'd10739,17'd10475,17'd24860,17'd14931,17'd14263,17'd24996,17'd17719,17'd17011,17'd15048,17'd9473,17'd15300,17'd25812,17'd15181,17'd16070,17'd11809,17'd9190,17'd15684,17'd8879,17'd8409,17'd8573,17'd8577,17'd21208,17'd25813,17'd8419,17'd25148,17'd8887,17'd21987,17'd11531,17'd12425,17'd25677,17'd9194,17'd10175,17'd8874,17'd10174,17'd13887,17'd15180,17'd17716,17'd25814,17'd25814,17'd17716,17'd24361,17'd10174,17'd9041,17'd8724,17'd8572,17'd9349,17'd19923,17'd19780,17'd8251,17'd8581,17'd16688,17'd16329,17'd16804,17'd19036,17'd10747,17'd7622,17'd14266,17'd25815,17'd15306,17'd7300,17'd18455,17'd8116,17'd25816,17'd25817,17'd25818,17'd25819,17'd25820,17'd25821,17'd25822,17'd25823,17'd25824,17'd24732,17'd25548,17'd24399,17'd24399,17'd24577,17'd25825,17'd25308,17'd25826,17'd25826,17'd25826,17'd25827,17'd25170,17'd25021,17'd25023,17'd25552,17'd25023,17'd24403,17'd24890,17'd25559,17'd25696,17'd25828,17'd25698,17'd25560,17'd25562,17'd23553,17'd24408,17'd25829,17'd25830,17'd25699,17'd25702,17'd25831,17'd25831,17'd25172,17'd25832,17'd24076,17'd24077,17'd23909,17'd24242,17'd25833,17'd25565,17'd24243,17'd25176,17'd25175,17'd25834,17'd25176,17'd25835,17'd25836,17'd25837,17'd25838,17'd25839,17'd21091,17'd25840,17'd25841,17'd25842,17'd25736,17'd25843,17'd25844,17'd25845,17'd24273,17'd25581,17'd25846,17'd25847,17'd25585,17'd25728,17'd25848,17'd25849,17'd25458,17'd25850,17'd25733,17'd25851,17'd25852,17'd25853,17'd25854,17'd24603,17'd25855,17'd25856,17'd25857,17'd25858,17'd25859,17'd25860,17'd25861,17'd25862,17'd25863,17'd18121,17'd18244,17'd19211,17'd25864,17'd25864,17'd19473,17'd19213,17'd25865,17'd19710,17'd19710,17'd25615,17'd25866,17'd24932,17'd25867,17'd25868,17'd25869,17'd25870,17'd21890,17'd20662,17'd20220,17'd25871,17'd25872,17'd25873,17'd25874,17'd25218,17'd25875,17'd25876,17'd24940,17'd24940,17'd21609,17'd25766,17'd25623,17'd25623,17'd25482,17'd25877,17'd24643,17'd25878,17'd22759,17'd8608,17'd25626,17'd6383,17'd5610,17'd5478,17'd4843,17'd4844,17'd5158,17'd6387,17'd6389,17'd6218,17'd5332,17'd5331,17'd5482,17'd5611,17'd5150,17'd4993,17'd4994,17'd5479,17'd25225,17'd25629,17'd5759,17'd5482,17'd6388,17'd6852,17'd12465,17'd25085,17'd13406,17'd13925,17'd14165,17'd14968,17'd15725,17'd15988,17'd16247,17'd16371,17'd16371,17'd16247,17'd18620,17'd18742,17'd19480,17'd20849,17'd25879,17'd21003,17'd25880,17'd22091,17'd25881,17'd25882,17'd25883,17'd25884,17'd25885,17'd25886,17'd25887,17'd25888,17'd25889,17'd25890,17'd25891,17'd25892,17'd25893,17'd25894,17'd9103,17'd2575,17'd941,17'd943,17'd945,17'd12645,17'd2396,17'd24668,17'd25642,17'd25642,17'd25895,17'd25896,17'd25100,17'd25100,17'd24503,17'd25376,17'd25897,17'd24823,17'd24823,17'd24503,17'd25240,17'd24959,17'd24824,17'd23482,17'd6723,17'd6723,17'd24175,17'd23820,17'd23996,17'd25647,17'd5780,17'd15622,17'd3399,17'd5635,17'd7193,17'd3720,17'd25898,17'd25899,17'd25900,17'd25901,17'd3242,17'd2416,17'd181,17'd182,17'd250,17'd15741
},
'{
17'd4892,17'd6420,17'd7214,17'd2590,17'd16747,17'd10260,17'd23,17'd4,17'd6,17'd6,17'd3753,17'd3753,17'd3594,17'd24,17'd21,17'd20,17'd2598,17'd2598,17'd11,17'd11,17'd11,17'd10,17'd21,17'd21,17'd22,17'd22,17'd22,17'd20,17'd11,17'd11,17'd18,17'd16,17'd289,17'd289,17'd3755,17'd3595,17'd4249,17'd4249,17'd5210,17'd25790,17'd25902,17'd4253,17'd3912,17'd4585,17'd25903,17'd5666,17'd11741,17'd9282,17'd6606,17'd7072,17'd6913,17'd22973,17'd25904,17'd25905,17'd25906,17'd4753,17'd25907,17'd18283,17'd25908,17'd25909,17'd25910,17'd25911,17'd25912,17'd24684,17'd21963,17'd18173,17'd19005,17'd17809,17'd13599,17'd13092,17'd16284,17'd12679,17'd12679,17'd14890,17'd12530,17'd12362,17'd12362,17'd12532,17'd12681,17'd17317,17'd16766,17'd19383,17'd17319,17'd19256,17'd15902,17'd16411,17'd16768,17'd16033,17'd17445,17'd17320,17'd16289,17'd16164,17'd16289,17'd16289,17'd15766,17'd15898,17'd15765,17'd10429,17'd9300,17'd5410,17'd6139,17'd8693,17'd25913,17'd25914,17'd9169,17'd10435,17'd9710,17'd16296,17'd22466,17'd25915,17'd25916,17'd10438,17'd23841,17'd9854,17'd10437,17'd25400,17'd25519,17'd12827,17'd9997,17'd25917,17'd25918,17'd9859,17'd25919,17'd17003,17'd16305,17'd25920,17'd13248,17'd11797,17'd25809,17'd11795,17'd11793,17'd25921,17'd24026,17'd12406,17'd12403,17'd11799,17'd25922,17'd25923,17'd25924,17'd10600,17'd20174,17'd10744,17'd9346,17'd9480,17'd14928,17'd11528,17'd14518,17'd13886,17'd10854,17'd11129,17'd11963,17'd14131,17'd13514,17'd15434,17'd12108,17'd19407,17'd14003,17'd23855,17'd18200,17'd25925,17'd25670,17'd25926,17'd20450,17'd20608,17'd21505,17'd24992,17'd24538,17'd24537,17'd25927,17'd23855,17'd17348,17'd12582,17'd17604,17'd12115,17'd13362,17'd11962,17'd20313,17'd11962,17'd11964,17'd11275,17'd22647,17'd14132,17'd11131,17'd10739,17'd10739,17'd24860,17'd14931,17'd19532,17'd10329,17'd17719,17'd12116,17'd12116,17'd18916,17'd25928,17'd15181,17'd17599,17'd18556,17'd10026,17'd16552,17'd8884,17'd8879,17'd8731,17'd8576,17'd21208,17'd10178,17'd14812,17'd21987,17'd9047,17'd8572,17'd8725,17'd8878,17'd16317,17'd10336,17'd8874,17'd10173,17'd11809,17'd11809,17'd11809,17'd11809,17'd11809,17'd11809,17'd16549,17'd11809,17'd22814,17'd10173,17'd9043,17'd8881,17'd8725,17'd8728,17'd8575,17'd9196,17'd10028,17'd11674,17'd8420,17'd17354,17'd15693,17'd25929,17'd14682,17'd25930,17'd11141,17'd17731,17'd24550,17'd25931,17'd25932,17'd8740,17'd25933,17'd25934,17'd25935,17'd25936,17'd25937,17'd25938,17'd25939,17'd25824,17'd25940,17'd25941,17'd25942,17'd24402,17'd24577,17'd25825,17'd25943,17'd25826,17'd25826,17'd25551,17'd25551,17'd25827,17'd25170,17'd24403,17'd25023,17'd25023,17'd25023,17'd25023,17'd25023,17'd25696,17'd25553,17'd25944,17'd25945,17'd25831,17'd24409,17'd23912,17'd25946,17'd23910,17'd25947,17'd25831,17'd25703,17'd25831,17'd25831,17'd25948,17'd24736,17'd24076,17'd24077,17'd24892,17'd24584,17'd25949,17'd25949,17'd24584,17'd23723,17'd25950,17'd25314,17'd23723,17'd25951,17'd25952,17'd25953,17'd25954,17'd25955,17'd25956,17'd25957,17'd25958,17'd25959,17'd25960,17'd25961,17'd25337,17'd25199,17'd25962,17'd25963,17'd25964,17'd25965,17'd25585,17'd24600,17'd25848,17'd25966,17'd25967,17'd25968,17'd25969,17'd25970,17'd25198,17'd25844,17'd25587,17'd25971,17'd25972,17'd25973,17'd25974,17'd25597,17'd24449,17'd25975,17'd25976,17'd25977,17'd25978,17'd18730,17'd25979,17'd25980,17'd18842,17'd25981,17'd18962,17'd19076,17'd25982,17'd25476,17'd18248,17'd25615,17'd25983,17'd25984,17'd25985,17'd24931,17'd25986,17'd25987,17'd23777,17'd20091,17'd23259,17'd25988,17'd25989,17'd25990,17'd25991,17'd25992,17'd25993,17'd25077,17'd24940,17'd24940,17'd24940,17'd24941,17'd25994,17'd25995,17'd25482,17'd25996,17'd25997,17'd25768,17'd25998,17'd25999,17'd6212,17'd23629,17'd5758,17'd5609,17'd5611,17'd4844,17'd5158,17'd6387,17'd6553,17'd6707,17'd6553,17'd5332,17'd5332,17'd5760,17'd4844,17'd5151,17'd5150,17'd5326,17'd25225,17'd5759,17'd5759,17'd5482,17'd6388,17'd6707,17'd12466,17'd14048,17'd13278,17'd13925,17'd13923,17'd14850,17'd15607,17'd15988,17'd16121,17'd16371,17'd16371,17'd16247,17'd18620,17'd18742,17'd19480,17'd18971,17'd20545,17'd25362,17'd23118,17'd19851,17'd26000,17'd26001,17'd26002,17'd26003,17'd15616,17'd26004,17'd20257,17'd24158,17'd2714,17'd26005,17'd26006,17'd26007,17'd26008,17'd26009,17'd7850,17'd2575,17'd941,17'd943,17'd945,17'd2100,17'd2396,17'd24955,17'd25642,17'd25643,17'd25784,17'd26010,17'd25644,17'd25099,17'd25376,17'd25376,17'd25897,17'd24672,17'd24672,17'd24503,17'd25240,17'd24957,17'd26011,17'd26012,17'd24169,17'd6723,17'd24175,17'd23820,17'd23996,17'd24963,17'd5637,17'd17293,17'd3227,17'd4407,17'd4718,17'd4564,17'd6578,17'd5369,17'd5043,17'd25901,17'd3093,17'd2111,17'd17551,17'd181,17'd213,17'd19241
},
'{
17'd4892,17'd4245,17'd1831,17'd2,17'd806,17'd2933,17'd4242,17'd2421,17'd5,17'd5,17'd3594,17'd3594,17'd22268,17'd284,17'd20,17'd1128,17'd20404,17'd20404,17'd1128,17'd1128,17'd11,17'd10,17'd21,17'd21,17'd22,17'd22,17'd22,17'd5518,17'd20,17'd1128,17'd18,17'd18,17'd289,17'd289,17'd4091,17'd3908,17'd5208,17'd4249,17'd5210,17'd5658,17'd4894,17'd4896,17'd5217,17'd26013,17'd26014,17'd12040,17'd26015,17'd6754,17'd11613,17'd7072,17'd8054,17'd26016,17'd12935,17'd25905,17'd4752,17'd26017,17'd4107,17'd18159,17'd26018,17'd26019,17'd26020,17'd26021,17'd25801,17'd25658,17'd21963,17'd18173,17'd19005,17'd13599,17'd13092,17'd13092,17'd12679,17'd12679,17'd12679,17'd12814,17'd12530,17'd12362,17'd12680,17'd12532,17'd12681,17'd17204,17'd18174,17'd18656,17'd16289,17'd17319,17'd24520,17'd16411,17'd15902,17'd16411,17'd17320,17'd16519,17'd21650,17'd21650,17'd16289,17'd16289,17'd15766,17'd15898,17'd15517,17'd10429,17'd8538,17'd5836,17'd6138,17'd26022,17'd7920,17'd26023,17'd9316,17'd9710,17'd9853,17'd9712,17'd25661,17'd25916,17'd12827,17'd23841,17'd9996,17'd11485,17'd13734,17'd26024,17'd13735,17'd26025,17'd26026,17'd26027,17'd26028,17'd26029,17'd24984,17'd16677,17'd13870,17'd25402,17'd19275,17'd11796,17'd25809,17'd11949,17'd26030,17'd25921,17'd25270,17'd12098,17'd12246,17'd24534,17'd26031,17'd26032,17'd26033,17'd26034,17'd10857,17'd23679,17'd10334,17'd18556,17'd11135,17'd10478,17'd10605,17'd10990,17'd11129,17'd11964,17'd11960,17'd12578,17'd12997,17'd12418,17'd13515,17'd13515,17'd12255,17'd18200,17'd18200,17'd25925,17'd24209,17'd26035,17'd20608,17'd21363,17'd22819,17'd23512,17'd24537,17'd25927,17'd26036,17'd16324,17'd15053,17'd12422,17'd12115,17'd12262,17'd12996,17'd13135,17'd12861,17'd11963,17'd10989,17'd11131,17'd14263,17'd11669,17'd11399,17'd11524,17'd14810,17'd14931,17'd16320,17'd16555,17'd10166,17'd9883,17'd11671,17'd21503,17'd10165,17'd17715,17'd26037,17'd11276,17'd10025,17'd9743,17'd17480,17'd8879,17'd8724,17'd8731,17'd21987,17'd10339,17'd12586,17'd8571,17'd16205,17'd8729,17'd15297,17'd24999,17'd16553,17'd24361,17'd9345,17'd10742,17'd11277,17'd16070,17'd11277,17'd17839,17'd17839,17'd11277,17'd11277,17'd12116,17'd12116,17'd12116,17'd10742,17'd9346,17'd8874,17'd15684,17'd26038,17'd26039,17'd9047,17'd9196,17'd23343,17'd13374,17'd11674,17'd16690,17'd12265,17'd15694,17'd7955,17'd26040,17'd14391,17'd10748,17'd15444,17'd26041,17'd26042,17'd26043,17'd26044,17'd26045,17'd26046,17'd26047,17'd26048,17'd26049,17'd26050,17'd26051,17'd25941,17'd26052,17'd26053,17'd25169,17'd25170,17'd25826,17'd25551,17'd26054,17'd25551,17'd25551,17'd25827,17'd25169,17'd25554,17'd25698,17'd25554,17'd25554,17'd25554,17'd25696,17'd25560,17'd26055,17'd25311,17'd25562,17'd26056,17'd25028,17'd26057,17'd26058,17'd26059,17'd26060,17'd26061,17'd25703,17'd25703,17'd25703,17'd25702,17'd25431,17'd23908,17'd24584,17'd23909,17'd23909,17'd26062,17'd26062,17'd23909,17'd24078,17'd25432,17'd26063,17'd24737,17'd26064,17'd26065,17'd26066,17'd26067,17'd26068,17'd26069,17'd26070,17'd26071,17'd26072,17'd26073,17'd26074,17'd26075,17'd25454,17'd26076,17'd26077,17'd26078,17'd26079,17'd26080,17'd24600,17'd25848,17'd25966,17'd26081,17'd25731,17'd26082,17'd25733,17'd26083,17'd26084,17'd26085,17'd26086,17'd26087,17'd25855,17'd26088,17'd25740,17'd26089,17'd26090,17'd20957,17'd26091,17'd26092,17'd18730,17'd25979,17'd26093,17'd18962,17'd18842,17'd18962,17'd18962,17'd19212,17'd19213,17'd26094,17'd24786,17'd26095,17'd26096,17'd26097,17'd26098,17'd26099,17'd26100,17'd26101,17'd26102,17'd19965,17'd26103,17'd26104,17'd26105,17'd26106,17'd26107,17'd26108,17'd26109,17'd24789,17'd24789,17'd26110,17'd24940,17'd25994,17'd25994,17'd22083,17'd25482,17'd25221,17'd26111,17'd22935,17'd25998,17'd7008,17'd23629,17'd24799,17'd5610,17'd5481,17'd5481,17'd5158,17'd5332,17'd6707,17'd9090,17'd9090,17'd6553,17'd6553,17'd6387,17'd5482,17'd5151,17'd5150,17'd5478,17'd5610,17'd5759,17'd5759,17'd5482,17'd5332,17'd6706,17'd10237,17'd25226,17'd13045,17'd14047,17'd14970,17'd15340,17'd15607,17'd15988,17'd15988,17'd16247,17'd18498,17'd18741,17'd18620,17'd18260,17'd19480,17'd26112,17'd26113,17'd23465,17'd19850,17'd23288,17'd26114,17'd19852,17'd26115,17'd25231,17'd15616,17'd18748,17'd26116,17'd23122,17'd26117,17'd26118,17'd26119,17'd26120,17'd26121,17'd26122,17'd799,17'd2905,17'd421,17'd417,17'd1949,17'd2100,17'd2395,17'd24955,17'd25642,17'd25642,17'd25895,17'd25896,17'd25099,17'd25099,17'd25376,17'd25376,17'd25376,17'd25376,17'd24503,17'd24503,17'd24816,17'd24501,17'd26123,17'd26124,17'd23482,17'd23482,17'd24963,17'd23996,17'd23996,17'd24963,17'd5637,17'd15738,17'd3400,17'd5635,17'd7193,17'd3720,17'd25898,17'd25899,17'd26125,17'd20568,17'd3093,17'd2416,17'd805,17'd181,17'd180,17'd26126
},
'{
17'd4243,17'd6420,17'd1831,17'd2,17'd806,17'd2933,17'd4242,17'd4242,17'd23,17'd5,17'd5,17'd5,17'd24,17'd5518,17'd1128,17'd20404,17'd20404,17'd26127,17'd20404,17'd20404,17'd1128,17'd11,17'd21,17'd21,17'd22,17'd22,17'd22,17'd20,17'd11,17'd1128,17'd18,17'd3905,17'd289,17'd289,17'd4091,17'd4091,17'd5208,17'd5208,17'd5379,17'd5806,17'd4742,17'd5380,17'd4744,17'd26013,17'd6116,17'd26128,17'd26015,17'd6754,17'd11613,17'd7072,17'd8054,17'd26129,17'd26130,17'd26131,17'd21336,17'd26132,17'd26133,17'd19743,17'd26134,17'd26135,17'd26020,17'd26021,17'd25911,17'd24840,17'd23324,17'd18173,17'd17809,17'd12954,17'd13092,17'd12679,17'd12679,17'd11626,17'd12065,17'd12530,17'd12361,17'd20424,17'd12531,17'd17317,17'd17204,17'd16766,17'd18656,17'd16289,17'd16289,17'd17445,17'd24520,17'd16033,17'd15902,17'd16033,17'd16519,17'd18060,17'd21185,17'd21650,17'd16164,17'd16164,17'd15898,17'd15898,17'd10429,17'd9300,17'd4767,17'd6138,17'd26022,17'd7918,17'd25514,17'd9169,17'd9852,17'd9853,17'd10436,17'd9592,17'd9854,17'd12827,17'd10820,17'd12687,17'd26136,17'd13223,17'd13856,17'd10438,17'd23841,17'd26137,17'd23673,17'd9858,17'd26138,17'd26139,17'd16675,17'd14917,17'd26140,17'd16903,17'd11659,17'd11658,17'd26141,17'd26142,17'd26143,17'd11940,17'd26144,17'd11944,17'd12851,17'd26145,17'd26146,17'd26147,17'd26148,17'd17011,17'd9346,17'd9620,17'd18556,17'd16561,17'd11400,17'd13886,17'd24860,17'd10853,17'd13516,17'd11806,17'd12414,17'd15434,17'd12859,17'd12417,17'd13515,17'd25279,17'd24991,17'd24856,17'd24707,17'd26149,17'd26150,17'd26151,17'd25926,17'd24209,17'd23512,17'd24030,17'd24856,17'd26036,17'd24207,17'd21505,17'd18443,17'd18444,17'd13516,17'd13362,17'd12858,17'd12858,17'd11962,17'd14262,17'd10990,17'd16555,17'd19282,17'd11132,17'd11524,17'd17236,17'd12720,17'd10990,17'd10475,17'd11133,17'd10741,17'd9883,17'd10331,17'd26152,17'd15052,17'd13886,17'd10478,17'd9884,17'd9480,17'd26153,17'd8884,17'd9195,17'd12425,17'd15429,17'd11811,17'd11967,17'd24368,17'd26154,17'd26154,17'd8885,17'd15944,17'd15187,17'd16549,17'd17011,17'd12116,17'd10479,17'd12863,17'd11670,17'd11670,17'd12863,17'd11527,17'd11527,17'd12863,17'd10330,17'd10329,17'd9884,17'd9741,17'd10742,17'd15569,17'd24361,17'd16067,17'd8569,17'd8731,17'd24711,17'd26155,17'd23173,17'd13373,17'd17240,17'd17127,17'd16333,17'd15693,17'd21508,17'd26156,17'd26157,17'd13259,17'd24217,17'd26158,17'd26159,17'd26160,17'd26161,17'd26162,17'd26163,17'd26164,17'd26165,17'd26166,17'd24887,17'd24732,17'd24401,17'd25021,17'd25169,17'd25826,17'd25551,17'd26054,17'd26054,17'd25551,17'd25551,17'd25170,17'd24578,17'd25698,17'd25698,17'd25554,17'd25558,17'd25554,17'd25554,17'd26167,17'd25311,17'd25948,17'd26168,17'd23556,17'd26169,17'd26170,17'd26171,17'd26169,17'd26172,17'd25947,17'd25829,17'd25703,17'd25561,17'd25702,17'd25561,17'd24583,17'd23553,17'd24584,17'd24891,17'd26062,17'd25949,17'd24891,17'd23909,17'd25433,17'd26173,17'd24737,17'd26174,17'd26175,17'd26176,17'd25953,17'd26177,17'd26178,17'd26179,17'd26180,17'd26181,17'd26073,17'd26182,17'd26183,17'd26184,17'd25199,17'd26185,17'd26186,17'd26187,17'd26188,17'd26189,17'd26190,17'd26191,17'd26192,17'd25342,17'd26082,17'd26193,17'd25590,17'd26194,17'd26195,17'd26196,17'd25050,17'd24273,17'd24267,17'd26197,17'd26198,17'd26199,17'd26200,17'd18234,17'd26201,17'd18122,17'd26202,17'd25980,17'd18962,17'd18842,17'd19473,17'd19473,17'd18962,17'd18734,17'd26094,17'd19330,17'd26203,17'd26204,17'd26205,17'd26206,17'd26207,17'd26208,17'd26209,17'd26210,17'd20817,17'd20366,17'd21289,17'd22728,17'd26211,17'd26212,17'd26213,17'd26214,17'd25993,17'd25077,17'd26110,17'd24940,17'd21452,17'd25994,17'd21766,17'd22083,17'd22413,17'd12443,17'd26215,17'd26216,17'd26217,17'd6212,17'd24799,17'd5759,17'd5482,17'd5760,17'd5331,17'd26218,17'd8154,17'd9394,17'd26219,17'd9090,17'd9090,17'd6852,17'd6388,17'd25770,17'd25770,17'd5478,17'd5610,17'd24799,17'd5759,17'd5758,17'd5760,17'd6706,17'd6852,17'd12466,17'd12306,17'd13165,17'd13558,17'd17655,17'd15606,17'd15988,17'd15725,17'd16121,17'd18741,17'd18741,17'd18620,17'd18260,17'd19480,17'd18375,17'd19848,17'd24486,17'd25630,17'd23981,17'd20699,17'd19852,17'd26220,17'd19351,17'd26221,17'd15100,17'd15732,17'd19723,17'd26222,17'd26223,17'd26224,17'd26225,17'd26226,17'd26227,17'd1115,17'd4084,17'd2589,17'd417,17'd1950,17'd26228,17'd2561,17'd24955,17'd25642,17'd25642,17'd25895,17'd26010,17'd25896,17'd25239,17'd26229,17'd26229,17'd26229,17'd25376,17'd24503,17'd24327,17'd24816,17'd26230,17'd26231,17'd26124,17'd23482,17'd23134,17'd25647,17'd24175,17'd24175,17'd24963,17'd26232,17'd17293,17'd3228,17'd4065,17'd7193,17'd3082,17'd6578,17'd26233,17'd26234,17'd20568,17'd20865,17'd2111,17'd404,17'd182,17'd182,17'd401
},
'{
17'd4891,17'd25384,17'd10535,17'd466,17'd2423,17'd8814,17'd2933,17'd4242,17'd23,17'd24,17'd24,17'd24,17'd284,17'd5517,17'd16636,17'd3430,17'd4089,17'd4089,17'd4089,17'd4089,17'd1128,17'd11,17'd21,17'd21,17'd21,17'd21,17'd20,17'd20,17'd980,17'd980,17'd653,17'd653,17'd289,17'd289,17'd4091,17'd4091,17'd5208,17'd5655,17'd5211,17'd5211,17'd4741,17'd5215,17'd26235,17'd26236,17'd5665,17'd26237,17'd26238,17'd26239,17'd11613,17'd7565,17'd23494,17'd26240,17'd26130,17'd26241,17'd3610,17'd26242,17'd26133,17'd19743,17'd26243,17'd26244,17'd26020,17'd26245,17'd26245,17'd24840,17'd21963,17'd19005,17'd13599,17'd12954,17'd12527,17'd12679,17'd12955,17'd12065,17'd12360,17'd11478,17'd11913,17'd10815,17'd11362,17'd17317,17'd17204,17'd18174,17'd18656,17'd16289,17'd17207,17'd16169,17'd16169,17'd16169,17'd17690,17'd17320,17'd21185,17'd21185,17'd21185,17'd21185,17'd16410,17'd16410,17'd10429,17'd10429,17'd9703,17'd7582,17'd5253,17'd6138,17'd25803,17'd25804,17'd25397,17'd10702,17'd9710,17'd26246,17'd15786,17'd10437,17'd25661,17'd12827,17'd10820,17'd10820,17'd14232,17'd14232,17'd9854,17'd23841,17'd26247,17'd26248,17'd26249,17'd26250,17'd26251,17'd17336,17'd26252,17'd26253,17'd26254,17'd13998,17'd11512,17'd19152,17'd11795,17'd17713,17'd26255,17'd12712,17'd25275,17'd26256,17'd11794,17'd26257,17'd24701,17'd17009,17'd18325,17'd13887,17'd9346,17'd9479,17'd16561,17'd19278,17'd12584,17'd11524,17'd10604,17'd10737,17'd13362,17'd12419,17'd15434,17'd12997,17'd13643,17'd14526,17'd13515,17'd19534,17'd25528,17'd24856,17'd24030,17'd24209,17'd26258,17'd26150,17'd23170,17'd23512,17'd12255,17'd24991,17'd25528,17'd25925,17'd16203,17'd21361,17'd16326,17'd11964,17'd11964,17'd11963,17'd12113,17'd13135,17'd13762,17'd11274,17'd10475,17'd10472,17'd10326,17'd11132,17'd17236,17'd11523,17'd11523,17'd11524,17'd19282,17'd10326,17'd10164,17'd10165,17'd11526,17'd15176,17'd14803,17'd10476,17'd11670,17'd9885,17'd9345,17'd10336,17'd8879,17'd16205,17'd8571,17'd11404,17'd9744,17'd24368,17'd9195,17'd17607,17'd16440,17'd16552,17'd16549,17'd9619,17'd11277,17'd11134,17'd11670,17'd10991,17'd11132,17'd16555,17'd10475,17'd10739,17'd10739,17'd14518,17'd10991,17'd10326,17'd10326,17'd10330,17'd9739,17'd17011,17'd15187,17'd15944,17'd9041,17'd8886,17'd26259,17'd24368,17'd26260,17'd24545,17'd26261,17'd25148,17'd26262,17'd11406,17'd15056,17'd16334,17'd26263,17'd26264,17'd26265,17'd26266,17'd26267,17'd26268,17'd26269,17'd26270,17'd26271,17'd26272,17'd26273,17'd26274,17'd26275,17'd25547,17'd25168,17'd24400,17'd25021,17'd25170,17'd25826,17'd25551,17'd26054,17'd26054,17'd26276,17'd26277,17'd26278,17'd25555,17'd25944,17'd25698,17'd25558,17'd25558,17'd25558,17'd25558,17'd26279,17'd25312,17'd25948,17'd23553,17'd24245,17'd26280,17'd26281,17'd26282,17'd26283,17'd26284,17'd23554,17'd26285,17'd25831,17'd25948,17'd25699,17'd25561,17'd25431,17'd26285,17'd24583,17'd24891,17'd23908,17'd24583,17'd24076,17'd23552,17'd23551,17'd26286,17'd25564,17'd25949,17'd26287,17'd26288,17'd26289,17'd26290,17'd26291,17'd26292,17'd26293,17'd26294,17'd26295,17'd26296,17'd26074,17'd26297,17'd25454,17'd26298,17'd26299,17'd26300,17'd25452,17'd26301,17'd26302,17'd26303,17'd26304,17'd25853,17'd25195,17'd25052,17'd26305,17'd26306,17'd25576,17'd26085,17'd26298,17'd25962,17'd26307,17'd26308,17'd20072,17'd26309,17'd19055,17'd26310,17'd26311,17'd19197,17'd18243,17'd18487,17'd18842,17'd18842,17'd18962,17'd18962,17'd18962,17'd18734,17'd26094,17'd19330,17'd26312,17'd26313,17'd26314,17'd26315,17'd26316,17'd26317,17'd26318,17'd26319,17'd26320,17'd20509,17'd26321,17'd26322,17'd22384,17'd26323,17'd26324,17'd26325,17'd20840,17'd25077,17'd26110,17'd24940,17'd21924,17'd25994,17'd21610,17'd22083,17'd26326,17'd11830,17'd26327,17'd8912,17'd7007,17'd6547,17'd5759,17'd26328,17'd5760,17'd5332,17'd5332,17'd5331,17'd6707,17'd9090,17'd10777,17'd26219,17'd9394,17'd10237,17'd6707,17'd5612,17'd25770,17'd4843,17'd5610,17'd24799,17'd24799,17'd5758,17'd5482,17'd6706,17'd6852,17'd12466,17'd14048,17'd25085,17'd13278,17'd14971,17'd14968,17'd21309,17'd15607,17'd15988,17'd18741,17'd18741,17'd18620,17'd18260,17'd19847,17'd20115,17'd26329,17'd24486,17'd23117,17'd24153,17'd20699,17'd25881,17'd25486,17'd26330,17'd26221,17'd14431,17'd26331,17'd20120,17'd26332,17'd26333,17'd26334,17'd26335,17'd26336,17'd26337,17'd26338,17'd1380,17'd602,17'd1672,17'd1950,17'd2101,17'd2395,17'd24955,17'd24668,17'd25642,17'd25895,17'd25895,17'd26339,17'd26339,17'd25644,17'd25644,17'd25644,17'd25644,17'd25376,17'd24327,17'd24816,17'd24670,17'd26123,17'd26124,17'd23482,17'd23134,17'd25647,17'd24963,17'd26340,17'd25105,17'd26232,17'd15738,17'd3400,17'd4065,17'd6243,17'd4069,17'd26233,17'd26233,17'd26234,17'd26341,17'd26342,17'd26343,17'd594,17'd639,17'd181,17'd1548
},
'{
17'd4425,17'd4243,17'd3252,17'd2595,17'd16636,17'd8814,17'd2933,17'd2591,17'd21,17'd23,17'd23,17'd22,17'd5518,17'd2598,17'd3430,17'd8971,17'd4089,17'd26344,17'd26344,17'd4089,17'd20404,17'd11,17'd21,17'd21,17'd21,17'd21,17'd20,17'd20,17'd980,17'd980,17'd653,17'd653,17'd289,17'd289,17'd4091,17'd4091,17'd3910,17'd5655,17'd5211,17'd5211,17'd4741,17'd5214,17'd5059,17'd26236,17'd5063,17'd26237,17'd26238,17'd26345,17'd26346,17'd26347,17'd25793,17'd26348,17'd26349,17'd21798,17'd15369,17'd21480,17'd26133,17'd26350,17'd26351,17'd26352,17'd26020,17'd26245,17'd26245,17'd26353,17'd21036,17'd19005,17'd12954,17'd12954,17'd12679,17'd12955,17'd12065,17'd12218,17'd11478,17'd11361,17'd10815,17'd17317,17'd17941,17'd19754,17'd19754,17'd18656,17'd16289,17'd18060,17'd16034,17'd16169,17'd16034,17'd24520,17'd22980,17'd16519,17'd21185,17'd21185,17'd21185,17'd21185,17'd16410,17'd10429,17'd10429,17'd9703,17'd9007,17'd5090,17'd6138,17'd8693,17'd26354,17'd25514,17'd13222,17'd12824,17'd15915,17'd15785,17'd15786,17'd26024,17'd10438,17'd12827,17'd23841,17'd9713,17'd11923,17'd11770,17'd11634,17'd11098,17'd26355,17'd26356,17'd26357,17'd26358,17'd26359,17'd26360,17'd26361,17'd26362,17'd11949,17'd26363,17'd26364,17'd19152,17'd11949,17'd26254,17'd25402,17'd12572,17'd26365,17'd26366,17'd26367,17'd10464,17'd26368,17'd10476,17'd9478,17'd9193,17'd10174,17'd11809,17'd9884,17'd26369,17'd11398,17'd11275,17'd20910,17'd15810,17'd12113,17'd12109,17'd12415,17'd16559,17'd13643,17'd14526,17'd14003,17'd24991,17'd26370,17'd26371,17'd24031,17'd26372,17'd26258,17'd26150,17'd24705,17'd23856,17'd23511,17'd26373,17'd25528,17'd24707,17'd24362,17'd18443,17'd11397,17'd11396,17'd13762,17'd11667,17'd11806,17'd12996,17'd11964,17'd10990,17'd10474,17'd26374,17'd10326,17'd11132,17'd17236,17'd13254,17'd11398,17'd11524,17'd19532,17'd10166,17'd17720,17'd10166,17'd17966,17'd15427,17'd10605,17'd21205,17'd10024,17'd9742,17'd10173,17'd9041,17'd8886,17'd12425,17'd8572,17'd8412,17'd24368,17'd9195,17'd17607,17'd9042,17'd16552,17'd19279,17'd9739,17'd9883,17'd11670,17'd10476,17'd10476,17'd11399,17'd10990,17'd14810,17'd10854,17'd10854,17'd10854,17'd10475,17'd19282,17'd19532,17'd19282,17'd19282,17'd20756,17'd9740,17'd9341,17'd9346,17'd8874,17'd15684,17'd16317,17'd8570,17'd26375,17'd26376,17'd26377,17'd26378,17'd26379,17'd26380,17'd25289,17'd26381,17'd26382,17'd26383,17'd26384,17'd26385,17'd26386,17'd26387,17'd26388,17'd26389,17'd26390,17'd26391,17'd26392,17'd26051,17'd26393,17'd25547,17'd25022,17'd25022,17'd25169,17'd25170,17'd25551,17'd25551,17'd26054,17'd26054,17'd26276,17'd26277,17'd26278,17'd25828,17'd26394,17'd25698,17'd25558,17'd25558,17'd25558,17'd25558,17'd26279,17'd25311,17'd25948,17'd23723,17'd23728,17'd26395,17'd26396,17'd26397,17'd26398,17'd26399,17'd24078,17'd24736,17'd25702,17'd25948,17'd26400,17'd25313,17'd25172,17'd25431,17'd24582,17'd24736,17'd24736,17'd24582,17'd23721,17'd24076,17'd25706,17'd25706,17'd26401,17'd25705,17'd25833,17'd26402,17'd26403,17'd26404,17'd26405,17'd26406,17'd26407,17'd26408,17'd26295,17'd26409,17'd26410,17'd26183,17'd25718,17'd26411,17'd26077,17'd26186,17'd25335,17'd26412,17'd26413,17'd26414,17'd25966,17'd26415,17'd25195,17'd26416,17'd26417,17'd26418,17'd25718,17'd26419,17'd26420,17'd25845,17'd23942,17'd26421,17'd26422,17'd26423,17'd26424,17'd26425,17'd26091,17'd26426,17'd18242,17'd26427,17'd25981,17'd19955,17'd24786,17'd24786,17'd19567,17'd19069,17'd26428,17'd26429,17'd26430,17'd26431,17'd26432,17'd26433,17'd26434,17'd26435,17'd26436,17'd26437,17'd26438,17'd26439,17'd26440,17'd20828,17'd26441,17'd26442,17'd26443,17'd26444,17'd26445,17'd25359,17'd25479,17'd21451,17'd25765,17'd21924,17'd26446,17'd21610,17'd26447,17'd11830,17'd26327,17'd26448,17'd26449,17'd6546,17'd5913,17'd26450,17'd26451,17'd5331,17'd5332,17'd6389,17'd8303,17'd8154,17'd10777,17'd10641,17'd26219,17'd26219,17'd9090,17'd26218,17'd26452,17'd4843,17'd5481,17'd24799,17'd24799,17'd5758,17'd5482,17'd6387,17'd6707,17'd26219,17'd25226,17'd14048,17'd13407,17'd13925,17'd14969,17'd15224,17'd15607,17'd15988,17'd18134,17'd18134,17'd18620,17'd18260,17'd19847,17'd18375,17'd19481,17'd19715,17'd20116,17'd26453,17'd26454,17'd21456,17'd26455,17'd20119,17'd26456,17'd22598,17'd26457,17'd20855,17'd26458,17'd26459,17'd26460,17'd26461,17'd26462,17'd26463,17'd26464,17'd2578,17'd24323,17'd194,17'd1672,17'd26228,17'd2243,17'd26465,17'd24668,17'd25642,17'd25895,17'd25895,17'd26339,17'd26339,17'd25644,17'd25644,17'd25644,17'd25644,17'd25376,17'd24327,17'd24816,17'd24816,17'd26011,17'd26124,17'd23482,17'd23134,17'd5636,17'd24963,17'd24330,17'd25105,17'd26232,17'd16257,17'd3228,17'd4065,17'd6243,17'd3082,17'd6252,17'd21162,17'd26234,17'd21945,17'd26466,17'd26467,17'd594,17'd405,17'd181,17'd402
},
'{
17'd4891,17'd4892,17'd3252,17'd1127,17'd3,17'd1275,17'd1275,17'd2933,17'd2933,17'd10260,17'd10260,17'd10260,17'd16747,17'd16636,17'd466,17'd2595,17'd2595,17'd2595,17'd8971,17'd3430,17'd1128,17'd11,17'd21,17'd21,17'd10,17'd11,17'd27,17'd980,17'd980,17'd980,17'd980,17'd1278,17'd652,17'd652,17'd4431,17'd5207,17'd26468,17'd5803,17'd12931,17'd26469,17'd4895,17'd26470,17'd26471,17'd6603,17'd26472,17'd26237,17'd26473,17'd11457,17'd26346,17'd26347,17'd26474,17'd26475,17'd26476,17'd13192,17'd3928,17'd26477,17'd26478,17'd26479,17'd15125,17'd24516,17'd26480,17'd26481,17'd26481,17'd23151,17'd18410,17'd19005,17'd13599,17'd13210,17'd12955,17'd12955,17'd12814,17'd12530,17'd11913,17'd11629,17'd17317,17'd16518,17'd19754,17'd19754,17'd17205,17'd17572,17'd19256,17'd16519,17'd16034,17'd24520,17'd16169,17'd16034,17'd17319,17'd16289,17'd21650,17'd21185,17'd21185,17'd21650,17'd16410,17'd10429,17'd10428,17'd10694,17'd7582,17'd5090,17'd6138,17'd8220,17'd7263,17'd26482,17'd9168,17'd7764,17'd16295,17'd26483,17'd25400,17'd13735,17'd10438,17'd9854,17'd10132,17'd11485,17'd11770,17'd26484,17'd26485,17'd26486,17'd10576,17'd24018,17'd25401,17'd26487,17'd16675,17'd26488,17'd15416,17'd26489,17'd13249,17'd14515,17'd26364,17'd19529,17'd16547,17'd26490,17'd11789,17'd12403,17'd11944,17'd13755,17'd10971,17'd26491,17'd25278,17'd11400,17'd9345,17'd9038,17'd25525,17'd19279,17'd10330,17'd11132,17'd25280,17'd11274,17'd10736,17'd15186,17'd12252,17'd26492,17'd14672,17'd21207,17'd15942,17'd14809,17'd12860,17'd18084,17'd25927,17'd26493,17'd26494,17'd26151,17'd26495,17'd26496,17'd24031,17'd24537,17'd25528,17'd17846,17'd18200,17'd14807,17'd15053,17'd18444,17'd11397,17'd14673,17'd13762,17'd11962,17'd12113,17'd11963,17'd11274,17'd24996,17'd10166,17'd10164,17'd11133,17'd13886,17'd17236,17'd11398,17'd11668,17'd11669,17'd19282,17'd11133,17'd10326,17'd11133,17'd17236,17'd26497,17'd20610,17'd12863,17'd12116,17'd9620,17'd8874,17'd16067,17'd8569,17'd8728,17'd8410,17'd8724,17'd25677,17'd15684,17'd10335,17'd9479,17'd15566,17'd11671,17'd10165,17'd10475,17'd16320,17'd14931,17'd14810,17'd16068,17'd16068,17'd16068,17'd11274,17'd10990,17'd10990,17'd14931,17'd11524,17'd11669,17'd11669,17'd11132,17'd10023,17'd10856,17'd10742,17'd15187,17'd24361,17'd17480,17'd26498,17'd24212,17'd26499,17'd26500,17'd26501,17'd26502,17'd26503,17'd26504,17'd26505,17'd26506,17'd26507,17'd26508,17'd26509,17'd26510,17'd26511,17'd26512,17'd26513,17'd26514,17'd26515,17'd26516,17'd26517,17'd26518,17'd26519,17'd26520,17'd24577,17'd26521,17'd25308,17'd25826,17'd25551,17'd25551,17'd26522,17'd26522,17'd26276,17'd26277,17'd26523,17'd25557,17'd25698,17'd25558,17'd25554,17'd26524,17'd26525,17'd25944,17'd26394,17'd26279,17'd25699,17'd24243,17'd24412,17'd26526,17'd26527,17'd23210,17'd26528,17'd23727,17'd23723,17'd23908,17'd25562,17'd25948,17'd25312,17'd26400,17'd25312,17'd25561,17'd25431,17'd25431,17'd24582,17'd24582,17'd24240,17'd26529,17'd23552,17'd23552,17'd24737,17'd24737,17'd26530,17'd26287,17'd26531,17'd26532,17'd26533,17'd26534,17'd26535,17'd26536,17'd26537,17'd26538,17'd26539,17'd26540,17'd26541,17'd26542,17'd26543,17'd26544,17'd26545,17'd25191,17'd25189,17'd26546,17'd25849,17'd26547,17'd26548,17'd26549,17'd26550,17'd26551,17'd26552,17'd26553,17'd25736,17'd25735,17'd26554,17'd26555,17'd22886,17'd20074,17'd26556,17'd26557,17'd26558,17'd26559,17'd19679,17'd26427,17'd26560,17'd25615,17'd26561,17'd19330,17'd19330,17'd26562,17'd26563,17'd26564,17'd26565,17'd22551,17'd26566,17'd26567,17'd26568,17'd26569,17'd26570,17'd26571,17'd26572,17'd26573,17'd20969,17'd26574,17'd26575,17'd26576,17'd26577,17'd26578,17'd26579,17'd26580,17'd21922,17'd24940,17'd21301,17'd25481,17'd21452,17'd26581,17'd26582,17'd26326,17'd26583,17'd26584,17'd8912,17'd6545,17'd6211,17'd6384,17'd24800,17'd26451,17'd6388,17'd6388,17'd6389,17'd8303,17'd10777,17'd11576,17'd10641,17'd12466,17'd9394,17'd6218,17'd5158,17'd5611,17'd5481,17'd5482,17'd5759,17'd5758,17'd5759,17'd24800,17'd24482,17'd24652,17'd12465,17'd25226,17'd12306,17'd14047,17'd14971,17'd22420,17'd26585,17'd26585,17'd16955,17'd18134,17'd18620,17'd18742,17'd22420,17'd19480,17'd19481,17'd22944,17'd21774,17'd19224,17'd26586,17'd26000,17'd26587,17'd24947,17'd19228,17'd16254,17'd26588,17'd18265,17'd26589,17'd26590,17'd26591,17'd26592,17'd26593,17'd26594,17'd18759,17'd2250,17'd26595,17'd1383,17'd777,17'd2100,17'd26596,17'd26465,17'd24668,17'd25642,17'd26597,17'd25895,17'd26339,17'd26339,17'd26598,17'd26598,17'd25896,17'd25896,17'd25644,17'd26599,17'd24816,17'd24670,17'd26123,17'd26012,17'd24168,17'd24169,17'd5781,17'd25105,17'd25105,17'd5781,17'd5945,17'd16960,17'd3400,17'd4233,17'd6243,17'd5037,17'd26600,17'd26233,17'd26601,17'd26602,17'd26603,17'd26467,17'd26604,17'd254,17'd18387,17'd15240
},
'{
17'd4891,17'd4892,17'd3252,17'd1127,17'd3,17'd1275,17'd1275,17'd1275,17'd2933,17'd2933,17'd2933,17'd8814,17'd2423,17'd3430,17'd4247,17'd4247,17'd4247,17'd2595,17'd8971,17'd3430,17'd1128,17'd11,17'd21,17'd21,17'd10,17'd11,17'd980,17'd980,17'd980,17'd980,17'd980,17'd1278,17'd652,17'd652,17'd4431,17'd5207,17'd26468,17'd5803,17'd12931,17'd26605,17'd26606,17'd26470,17'd26471,17'd6603,17'd26472,17'd26237,17'd11346,17'd11457,17'd11613,17'd26607,17'd26474,17'd26348,17'd5067,17'd13309,17'd3448,17'd26608,17'd26609,17'd18766,17'd26610,17'd26611,17'd26612,17'd26481,17'd26481,17'd23151,17'd18410,17'd17809,17'd13599,17'd13093,17'd12955,17'd13094,17'd12218,17'd11764,17'd11629,17'd19621,17'd19754,17'd16766,17'd16518,17'd21649,17'd17572,17'd16289,17'd18060,17'd18776,17'd16169,17'd16169,17'd16169,17'd24348,17'd17319,17'd16289,17'd21650,17'd21650,17'd21650,17'd16164,17'd10565,17'd9703,17'd10694,17'd12534,17'd4767,17'd5089,17'd8846,17'd26354,17'd7920,17'd7924,17'd9020,17'd12824,17'd16295,17'd26483,17'd25516,17'd25400,17'd25661,17'd13615,17'd11485,17'd14232,17'd9593,17'd26613,17'd26614,17'd23842,17'd26027,17'd26615,17'd26616,17'd26617,17'd26618,17'd26619,17'd26620,17'd26621,17'd11510,17'd26622,17'd11511,17'd11659,17'd16547,17'd11504,17'd12099,17'd26623,17'd12851,17'd26624,17'd10725,17'd26625,17'd19156,17'd10329,17'd9344,17'd26626,17'd18080,17'd15048,17'd10326,17'd10854,17'd11397,17'd13516,17'd19157,17'd12861,17'd12577,17'd13884,17'd14930,17'd26627,17'd21207,17'd12416,17'd18200,17'd25927,17'd26371,17'd24857,17'd26628,17'd26150,17'd26495,17'd24031,17'd24537,17'd24856,17'd26629,17'd26373,17'd12254,17'd19408,17'd18443,17'd13516,17'd11396,17'd16069,17'd11667,17'd13253,17'd11962,17'd12115,17'd10854,17'd24996,17'd10166,17'd11133,17'd10991,17'd13886,17'd17236,17'd11398,17'd11398,17'd21206,17'd19282,17'd10991,17'd11133,17'd10476,17'd17838,17'd24035,17'd26630,17'd11276,17'd9620,17'd9346,17'd8874,17'd9348,17'd8725,17'd8726,17'd8724,17'd9040,17'd15684,17'd10174,17'd9620,17'd9741,17'd11671,17'd11670,17'd10475,17'd10990,17'd14810,17'd14673,17'd14673,17'd16068,17'd11522,17'd11522,17'd16068,17'd14673,17'd14931,17'd14931,17'd11399,17'd11399,17'd11399,17'd13886,17'd11133,17'd10741,17'd9739,17'd15048,17'd16065,17'd14674,17'd16552,17'd26631,17'd26632,17'd26633,17'd26634,17'd26635,17'd26636,17'd26637,17'd26638,17'd26639,17'd26640,17'd26641,17'd26642,17'd26643,17'd26644,17'd26645,17'd26646,17'd26647,17'd26648,17'd26649,17'd26650,17'd26651,17'd24888,17'd25424,17'd25825,17'd26521,17'd25308,17'd25826,17'd25551,17'd25551,17'd26522,17'd26522,17'd26276,17'd26652,17'd26523,17'd25557,17'd25698,17'd25558,17'd25554,17'd26524,17'd26524,17'd25944,17'd26653,17'd26279,17'd25702,17'd24892,17'd26654,17'd26655,17'd26281,17'd26656,17'd26657,17'd23727,17'd26658,17'd25832,17'd25704,17'd25313,17'd25945,17'd25429,17'd25312,17'd25312,17'd25561,17'd25172,17'd25704,17'd25172,17'd23718,17'd24240,17'd26659,17'd26660,17'd24891,17'd24891,17'd26530,17'd26174,17'd26661,17'd26662,17'd26663,17'd26664,17'd26665,17'd23752,17'd26666,17'd26667,17'd26668,17'd26669,17'd26670,17'd26671,17'd25735,17'd26544,17'd26672,17'd26673,17'd26674,17'd26675,17'd26676,17'd26547,17'd26677,17'd26678,17'd26550,17'd26679,17'd26680,17'd26085,17'd25736,17'd26084,17'd26681,17'd26682,17'd26683,17'd26684,17'd26685,17'd26686,17'd26687,17'd26311,17'd19327,17'd18010,17'd19680,17'd18728,17'd19330,17'd26562,17'd19069,17'd26688,17'd26689,17'd26690,17'd26691,17'd26692,17'd26693,17'd26694,17'd26695,17'd26696,17'd26697,17'd26698,17'd26699,17'd26700,17'd26701,17'd20231,17'd26702,17'd26703,17'd26704,17'd26705,17'd26706,17'd26445,17'd26707,17'd25078,17'd24940,17'd25765,17'd21301,17'd21141,17'd26581,17'd12136,17'd11692,17'd26584,17'd10196,17'd9907,17'd6547,17'd5914,17'd26451,17'd24800,17'd6388,17'd6218,17'd26708,17'd26709,17'd10513,17'd10641,17'd10641,17'd10641,17'd26219,17'd8303,17'd5159,17'd5612,17'd5611,17'd5482,17'd5759,17'd5758,17'd5759,17'd24800,17'd6706,17'd24652,17'd12466,17'd12465,17'd12306,17'd13165,17'd14970,17'd22420,17'd17066,17'd26585,17'd26710,17'd19590,17'd18260,17'd18742,17'd22420,17'd19480,17'd19848,17'd26711,17'd21311,17'd25088,17'd23981,17'd26712,17'd26713,17'd26220,17'd18378,17'd25775,17'd26714,17'd23292,17'd26715,17'd26716,17'd26717,17'd26718,17'd26719,17'd26720,17'd26721,17'd3587,17'd4084,17'd413,17'd777,17'd26228,17'd2244,17'd26465,17'd24668,17'd26722,17'd26723,17'd26724,17'd26725,17'd26725,17'd26598,17'd26598,17'd26726,17'd25896,17'd25644,17'd26599,17'd23993,17'd23993,17'd26727,17'd26124,17'd24168,17'd24169,17'd5781,17'd25105,17'd24330,17'd25105,17'd5945,17'd16257,17'd3228,17'd3574,17'd4407,17'd6249,17'd3579,17'd6252,17'd4076,17'd26602,17'd26603,17'd2112,17'd2588,17'd456,17'd26728,17'd17789
},
'{
17'd4425,17'd4892,17'd3252,17'd1127,17'd12,17'd806,17'd806,17'd806,17'd806,17'd8814,17'd8814,17'd16747,17'd16636,17'd8971,17'd2594,17'd2594,17'd4247,17'd2595,17'd8971,17'd13,17'd1128,17'd11,17'd21,17'd21,17'd11,17'd11,17'd652,17'd652,17'd652,17'd652,17'd980,17'd980,17'd652,17'd652,17'd4430,17'd26729,17'd26730,17'd5973,17'd26731,17'd5810,17'd26732,17'd26733,17'd6444,17'd26734,17'd26735,17'd11346,17'd11457,17'd6754,17'd26736,17'd12041,17'd26737,17'd26738,17'd26739,17'd3766,17'd3448,17'd21480,17'd20281,17'd18525,17'd18402,17'd26611,17'd26740,17'd23668,17'd26741,17'd23151,17'd18532,17'd17809,17'd17096,17'd17096,17'd13211,17'd13094,17'd12530,17'd11764,17'd11362,17'd19621,17'd16766,17'd16986,17'd15765,17'd16289,17'd18657,17'd16164,17'd17320,17'd17448,17'd17690,17'd17690,17'd18657,17'd17207,17'd18656,17'd17206,17'd21650,17'd21650,17'd16164,17'd16164,17'd10565,17'd9703,17'd10694,17'd10430,17'd5254,17'd6138,17'd25803,17'd8076,17'd26742,17'd8857,17'd9315,17'd9589,17'd25131,17'd15405,17'd25516,17'd25400,17'd10131,17'd11097,17'd11485,17'd11923,17'd12075,17'd26743,17'd23330,17'd26744,17'd26745,17'd26746,17'd26747,17'd17464,17'd26748,17'd26749,17'd26750,17'd25922,17'd26751,17'd26752,17'd26753,17'd11506,17'd11793,17'd13248,17'd19275,17'd12851,17'd15043,17'd11117,17'd26754,17'd10986,17'd10325,17'd17012,17'd9339,17'd15180,17'd24037,17'd9739,17'd11132,17'd11274,17'd13516,17'd12422,17'd11962,17'd12718,17'd12256,17'd12859,17'd14003,17'd26755,17'd21504,17'd19534,17'd18084,17'd24991,17'd24859,17'd26756,17'd26628,17'd26372,17'd24705,17'd24031,17'd24856,17'd26757,17'd26758,17'd23855,17'd14807,17'd17603,17'd16204,17'd13516,17'd13762,17'd11667,17'd13253,17'd13253,17'd11395,17'd20910,17'd19532,17'd10329,17'd10165,17'd10991,17'd10603,17'd16320,17'd14931,17'd11808,17'd11524,17'd21206,17'd19282,17'd11132,17'd10476,17'd13001,17'd12862,17'd13138,17'd26037,17'd9741,17'd23679,17'd9347,17'd8873,17'd8566,17'd8882,17'd15297,17'd24999,17'd23859,17'd15807,17'd9479,17'd9741,17'd17719,17'd10164,17'd10603,17'd10604,17'd11519,17'd11519,17'd11395,17'd11395,17'd13762,17'd11807,17'd13762,17'd16069,17'd16069,17'd12720,17'd14810,17'd17236,17'd17236,17'd17236,17'd10605,17'd10991,17'd17720,17'd11528,17'd26759,17'd24998,17'd25408,17'd15807,17'd16552,17'd26760,17'd26761,17'd26762,17'd26763,17'd26764,17'd26765,17'd26766,17'd26767,17'd26768,17'd26769,17'd26770,17'd26771,17'd26772,17'd26773,17'd26774,17'd26775,17'd26776,17'd26649,17'd26777,17'd26778,17'd26779,17'd25548,17'd24402,17'd24577,17'd25308,17'd25551,17'd25551,17'd25551,17'd26522,17'd26522,17'd26277,17'd26652,17'd26780,17'd25557,17'd25698,17'd25558,17'd25554,17'd25558,17'd26780,17'd25557,17'd26394,17'd26167,17'd26400,17'd24891,17'd24739,17'd23729,17'd23382,17'd24083,17'd24899,17'd23726,17'd26658,17'd25434,17'd25431,17'd25948,17'd25311,17'd26279,17'd26781,17'd26782,17'd25561,17'd25172,17'd25172,17'd25430,17'd24239,17'd23719,17'd26168,17'd24408,17'd24583,17'd23908,17'd24736,17'd24582,17'd25708,17'd26783,17'd26784,17'd26785,17'd26786,17'd26787,17'd26788,17'd26789,17'd26790,17'd26791,17'd26792,17'd26793,17'd25342,17'd26794,17'd26795,17'd26796,17'd24756,17'd26797,17'd26675,17'd25843,17'd26798,17'd26551,17'd26799,17'd25589,17'd25845,17'd26800,17'd26195,17'd25853,17'd25852,17'd26801,17'd26802,17'd23764,17'd19437,17'd22367,17'd26803,17'd26804,17'd26805,17'd17769,17'd19567,17'd26562,17'd26806,17'd19816,17'd25616,17'd26806,17'd26807,17'd26808,17'd26809,17'd26810,17'd26811,17'd26812,17'd26813,17'd26814,17'd26815,17'd26816,17'd26817,17'd26818,17'd26819,17'd26820,17'd26821,17'd26822,17'd26823,17'd26824,17'd26825,17'd26444,17'd26707,17'd21608,17'd24940,17'd21451,17'd21301,17'd21452,17'd26581,17'd12136,17'd12741,17'd26826,17'd10196,17'd9907,17'd26827,17'd5913,17'd26451,17'd24800,17'd6387,17'd6387,17'd6218,17'd26709,17'd8304,17'd10513,17'd10777,17'd11576,17'd10641,17'd8154,17'd6389,17'd5158,17'd5611,17'd5481,17'd5482,17'd5481,17'd5759,17'd5760,17'd26828,17'd6392,17'd24652,17'd26829,17'd25226,17'd24653,17'd13925,17'd15476,17'd17904,17'd17904,17'd26585,17'd16955,17'd18260,17'd18022,17'd22420,17'd19480,17'd19223,17'd26711,17'd19849,17'd25088,17'd26830,17'd22091,17'd26831,17'd25486,17'd26832,17'd25775,17'd26714,17'd14431,17'd22949,17'd26833,17'd26834,17'd26718,17'd26835,17'd26836,17'd26837,17'd26838,17'd1380,17'd602,17'd777,17'd26839,17'd26596,17'd2396,17'd24500,17'd24668,17'd26840,17'd26841,17'd26725,17'd26722,17'd26842,17'd26598,17'd26842,17'd26842,17'd25896,17'd24326,17'd23993,17'd23818,17'd26843,17'd24824,17'd5782,17'd23482,17'd5781,17'd25105,17'd24330,17'd25105,17'd5945,17'd16257,17'd3228,17'd3574,17'd4407,17'd5037,17'd26844,17'd4414,17'd4076,17'd26602,17'd26845,17'd21161,17'd2588,17'd460,17'd1123,17'd26728
},
'{
17'd4425,17'd4243,17'd3252,17'd1127,17'd12,17'd2423,17'd806,17'd806,17'd806,17'd806,17'd806,17'd2423,17'd3430,17'd2595,17'd1831,17'd1831,17'd4247,17'd4247,17'd466,17'd13,17'd1128,17'd11,17'd21,17'd21,17'd11,17'd1128,17'd652,17'd652,17'd652,17'd652,17'd980,17'd980,17'd652,17'd28,17'd6744,17'd6438,17'd5973,17'd26846,17'd5977,17'd5810,17'd26732,17'd26847,17'd6444,17'd6603,17'd26472,17'd6753,17'd26238,17'd6754,17'd6447,17'd4266,17'd26848,17'd26738,17'd22792,17'd3766,17'd2626,17'd26849,17'd4108,17'd18999,17'd26850,17'd26851,17'd26852,17'd26853,17'd26854,17'd23152,17'd25802,17'd17809,17'd23325,17'd17096,17'd13094,17'd12362,17'd11764,17'd11362,17'd17204,17'd19754,17'd21649,17'd16986,17'd16164,17'd17207,17'd18657,17'd19256,17'd17448,17'd17810,17'd17690,17'd17445,17'd17207,17'd17319,17'd17206,17'd17206,17'd21650,17'd21650,17'd16164,17'd15766,17'd10113,17'd9007,17'd10430,17'd9302,17'd5252,17'd8846,17'd26855,17'd8385,17'd26856,17'd8856,17'd9589,17'd16180,17'd15540,17'd15405,17'd26857,17'd26024,17'd11097,17'd26858,17'd11923,17'd12074,17'd21196,17'd9714,17'd26859,17'd26860,17'd26861,17'd26862,17'd26863,17'd26748,17'd26864,17'd26865,17'd11258,17'd12852,17'd22471,17'd13878,17'd26363,17'd11505,17'd11793,17'd12246,17'd26866,17'd18075,17'd11258,17'd26867,17'd26868,17'd26869,17'd26870,17'd10857,17'd10857,17'd10742,17'd25673,17'd10022,17'd10990,17'd11964,17'd17604,17'd16204,17'd11961,17'd12413,17'd12578,17'd12417,17'd13515,17'd25279,17'd19534,17'd24991,17'd25528,17'd24856,17'd25526,17'd26494,17'd26628,17'd26871,17'd24031,17'd24537,17'd26872,17'd26873,17'd26758,17'd20452,17'd17602,17'd18917,17'd12996,17'd13762,17'd13762,17'd11667,17'd13253,17'd11666,17'd10737,17'd10475,17'd10166,17'd10330,17'd11133,17'd10476,17'd10739,17'd10990,17'd11808,17'd11808,17'd11524,17'd21206,17'd19282,17'd11132,17'd10605,17'd26497,17'd12862,17'd13886,17'd11134,17'd9479,17'd9346,17'd9347,17'd8720,17'd26874,17'd9045,17'd17123,17'd24361,17'd15807,17'd9479,17'd11277,17'd11134,17'd10326,17'd10603,17'd24860,17'd11519,17'd11520,17'd11520,17'd13762,17'd13762,17'd11807,17'd11667,17'd11807,17'd16069,17'd13000,17'd15182,17'd12720,17'd13138,17'd13138,17'd17236,17'd11399,17'd11132,17'd10991,17'd12863,17'd10479,17'd14928,17'd15566,17'd17965,17'd26875,17'd26876,17'd26877,17'd26878,17'd26879,17'd26880,17'd26881,17'd26882,17'd26883,17'd26884,17'd26885,17'd26886,17'd26887,17'd26888,17'd26889,17'd26890,17'd26891,17'd26892,17'd26893,17'd26894,17'd26895,17'd26896,17'd26779,17'd24889,17'd24399,17'd25170,17'd25551,17'd25551,17'd25551,17'd26897,17'd26522,17'd26277,17'd26652,17'd26780,17'd25828,17'd25554,17'd25558,17'd25558,17'd26780,17'd26780,17'd25557,17'd26898,17'd25429,17'd25945,17'd24736,17'd25176,17'd26899,17'd24741,17'd24900,17'd26900,17'd25028,17'd23910,17'd24737,17'd24582,17'd25561,17'd25312,17'd26167,17'd26901,17'd26902,17'd25948,17'd25561,17'd25430,17'd25313,17'd23907,17'd23907,17'd25562,17'd26168,17'd26168,17'd25431,17'd25172,17'd25561,17'd26903,17'd26904,17'd26905,17'd26906,17'd26907,17'd26908,17'd25188,17'd26909,17'd26910,17'd26911,17'd26912,17'd26670,17'd26913,17'd26914,17'd26795,17'd26915,17'd26916,17'd26917,17'd26918,17'd25843,17'd25342,17'd26919,17'd26678,17'd26417,17'd25338,17'd25737,17'd26540,17'd26920,17'd26194,17'd26921,17'd26922,17'd26923,17'd26924,17'd26925,17'd26926,17'd26927,17'd26928,17'd18007,17'd17771,17'd26562,17'd18735,17'd19681,17'd19710,17'd26929,17'd26930,17'd26931,17'd26932,17'd26810,17'd26933,17'd26934,17'd26935,17'd26936,17'd26937,17'd26938,17'd26939,17'd26940,17'd26941,17'd26942,17'd26943,17'd26944,17'd26945,17'd26946,17'd21918,17'd26947,17'd26948,17'd26707,17'd25479,17'd25480,17'd25765,17'd21301,17'd26446,17'd26581,17'd26582,17'd12741,17'd26826,17'd9907,17'd6546,17'd6548,17'd5482,17'd24800,17'd6387,17'd6387,17'd6553,17'd26709,17'd8303,17'd9657,17'd10513,17'd11576,17'd11576,17'd10513,17'd26709,17'd5159,17'd5612,17'd5481,17'd5482,17'd5481,17'd5758,17'd5482,17'd26949,17'd6221,17'd10237,17'd24652,17'd12465,17'd25085,17'd13558,17'd15340,17'd15476,17'd15476,17'd26585,17'd16955,17'd18742,17'd18022,17'd22420,17'd19480,17'd18853,17'd12163,17'd19849,17'd26950,17'd26951,17'd26454,17'd26952,17'd26953,17'd26954,17'd26955,17'd26956,17'd24157,17'd26957,17'd26958,17'd26959,17'd26960,17'd26961,17'd26962,17'd26963,17'd26964,17'd1678,17'd412,17'd26965,17'd26966,17'd2244,17'd2395,17'd24499,17'd26722,17'd26723,17'd26723,17'd26967,17'd26967,17'd26968,17'd26969,17'd26842,17'd26725,17'd25896,17'd24326,17'd24171,17'd23993,17'd23994,17'd23995,17'd23133,17'd23482,17'd5780,17'd25105,17'd24330,17'd25105,17'd26970,17'd16257,17'd3228,17'd3398,17'd4062,17'd4064,17'd12486,17'd4414,17'd4076,17'd3238,17'd23301,17'd21161,17'd2588,17'd967,17'd965,17'd26728
},
'{
17'd4425,17'd4243,17'd3252,17'd1127,17'd2,17'd13,17'd12,17'd3,17'd3,17'd806,17'd806,17'd2423,17'd3430,17'd15745,17'd1831,17'd1688,17'd4247,17'd2595,17'd3430,17'd13,17'd1128,17'd20,17'd21,17'd20,17'd11,17'd1128,17'd652,17'd652,17'd652,17'd652,17'd980,17'd980,17'd652,17'd6744,17'd6437,17'd6438,17'd5973,17'd26971,17'd5977,17'd26972,17'd26973,17'd26974,17'd5225,17'd26734,17'd26735,17'd26975,17'd11457,17'd26976,17'd26977,17'd26978,17'd26979,17'd26980,17'd26981,17'd2625,17'd14197,17'd26982,17'd18524,17'd26983,17'd18050,17'd26984,17'd26985,17'd26853,17'd26854,17'd23836,17'd25802,17'd17096,17'd17096,17'd17096,17'd12362,17'd13969,17'd12681,17'd17204,17'd23155,17'd16986,17'd21649,17'd19384,17'd17319,17'd17207,17'd17319,17'd18060,17'd17810,17'd17810,17'd17445,17'd17320,17'd19255,17'd18656,17'd18174,17'd17205,17'd16986,17'd16986,17'd19384,17'd15766,17'd10113,17'd9007,17'd9302,17'd5254,17'd5252,17'd8846,17'd8076,17'd7761,17'd8078,17'd8856,17'd9589,17'd26986,17'd26987,17'd15405,17'd14783,17'd13734,17'd11485,17'd11923,17'd26988,17'd26989,17'd25266,17'd26990,17'd26991,17'd26992,17'd26993,17'd9326,17'd26994,17'd26619,17'd15416,17'd26995,17'd10972,17'd12991,17'd26996,17'd18190,17'd18438,17'd26997,17'd11652,17'd18912,17'd11795,17'd26998,17'd26999,17'd27000,17'd27001,17'd27002,17'd27003,17'd9341,17'd10743,17'd17011,17'd25673,17'd10606,17'd14673,17'd18444,17'd16204,17'd12858,17'd12110,17'd13514,17'd15434,17'd14807,17'd19407,17'd12255,17'd25528,17'd25528,17'd25528,17'd24537,17'd24705,17'd26494,17'd26871,17'd24031,17'd24537,17'd27004,17'd26757,17'd27005,17'd25925,17'd20314,17'd12582,17'd16204,17'd13362,17'd11963,17'd12996,17'd13135,17'd11667,17'd11395,17'd10739,17'd10326,17'd26152,17'd11670,17'd11132,17'd11399,17'd11808,17'd11965,17'd10990,17'd10990,17'd11132,17'd19282,17'd11525,17'd11399,17'd17838,17'd15432,17'd11519,17'd16555,17'd9741,17'd9345,17'd9346,17'd9043,17'd9044,17'd9044,17'd10174,17'd14674,17'd9479,17'd9885,17'd9884,17'd12863,17'd11132,17'd10739,17'd10604,17'd16435,17'd15186,17'd11963,17'd11963,17'd12996,17'd12996,17'd11806,17'd13646,17'd11667,17'd11520,17'd11666,17'd12862,17'd14810,17'd17236,17'd13138,17'd17236,17'd11399,17'd11131,17'd10475,17'd11133,17'd10479,17'd11134,17'd11277,17'd12116,17'd17841,17'd27006,17'd27007,17'd27008,17'd27009,17'd27010,17'd27011,17'd27012,17'd27013,17'd27014,17'd27015,17'd27016,17'd27017,17'd27018,17'd27019,17'd27020,17'd27021,17'd27022,17'd27023,17'd26165,17'd27024,17'd26896,17'd26779,17'd24400,17'd24402,17'd25170,17'd25551,17'd25551,17'd25826,17'd25826,17'd25826,17'd26652,17'd25697,17'd25555,17'd25554,17'd25558,17'd26524,17'd26523,17'd26523,17'd26780,17'd25828,17'd25429,17'd25429,17'd25945,17'd27025,17'd23909,17'd27026,17'd24894,17'd23560,17'd23727,17'd23725,17'd23910,17'd25434,17'd24891,17'd24736,17'd25172,17'd26400,17'd27027,17'd26902,17'd25948,17'd25561,17'd24239,17'd24073,17'd25945,17'd25311,17'd25562,17'd25562,17'd25562,17'd25703,17'd25311,17'd25312,17'd25702,17'd27028,17'd27029,17'd27030,17'd27031,17'd27032,17'd27033,17'd27034,17'd27035,17'd27036,17'd27037,17'd27038,17'd26792,17'd27039,17'd27040,17'd27041,17'd25049,17'd27042,17'd27043,17'd27044,17'd25736,17'd27045,17'd27046,17'd26678,17'd27047,17'd27048,17'd27049,17'd26540,17'd27050,17'd27051,17'd27052,17'd27053,17'd27054,17'd27055,17'd27056,17'd27057,17'd27058,17'd27059,17'd17771,17'd18728,17'd18605,17'd18014,17'd19451,17'd25616,17'd27060,17'd27061,17'd20986,17'd27062,17'd27063,17'd27064,17'd27065,17'd27066,17'd27067,17'd27068,17'd26816,17'd27069,17'd27070,17'd27071,17'd27072,17'd27073,17'd27074,17'd27075,17'd27076,17'd21762,17'd27077,17'd26580,17'd25479,17'd25480,17'd21451,17'd21924,17'd21766,17'd27078,17'd27079,17'd27080,17'd11294,17'd10196,17'd6545,17'd26827,17'd5610,17'd5760,17'd6387,17'd6387,17'd6706,17'd6218,17'd8303,17'd8154,17'd10513,17'd11576,17'd11853,17'd10777,17'd8154,17'd6389,17'd5158,17'd5158,17'd5482,17'd5481,17'd5758,17'd5482,17'd26949,17'd27081,17'd6852,17'd10237,17'd12465,17'd25226,17'd14301,17'd18621,17'd15476,17'd15340,17'd17904,17'd18022,17'd18742,17'd18022,17'd22420,17'd19480,17'd27082,17'd12308,17'd24804,17'd27083,17'd27084,17'd23288,17'd26000,17'd17411,17'd27085,17'd14430,17'd27086,17'd18379,17'd27087,17'd27088,17'd25491,17'd27089,17'd27090,17'd27091,17'd27092,17'd27093,17'd16858,17'd2740,17'd27094,17'd1950,17'd2100,17'd2395,17'd2396,17'd24668,17'd26840,17'd26723,17'd27095,17'd26967,17'd26723,17'd26968,17'd26725,17'd26725,17'd25643,17'd24326,17'd23993,17'd23818,17'd27096,17'd23995,17'd23133,17'd23134,17'd5780,17'd5781,17'd25646,17'd24824,17'd27096,17'd16257,17'd3228,17'd3399,17'd4232,17'd5037,17'd26844,17'd4414,17'd3732,17'd3238,17'd9662,17'd21161,17'd263,17'd264,17'd254,17'd26728
},
'{
17'd27097,17'd4892,17'd2422,17'd1127,17'd2,17'd13,17'd13,17'd12,17'd12,17'd3,17'd806,17'd13,17'd2595,17'd2594,17'd1831,17'd3250,17'd1688,17'd4247,17'd466,17'd13,17'd1128,17'd20,17'd20,17'd20,17'd1128,17'd1128,17'd652,17'd652,17'd652,17'd652,17'd980,17'd980,17'd652,17'd28,17'd6744,17'd6438,17'd5973,17'd26971,17'd5977,17'd5810,17'd5661,17'd5524,17'd27098,17'd6603,17'd26472,17'd26975,17'd11457,17'd11613,17'd6448,17'd27099,17'd27100,17'd3765,17'd27101,17'd27102,17'd27103,17'd26133,17'd18525,17'd18768,17'd27104,17'd27105,17'd26985,17'd26853,17'd24840,17'd27106,17'd17940,17'd13211,17'd17096,17'd13094,17'd12361,17'd12681,17'd17941,17'd19893,17'd27107,17'd17206,17'd19384,17'd16164,17'd18657,17'd17207,17'd16289,17'd17445,17'd17942,17'd17575,17'd18776,17'd17319,17'd17206,17'd17206,17'd18174,17'd18174,17'd16986,17'd16986,17'd19384,17'd15898,17'd9703,17'd8066,17'd5254,17'd5252,17'd8846,17'd8542,17'd7760,17'd7264,17'd8855,17'd15402,17'd16531,17'd25131,17'd26987,17'd14642,17'd10437,17'd11097,17'd27108,17'd26988,17'd27109,17'd27110,17'd21353,17'd27111,17'd24690,17'd27112,17'd9458,17'd27113,17'd27114,17'd27115,17'd26620,17'd26750,17'd15937,17'd18555,17'd26996,17'd18190,17'd11950,17'd15043,17'd11507,17'd11949,17'd27116,17'd27117,17'd27118,17'd27119,17'd27120,17'd10741,17'd9341,17'd10743,17'd10742,17'd9741,17'd11134,17'd13886,17'd11522,17'd18444,17'd12996,17'd12857,17'd12414,17'd15434,17'd12253,17'd14807,17'd12108,17'd23855,17'd25528,17'd27121,17'd24856,17'd24030,17'd23170,17'd23170,17'd27122,17'd24857,17'd27121,17'd26629,17'd26757,17'd27123,17'd24030,17'd18559,17'd18806,17'd12262,17'd12262,17'd11963,17'd13135,17'd11806,17'd11667,17'd11274,17'd19532,17'd10023,17'd11134,17'd11527,17'd10476,17'd11275,17'd13516,17'd13645,17'd11275,17'd10990,17'd19282,17'd19532,17'd12423,17'd24364,17'd24035,17'd15182,17'd10737,17'd10473,17'd9741,17'd9344,17'd9189,17'd15682,17'd8720,17'd10174,17'd14674,17'd9479,17'd9884,17'd10329,17'd11400,17'd11399,17'd14931,17'd14262,17'd11395,17'd15186,17'd11963,17'd11962,17'd13135,17'd13135,17'd11806,17'd11961,17'd13646,17'd13520,17'd11807,17'd11395,17'd14931,17'd10854,17'd21206,17'd11399,17'd11524,17'd11524,17'd10854,17'd10854,17'd11132,17'd11133,17'd10326,17'd10479,17'd11134,17'd17847,17'd17479,17'd27124,17'd27125,17'd27126,17'd27127,17'd27128,17'd27129,17'd27130,17'd27131,17'd27132,17'd27133,17'd27134,17'd27135,17'd27136,17'd27137,17'd27138,17'd27139,17'd27140,17'd27141,17'd27142,17'd27143,17'd25548,17'd27144,17'd26053,17'd25170,17'd25551,17'd25551,17'd25826,17'd25826,17'd25826,17'd26652,17'd26780,17'd25554,17'd25554,17'd25558,17'd26524,17'd26523,17'd26523,17'd26652,17'd26780,17'd25553,17'd25559,17'd25698,17'd27145,17'd25832,17'd24078,17'd23557,17'd26899,17'd23913,17'd23725,17'd24078,17'd24892,17'd24891,17'd24891,17'd24582,17'd25699,17'd27027,17'd27027,17'd25702,17'd25948,17'd23907,17'd24073,17'd26394,17'd25429,17'd25561,17'd25562,17'd25703,17'd25702,17'd26279,17'd26279,17'd26279,17'd27146,17'd27147,17'd27148,17'd27149,17'd27150,17'd27151,17'd27152,17'd27153,17'd27154,17'd27034,17'd27155,17'd27156,17'd26303,17'd27157,17'd27040,17'd27158,17'd27159,17'd27160,17'd25843,17'd27161,17'd27162,17'd27163,17'd27164,17'd27165,17'd25593,17'd27166,17'd27167,17'd27168,17'd27169,17'd27170,17'd26683,17'd27171,17'd27172,17'd27173,17'd27174,17'd27175,17'd27176,17'd17647,17'd19567,17'd27177,17'd18014,17'd19568,17'd19817,17'd27178,17'd24465,17'd27179,17'd27180,17'd27181,17'd27182,17'd27183,17'd27184,17'd27185,17'd27186,17'd27187,17'd27188,17'd27189,17'd27190,17'd27191,17'd27192,17'd27193,17'd22907,17'd27194,17'd27195,17'd21763,17'd21139,17'd21300,17'd27196,17'd21451,17'd21451,17'd21924,17'd21610,17'd12281,17'd27197,17'd11013,17'd9503,17'd6545,17'd5148,17'd4843,17'd5482,17'd6387,17'd6387,17'd24482,17'd6387,17'd6553,17'd8154,17'd9657,17'd10641,17'd11853,17'd10641,17'd9394,17'd26709,17'd26218,17'd5331,17'd5482,17'd5481,17'd5610,17'd5481,17'd5762,17'd26828,17'd6852,17'd10237,17'd12466,17'd12465,17'd12760,17'd27198,17'd15340,17'd15340,17'd15476,17'd22420,17'd18022,17'd18022,17'd22420,17'd19480,17'd27199,17'd13408,17'd24804,17'd27083,17'd24313,17'd27200,17'd19718,17'd17286,17'd18377,17'd14974,17'd27201,17'd18379,17'd26004,17'd27202,17'd27203,17'd27089,17'd27204,17'd27205,17'd27206,17'd27207,17'd1239,17'd6407,17'd5631,17'd1949,17'd2100,17'd2242,17'd2396,17'd2563,17'd27208,17'd27209,17'd27095,17'd27095,17'd27209,17'd26723,17'd26725,17'd26725,17'd25643,17'd25644,17'd23993,17'd23993,17'd23994,17'd23995,17'd23133,17'd23134,17'd5637,17'd5781,17'd24824,17'd23995,17'd27096,17'd24167,17'd23989,17'd3399,17'd4232,17'd4408,17'd3234,17'd26844,17'd9249,17'd9533,17'd9662,17'd10073,17'd257,17'd263,17'd456,17'd965
},
'{
17'd27097,17'd4892,17'd2422,17'd1127,17'd466,17'd3430,17'd3430,17'd13,17'd13,17'd12,17'd12,17'd3430,17'd15745,17'd17917,17'd7545,17'd7711,17'd1831,17'd2595,17'd3430,17'd16636,17'd2598,17'd20,17'd20,17'd20,17'd980,17'd980,17'd653,17'd653,17'd652,17'd652,17'd980,17'd980,17'd652,17'd6744,17'd6437,17'd5973,17'd26971,17'd26971,17'd27210,17'd26972,17'd27211,17'd5523,17'd5387,17'd27212,17'd27213,17'd11346,17'd26345,17'd26736,17'd5527,17'd27214,17'd27100,17'd3765,17'd3447,17'd13442,17'd27215,17'd4107,17'd25255,17'd14997,17'd24010,17'd27216,17'd26985,17'd26612,17'd25658,17'd27106,17'd17940,17'd17940,17'd12815,17'd12362,17'd13969,17'd27217,17'd27218,17'd17204,17'd16766,17'd16986,17'd16164,17'd16519,17'd17690,17'd17320,17'd15899,17'd17690,17'd17942,17'd27219,17'd19011,17'd21185,17'd17206,17'd18174,17'd18655,17'd18655,17'd17206,17'd16986,17'd19384,17'd15898,17'd9703,17'd4611,17'd5254,17'd6138,17'd24841,17'd8382,17'd7761,17'd27220,17'd8856,17'd15402,17'd16531,17'd26987,17'd15405,17'd14642,17'd27221,17'd13855,17'd12223,17'd26989,17'd27222,17'd27223,17'd26744,17'd23158,17'd27224,17'd27225,17'd27226,17'd27227,17'd15417,17'd27228,17'd27229,17'd27230,17'd16904,17'd11265,17'd26996,17'd27231,17'd26367,17'd11794,17'd11660,17'd18075,17'd11258,17'd26999,17'd27232,17'd27233,17'd9882,17'd9741,17'd13255,17'd9480,17'd17011,17'd9739,17'd10991,17'd17236,17'd18327,17'd19158,17'd11806,17'd12718,17'd12578,17'd12253,17'd14807,17'd14807,17'd18564,17'd18200,17'd26872,17'd26370,17'd24537,17'd23512,17'd24209,17'd24209,17'd24538,17'd24537,17'd27234,17'd27235,17'd26629,17'd24537,17'd23170,17'd22472,17'd19158,17'd15810,17'd19157,17'd12999,17'd12113,17'd13135,17'd13762,17'd11130,17'd10166,17'd9883,17'd11528,17'd26037,17'd11524,17'd11275,17'd13516,17'd13645,17'd11275,17'd10854,17'd11132,17'd19282,17'd16687,17'd24035,17'd13000,17'd16068,17'd25144,17'd27236,17'd10742,17'd9743,17'd9043,17'd8874,17'd15944,17'd17716,17'd16549,17'd19531,17'd19155,17'd12584,17'd11398,17'd11274,17'd14262,17'd15186,17'd16797,17'd11957,17'd11957,17'd12113,17'd12857,17'd12857,17'd11960,17'd11960,17'd11806,17'd12996,17'd13762,17'd11965,17'd11131,17'd14263,17'd14263,17'd11131,17'd11399,17'd17236,17'd11808,17'd10737,17'd10990,17'd10739,17'd10603,17'd14518,17'd11527,17'd12585,17'd17479,17'd27237,17'd27238,17'd27239,17'd27240,17'd27241,17'd27242,17'd27243,17'd27244,17'd27245,17'd27246,17'd27247,17'd27248,17'd27136,17'd27249,17'd27250,17'd27251,17'd27252,17'd27253,17'd27254,17'd25307,17'd25548,17'd27255,17'd25825,17'd25826,17'd25551,17'd25551,17'd25826,17'd25826,17'd25826,17'd25169,17'd24578,17'd25554,17'd25558,17'd25558,17'd26524,17'd26523,17'd26278,17'd26277,17'd26278,17'd25559,17'd26055,17'd25944,17'd27145,17'd27256,17'd27257,17'd25176,17'd27026,17'd23912,17'd23911,17'd23910,17'd24892,17'd24584,17'd23908,17'd25431,17'd25699,17'd27027,17'd27258,17'd25831,17'd25702,17'd23904,17'd23906,17'd26394,17'd26394,17'd26782,17'd27259,17'd27259,17'd26902,17'd25698,17'd25698,17'd25552,17'd26055,17'd27260,17'd27261,17'd27262,17'd27263,17'd27264,17'd27265,17'd27266,17'd27267,17'd26911,17'd27268,17'd27269,17'd27270,17'd25452,17'd27271,17'd27272,17'd25335,17'd27160,17'd25843,17'd26304,17'd26920,17'd27273,17'd27164,17'd27274,17'd25343,17'd27166,17'd27275,17'd27276,17'd27277,17'd26550,17'd27278,17'd27279,17'd27280,17'd27281,17'd27282,17'd27283,17'd27284,17'd17770,17'd19449,17'd27177,17'd18014,17'd19568,17'd25606,17'd27285,17'd24466,17'd20087,17'd27286,17'd27287,17'd27288,17'd27289,17'd27290,17'd27291,17'd27292,17'd27293,17'd27294,17'd27295,17'd27296,17'd27297,17'd27298,17'd27299,17'd27300,17'd20678,17'd27301,17'd27302,17'd27303,17'd21139,17'd21300,17'd21451,17'd21451,17'd25481,17'd21610,17'd12281,17'd27304,17'd27305,17'd7824,17'd24480,17'd6546,17'd5150,17'd5481,17'd6388,17'd6706,17'd24482,17'd6706,17'd6707,17'd8154,17'd8304,17'd10777,17'd11576,17'd10641,17'd26219,17'd6707,17'd5332,17'd5332,17'd5482,17'd5611,17'd5611,17'd5481,17'd5762,17'd26828,17'd5919,17'd6221,17'd9394,17'd12466,17'd11854,17'd14423,17'd17655,17'd15094,17'd17655,17'd17904,17'd18022,17'd22420,17'd22420,17'd18852,17'd27306,17'd27307,17'd24804,17'd27083,17'd27308,17'd27200,17'd27309,17'd17286,17'd18377,17'd15099,17'd27310,17'd18138,17'd16379,17'd27311,17'd27312,17'd27313,17'd27314,17'd27315,17'd27316,17'd25783,17'd27317,17'd4084,17'd14178,17'd27318,17'd2100,17'd2242,17'd2398,17'd24500,17'd26722,17'd26723,17'd27095,17'd27095,17'd27319,17'd27320,17'd26725,17'd26725,17'd25643,17'd25644,17'd24171,17'd23993,17'd23994,17'd24174,17'd5638,17'd23134,17'd5637,17'd5780,17'd24824,17'd23995,17'd27096,17'd16257,17'd3228,17'd3400,17'd4404,17'd4067,17'd26600,17'd26844,17'd9249,17'd27321,17'd9662,17'd10073,17'd257,17'd263,17'd1271,17'd1270
},
'{
17'd27097,17'd4892,17'd2784,17'd1689,17'd466,17'd8971,17'd3430,17'd13,17'd13,17'd13,17'd13,17'd466,17'd15745,17'd17917,17'd7545,17'd7711,17'd2594,17'd2595,17'd3430,17'd13,17'd1128,17'd20,17'd20,17'd1128,17'd980,17'd980,17'd653,17'd653,17'd652,17'd652,17'd980,17'd980,17'd652,17'd6744,17'd6437,17'd6437,17'd5972,17'd26971,17'd27210,17'd27322,17'd5812,17'd5386,17'd6751,17'd27212,17'd26237,17'd11457,17'd26346,17'd27323,17'd4101,17'd27214,17'd27324,17'd27325,17'd3447,17'd14083,17'd27326,17'd25797,17'd25392,17'd18288,17'd24010,17'd27216,17'd26985,17'd26853,17'd25658,17'd20885,17'd17940,17'd12815,17'd12362,17'd12680,17'd11764,17'd27218,17'd19753,17'd19754,17'd17206,17'd16164,17'd18060,17'd17690,17'd17445,17'd16519,17'd16034,17'd17942,17'd19010,17'd27219,17'd19011,17'd21650,17'd16986,17'd18174,17'd18655,17'd17206,17'd17206,17'd16164,17'd19384,17'd15898,17'd9007,17'd4611,17'd5253,17'd9160,17'd27327,17'd25260,17'd27328,17'd27329,17'd9020,17'd15538,17'd26986,17'd26987,17'd15405,17'd15786,17'd10819,17'd27108,17'd27330,17'd27331,17'd27332,17'd9595,17'd27333,17'd24690,17'd27334,17'd27335,17'd27336,17'd27337,17'd27338,17'd27339,17'd27340,17'd26257,17'd27341,17'd11264,17'd11266,17'd11389,17'd27342,17'd16310,17'd18438,17'd26367,17'd27117,17'd27343,17'd27344,17'd27345,17'd22131,17'd9742,17'd13370,17'd9742,17'd9885,17'd11134,17'd13886,17'd11274,17'd21985,17'd16325,17'd11960,17'd12577,17'd15434,17'd12579,17'd17348,17'd12579,17'd16685,17'd18084,17'd26872,17'd27346,17'd27347,17'd24705,17'd24209,17'd24992,17'd24030,17'd24856,17'd27348,17'd27349,17'd26758,17'd23512,17'd21362,17'd18443,17'd19158,17'd11964,17'd11963,17'd12112,17'd12113,17'd16204,17'd13645,17'd14132,17'd10329,17'd11134,17'd20756,17'd14666,17'd14931,17'd19533,17'd13516,17'd13516,17'd11275,17'd10475,17'd11132,17'd19282,17'd17236,17'd16199,17'd15432,17'd14810,17'd10474,17'd10168,17'd9340,17'd9190,17'd9189,17'd17716,17'd25408,17'd16549,17'd11276,17'd14668,17'd27350,17'd13367,17'd11522,17'd11964,17'd13362,17'd11962,17'd12999,17'd12858,17'd12857,17'd12111,17'd12111,17'd12419,17'd13761,17'd11960,17'd13520,17'd11964,17'd10989,17'd11130,17'd14263,17'd16555,17'd10475,17'd11131,17'd10854,17'd10990,17'd10737,17'd14262,17'd14673,17'd14931,17'd16320,17'd13886,17'd10991,17'd11670,17'd27351,17'd27237,17'd27352,17'd27353,17'd27354,17'd27355,17'd27356,17'd27357,17'd27358,17'd27359,17'd27360,17'd27361,17'd27248,17'd27362,17'd27363,17'd27364,17'd27251,17'd27365,17'd27366,17'd27367,17'd25168,17'd24397,17'd25825,17'd25022,17'd25826,17'd25551,17'd25551,17'd25826,17'd25826,17'd25826,17'd25169,17'd24578,17'd25554,17'd25558,17'd26523,17'd26523,17'd26278,17'd26278,17'd26277,17'd26276,17'd27368,17'd27369,17'd25944,17'd25945,17'd25704,17'd24891,17'd25176,17'd24080,17'd23725,17'd24585,17'd27370,17'd26658,17'd24892,17'd24891,17'd24736,17'd25948,17'd27027,17'd27027,17'd25699,17'd25699,17'd23904,17'd23906,17'd26394,17'd26394,17'd27027,17'd27371,17'd27371,17'd26782,17'd25944,17'd25828,17'd25428,17'd25554,17'd27372,17'd27373,17'd27374,17'd27375,17'd27376,17'd27377,17'd27266,17'd27267,17'd27378,17'd27156,17'd27379,17'd27380,17'd27381,17'd27382,17'd27383,17'd27384,17'd27385,17'd26918,17'd26191,17'd27386,17'd27387,17'd27388,17'd27389,17'd25194,17'd26540,17'd27275,17'd27390,17'd27391,17'd27392,17'd27393,17'd27394,17'd27395,17'd27396,17'd27397,17'd27398,17'd27399,17'd27400,17'd27401,17'd19449,17'd18605,17'd27402,17'd27403,17'd19681,17'd27404,17'd27405,17'd27406,17'd27407,17'd27408,17'd27409,17'd27410,17'd27411,17'd19547,17'd27412,17'd27413,17'd27414,17'd27415,17'd27416,17'd27417,17'd27418,17'd27419,17'd22725,17'd27420,17'd27421,17'd27422,17'd21299,17'd26580,17'd21608,17'd21451,17'd25481,17'd21766,17'd12281,17'd27423,17'd27424,17'd23458,17'd7165,17'd27425,17'd27426,17'd5611,17'd6388,17'd6706,17'd10237,17'd6852,17'd6852,17'd9090,17'd8154,17'd10777,17'd11576,17'd10641,17'd10641,17'd9090,17'd6218,17'd6388,17'd5331,17'd5611,17'd5611,17'd5330,17'd5333,17'd26949,17'd5615,17'd5919,17'd9090,17'd26219,17'd14049,17'd16123,17'd15094,17'd15094,17'd15094,17'd15476,17'd22420,17'd22420,17'd17904,17'd18852,17'd27427,17'd12308,17'd27428,17'd27083,17'd27308,17'd23981,17'd25228,17'd27429,17'd12766,17'd26832,17'd27430,17'd27431,17'd27432,17'd27433,17'd27434,17'd27435,17'd27436,17'd27437,17'd27438,17'd27439,17'd1958,17'd1667,17'd2589,17'd27318,17'd2100,17'd2244,17'd2397,17'd2563,17'd26722,17'd26723,17'd27319,17'd27320,17'd27319,17'd27208,17'd26725,17'd26725,17'd25895,17'd25644,17'd24171,17'd23993,17'd24501,17'd24174,17'd5638,17'd24168,17'd5637,17'd5780,17'd24824,17'd23995,17'd27096,17'd24167,17'd17293,17'd3400,17'd4404,17'd4408,17'd3234,17'd26844,17'd21326,17'd27440,17'd3239,17'd9942,17'd257,17'd256,17'd459,17'd1271
},
'{
17'd27441,17'd4088,17'd4577,17'd7545,17'd2594,17'd2595,17'd3430,17'd12,17'd13,17'd13,17'd466,17'd4247,17'd17917,17'd10535,17'd2422,17'd1688,17'd27442,17'd26344,17'd4089,17'd18,17'd1128,17'd1128,17'd1128,17'd20404,17'd1128,17'd18,17'd652,17'd652,17'd980,17'd980,17'd27443,17'd27443,17'd27444,17'd6745,17'd6437,17'd6437,17'd5803,17'd27445,17'd27210,17'd5978,17'd27446,17'd27447,17'd27448,17'd27449,17'd26975,17'd6754,17'd27450,17'd27323,17'd27451,17'd27452,17'd2799,17'd27325,17'd22791,17'd27453,17'd27454,17'd18766,17'd26983,17'd18288,17'd27455,17'd17679,17'd27456,17'd27457,17'd21963,17'd12362,17'd27458,17'd12362,17'd20885,17'd12531,17'd20423,17'd17941,17'd16766,17'd17318,17'd17318,17'd15766,17'd16169,17'd24520,17'd17322,17'd15524,17'd24192,17'd17810,17'd27459,17'd27460,17'd27461,17'd19007,17'd17205,17'd18174,17'd17206,17'd17206,17'd21185,17'd19256,17'd16028,17'd13972,17'd9007,17'd4611,17'd5253,17'd25396,17'd27462,17'd27463,17'd7264,17'd26023,17'd9316,17'd27464,17'd15918,17'd27465,17'd26987,17'd10437,17'd11769,17'd27330,17'd27466,17'd27467,17'd27332,17'd27468,17'd27469,17'd27470,17'd26993,17'd27471,17'd27472,17'd27473,17'd27474,17'd27475,17'd27476,17'd11953,17'd27477,17'd25406,17'd12102,17'd12101,17'd27478,17'd26624,17'd13998,17'd27479,17'd10969,17'd27480,17'd27481,17'd27482,17'd16549,17'd9620,17'd9480,17'd10743,17'd16796,17'd11133,17'd14931,17'd13762,17'd15185,17'd15053,17'd12579,17'd15434,17'd12418,17'd13252,17'd13252,17'd12418,17'd18200,17'd24991,17'd26872,17'd27483,17'd25526,17'd26756,17'd24705,17'd24030,17'd18084,17'd27484,17'd27485,17'd27486,17'd12108,17'd18198,17'd16442,17'd18327,17'd16326,17'd19158,17'd13883,17'd11806,17'd11962,17'd18560,17'd14132,17'd27487,17'd10331,17'd27488,17'd21205,17'd11132,17'd11808,17'd11964,17'd13645,17'd11965,17'd10990,17'd11132,17'd19282,17'd13886,17'd15182,17'd15805,17'd15182,17'd10476,17'd17847,17'd17965,17'd27489,17'd22813,17'd15944,17'd22814,17'd16549,17'd11276,17'd16687,17'd17343,17'd23513,17'd16325,17'd13646,17'd11961,17'd12861,17'd12861,17'd11806,17'd12420,17'd12110,17'd13365,17'd12419,17'd12577,17'd13882,17'd13646,17'd11396,17'd11274,17'd11131,17'd10326,17'd10606,17'd22296,17'd10472,17'd10473,17'd10990,17'd11519,17'd11665,17'd11665,17'd14673,17'd25280,17'd11398,17'd11399,17'd11133,17'd10479,17'd27490,17'd27491,17'd27492,17'd27493,17'd27494,17'd27495,17'd27496,17'd27497,17'd27498,17'd27499,17'd27500,17'd27501,17'd27502,17'd27503,17'd27504,17'd27505,17'd27506,17'd27507,17'd25168,17'd24402,17'd24402,17'd25023,17'd24578,17'd25169,17'd25826,17'd27508,17'd27508,17'd25826,17'd26277,17'd26652,17'd26780,17'd25558,17'd25558,17'd26523,17'd26652,17'd26277,17'd26523,17'd26652,17'd26897,17'd26522,17'd26276,17'd26523,17'd25558,17'd25429,17'd25948,17'd24242,17'd27509,17'd27510,17'd27511,17'd27512,17'd25568,17'd25709,17'd27513,17'd26174,17'd27514,17'd27515,17'd25948,17'd25311,17'd26400,17'd26400,17'd26279,17'd26279,17'd26279,17'd26279,17'd26279,17'd25311,17'd25312,17'd27145,17'd25554,17'd26524,17'd25557,17'd27368,17'd27516,17'd27517,17'd27518,17'd27519,17'd27520,17'd27521,17'd27522,17'd27153,17'd27268,17'd27523,17'd26790,17'd26909,17'd27524,17'd27525,17'd27526,17'd27527,17'd27528,17'd26675,17'd27529,17'd27386,17'd27530,17'd27531,17'd26551,17'd27532,17'd27533,17'd27534,17'd27535,17'd26081,17'd27536,17'd27537,17'd27538,17'd27539,17'd27540,17'd27541,17'd27174,17'd20352,17'd27542,17'd27543,17'd27544,17'd27545,17'd27546,17'd27546,17'd18014,17'd19449,17'd27547,17'd19461,17'd24129,17'd27548,17'd27549,17'd27550,17'd27551,17'd27552,17'd27553,17'd27554,17'd27555,17'd27556,17'd27557,17'd27558,17'd27559,17'd27560,17'd27561,17'd27562,17'd27563,17'd27564,17'd27565,17'd26948,17'd27566,17'd21451,17'd21924,17'd27567,17'd21142,17'd12281,17'd27568,17'd22245,17'd7166,17'd6548,17'd27569,17'd5613,17'd26451,17'd6706,17'd6852,17'd26219,17'd26219,17'd8154,17'd8154,17'd9394,17'd10641,17'd10641,17'd12160,17'd8780,17'd9091,17'd6390,17'd5335,17'd5330,17'd27570,17'd27570,17'd5334,17'd27571,17'd27081,17'd26949,17'd6553,17'd12466,17'd14049,17'd14301,17'd27198,17'd17535,17'd14971,17'd17655,17'd22420,17'd22420,17'd15476,17'd18375,17'd18971,17'd22944,17'd15856,17'd25088,17'd18622,17'd27572,17'd26454,17'd20548,17'd17287,17'd27573,17'd25775,17'd24660,17'd19352,17'd25490,17'd27574,17'd27575,17'd27576,17'd27577,17'd27578,17'd27579,17'd610,17'd952,17'd602,17'd25374,17'd27580,17'd27581,17'd12645,17'd14979,17'd27582,17'd26840,17'd27319,17'd27583,17'd27320,17'd27320,17'd26723,17'd26725,17'd26842,17'd26842,17'd27584,17'd27585,17'd23994,17'd26843,17'd5637,17'd5637,17'd5637,17'd5780,17'd23995,17'd23995,17'd27586,17'd27587,17'd16257,17'd3401,17'd3402,17'd27588,17'd27589,17'd4074,17'd3885,17'd27440,17'd10389,17'd458,17'd268,17'd459,17'd460,17'd456
},
'{
17'd27590,17'd4088,17'd27591,17'd7545,17'd1831,17'd4247,17'd466,17'd13,17'd13,17'd466,17'd1127,17'd2594,17'd10535,17'd10535,17'd2422,17'd1688,17'd27442,17'd26344,17'd3905,17'd18,17'd1128,17'd1128,17'd1128,17'd1128,17'd18,17'd18,17'd652,17'd652,17'd980,17'd980,17'd27443,17'd27443,17'd6745,17'd6745,17'd6437,17'd6437,17'd6746,17'd11211,17'd27592,17'd6442,17'd27593,17'd27447,17'd27594,17'd27595,17'd26975,17'd6754,17'd26736,17'd26977,17'd3606,17'd3272,17'd27596,17'd23661,17'd27102,17'd27597,17'd27598,17'd18525,17'd18646,17'd26850,17'd27599,17'd27600,17'd27456,17'd23151,17'd14470,17'd13094,17'd24347,17'd12362,17'd12531,17'd12532,17'd17941,17'd16766,17'd16410,17'd16289,17'd16880,17'd15899,17'd16169,17'd16169,17'd16769,17'd15902,17'd16768,17'd17810,17'd27460,17'd27601,17'd18774,17'd18774,17'd17205,17'd17205,17'd17206,17'd21185,17'd18060,17'd16028,17'd23837,17'd14769,17'd8539,17'd4926,17'd6138,17'd24976,17'd27602,17'd13612,17'd7923,17'd27603,17'd9449,17'd25660,17'd15918,17'd15918,17'd15405,17'd27604,17'd12223,17'd27605,17'd27606,17'd27607,17'd27332,17'd27468,17'd27608,17'd27609,17'd27610,17'd27611,17'd27612,17'd27613,17'd26620,17'd27614,17'd17465,17'd11802,17'd16062,17'd25140,17'd27615,17'd27616,17'd12100,17'd27478,17'd26367,17'd27617,17'd27618,17'd27619,17'd27620,17'd14928,17'd9479,17'd16328,17'd9345,17'd10743,17'd17719,17'd10475,17'd14262,17'd13762,17'd12996,17'd13883,17'd12579,17'd12108,17'd12417,17'd13252,17'd12417,17'd12860,17'd18083,17'd26872,17'd27621,17'd27483,17'd27622,17'd26756,17'd23512,17'd24537,17'd26758,17'd27349,17'd27349,17'd18200,17'd11959,17'd15053,17'd19158,17'd11522,17'd19158,17'd16442,17'd11960,17'd13883,17'd13362,17'd20910,17'd26374,17'd26152,17'd12585,17'd27488,17'd26037,17'd10476,17'd11274,17'd11964,17'd13516,17'd11129,17'd11131,17'd19282,17'd10476,17'd12720,17'd21986,17'd15432,17'd24860,17'd12863,17'd17965,17'd22812,17'd9190,17'd10335,17'd14674,17'd11809,17'd11276,17'd12721,17'd11521,17'd19920,17'd21361,17'd18198,17'd11960,17'd13363,17'd13363,17'd13363,17'd13761,17'd12109,17'd16321,17'd12578,17'd13514,17'd13882,17'd13646,17'd11521,17'd11398,17'd27623,17'd19532,17'd10991,17'd17720,17'd17124,17'd27236,17'd24860,17'd15047,17'd16435,17'd21982,17'd16435,17'd11522,17'd13367,17'd23337,17'd11398,17'd10991,17'd10479,17'd19531,17'd27006,17'd27492,17'd27624,17'd27625,17'd27626,17'd27627,17'd27496,17'd27628,17'd27629,17'd27630,17'd27631,17'd27502,17'd27632,17'd27633,17'd27505,17'd27634,17'd26166,17'd25307,17'd24402,17'd25023,17'd25023,17'd24578,17'd25308,17'd25310,17'd27635,17'd25551,17'd25308,17'd27636,17'd26652,17'd25555,17'd25554,17'd25558,17'd26523,17'd26652,17'd26652,17'd26523,17'd26523,17'd26897,17'd26522,17'd26522,17'd26652,17'd25554,17'd26400,17'd25699,17'd23553,17'd23726,17'd24412,17'd27637,17'd25178,17'd25178,17'd27512,17'd27638,17'd25949,17'd27639,17'd27640,17'd25312,17'd25311,17'd26279,17'd26279,17'd26279,17'd26279,17'd26279,17'd26279,17'd26279,17'd25429,17'd25429,17'd27641,17'd25554,17'd26525,17'd25555,17'd27642,17'd27643,17'd27644,17'd27645,17'd27646,17'd27647,17'd27648,17'd27649,17'd27650,17'd27268,17'd27523,17'd27651,17'd27652,17'd27653,17'd27654,17'd27526,17'd27655,17'd27656,17'd27657,17'd27658,17'd27659,17'd27660,17'd27661,17'd27163,17'd27662,17'd27045,17'd27663,17'd26296,17'd27664,17'd27665,17'd27666,17'd24925,17'd27667,17'd21558,17'd27668,17'd27669,17'd17265,17'd27670,17'd27671,17'd17769,17'd17772,17'd18727,17'd27672,17'd18014,17'd27673,17'd25605,17'd19580,17'd20220,17'd27674,17'd27675,17'd27676,17'd27677,17'd27678,17'd27679,17'd27680,17'd27681,17'd27682,17'd27683,17'd27684,17'd27685,17'd27686,17'd21277,17'd22382,17'd27687,17'd27688,17'd23613,17'd27689,17'd27566,17'd27690,17'd25481,17'd27691,17'd27692,17'd27693,17'd27694,17'd10499,17'd9219,17'd6844,17'd27695,17'd5613,17'd5482,17'd6706,17'd9394,17'd10513,17'd10777,17'd10513,17'd9090,17'd9657,17'd10777,17'd11181,17'd11037,17'd10515,17'd27696,17'd9091,17'd5614,17'd5160,17'd27697,17'd27697,17'd5330,17'd5333,17'd26828,17'd5762,17'd6218,17'd24652,17'd12465,17'd12760,17'd14423,17'd27198,17'd14971,17'd17655,17'd17904,17'd22420,17'd15476,17'd15476,17'd20115,17'd22944,17'd15856,17'd18972,17'd18622,17'd17906,17'd26454,17'd20548,17'd27698,17'd13415,17'd27699,17'd26331,17'd17072,17'd27700,17'd27701,17'd27702,17'd27703,17'd27704,17'd27705,17'd27706,17'd403,17'd1098,17'd602,17'd26965,17'd27707,17'd27708,17'd27709,17'd14979,17'd24668,17'd26840,17'd27710,17'd27711,17'd27320,17'd27320,17'd26723,17'd26968,17'd26725,17'd26842,17'd26598,17'd27585,17'd24501,17'd26843,17'd5637,17'd5637,17'd5637,17'd5780,17'd23995,17'd24174,17'd27586,17'd27587,17'd16257,17'd3401,17'd3402,17'd2105,17'd3728,17'd4074,17'd3885,17'd27712,17'd10389,17'd458,17'd257,17'd265,17'd456,17'd254
},
'{
17'd27713,17'd4733,17'd4577,17'd5508,17'd1831,17'd4247,17'd2595,17'd466,17'd466,17'd466,17'd4247,17'd2594,17'd27714,17'd27714,17'd1831,17'd4247,17'd22965,17'd26344,17'd3905,17'd18,17'd1128,17'd1128,17'd1128,17'd1128,17'd18,17'd18,17'd652,17'd652,17'd980,17'd980,17'd27443,17'd20570,17'd6745,17'd6745,17'd6437,17'd6903,17'd6439,17'd10672,17'd6112,17'd6442,17'd27715,17'd27716,17'd27594,17'd27595,17'd26975,17'd26239,17'd27323,17'd24002,17'd3606,17'd3272,17'd2622,17'd23661,17'd27717,17'd26849,17'd4108,17'd25255,17'd15125,17'd26850,17'd27718,17'd27719,17'd26853,17'd23151,17'd14470,17'd13094,17'd12815,17'd12362,17'd12532,17'd20423,17'd17941,17'd17205,17'd17318,17'd16289,17'd16880,17'd16034,17'd16169,17'd15902,17'd18776,17'd17810,17'd17810,17'd19257,17'd27461,17'd19128,17'd17689,17'd18774,17'd18174,17'd17205,17'd16410,17'd17318,17'd16164,17'd19256,17'd23501,17'd9704,17'd4611,17'd5253,17'd9842,17'd8694,17'd27463,17'd14640,17'd27220,17'd10295,17'd27720,17'd25660,17'd26987,17'd26987,17'd14642,17'd10819,17'd27721,17'd27722,17'd27723,17'd27607,17'd27724,17'd27608,17'd27725,17'd27726,17'd27727,17'd9327,17'd27728,17'd27729,17'd27730,17'd27731,17'd10839,17'd12248,17'd27732,17'd10983,17'd27733,17'd11386,17'd11952,17'd12100,17'd17465,17'd27734,17'd10723,17'd9879,17'd27735,17'd17011,17'd9344,17'd10173,17'd9480,17'd9885,17'd10329,17'd10990,17'd14262,17'd13362,17'd12858,17'd12419,17'd12579,17'd14807,17'd13517,17'd13517,17'd12415,17'd16558,17'd27736,17'd27737,17'd27004,17'd24857,17'd26756,17'd24031,17'd24537,17'd25528,17'd27348,17'd27349,17'd26758,17'd12254,17'd18198,17'd16204,17'd13762,17'd13762,17'd15185,17'd13520,17'd13366,17'd11667,17'd10853,17'd27738,17'd27739,17'd10165,17'd12863,17'd15176,17'd14134,17'd17236,17'd14810,17'd14810,17'd10736,17'd20910,17'd14263,17'd11131,17'd14931,17'd15182,17'd21986,17'd12720,17'd11133,17'd17719,17'd9620,17'd9481,17'd9743,17'd15187,17'd16549,17'd11671,17'd15176,17'd27740,17'd27741,17'd15055,17'd16203,17'd12579,17'd12109,17'd12110,17'd12577,17'd12414,17'd15434,17'd15434,17'd12579,17'd12414,17'd12577,17'd13363,17'd11807,17'd10990,17'd19282,17'd19532,17'd10991,17'd10328,17'd27742,17'd27743,17'd10853,17'd13885,17'd15679,17'd16797,17'd11666,17'd11666,17'd11962,17'd13520,17'd13762,17'd11274,17'd10991,17'd10479,17'd12116,17'd27744,17'd27745,17'd27746,17'd27747,17'd27748,17'd27749,17'd27355,17'd27750,17'd27751,17'd27752,17'd27753,17'd27754,17'd27755,17'd27756,17'd27757,17'd27758,17'd27759,17'd27760,17'd25307,17'd24399,17'd24402,17'd25169,17'd25169,17'd25551,17'd25551,17'd25169,17'd24578,17'd26652,17'd26652,17'd25555,17'd25554,17'd25558,17'd26780,17'd26652,17'd26652,17'd26523,17'd26523,17'd26276,17'd27761,17'd26277,17'd26523,17'd25698,17'd26167,17'd25700,17'd26061,17'd23725,17'd27762,17'd27763,17'd25180,17'd25178,17'd27764,17'd27765,17'd27766,17'd27767,17'd27514,17'd25948,17'd25312,17'd26279,17'd26279,17'd26279,17'd26279,17'd26279,17'd26279,17'd26167,17'd25429,17'd26279,17'd25429,17'd25554,17'd27368,17'd27768,17'd27642,17'd27769,17'd27770,17'd27771,17'd27772,17'd27519,17'd27773,17'd27774,17'd27775,17'd27776,17'd27037,17'd27651,17'd27777,17'd27778,17'd27779,17'd27780,17'd27781,17'd24755,17'd25334,17'd26414,17'd27658,17'd26410,17'd27782,17'd27783,17'd27532,17'd27784,17'd26297,17'd26296,17'd27664,17'd27785,17'd27786,17'd27787,17'd27788,17'd27789,17'd20645,17'd27790,17'd27174,17'd27791,17'd27792,17'd27793,17'd19680,17'd19199,17'd18841,17'd18735,17'd27794,17'd27795,17'd27796,17'd19689,17'd27797,17'd27798,17'd27799,17'd27800,17'd27801,17'd27802,17'd27803,17'd27804,17'd27805,17'd27806,17'd27807,17'd27808,17'd27809,17'd27810,17'd20826,17'd27811,17'd22558,17'd27812,17'd23786,17'd21765,17'd27690,17'd25481,17'd27691,17'd27813,17'd27814,17'd11159,17'd10766,17'd8913,17'd6846,17'd5915,17'd5613,17'd5481,17'd6387,17'd26219,17'd10513,17'd10777,17'd10777,17'd10513,17'd8304,17'd10513,17'd11181,17'd10642,17'd10642,17'd27815,17'd7668,17'd5919,17'd5335,17'd4845,17'd27570,17'd5330,17'd5334,17'd26949,17'd5336,17'd6389,17'd6852,17'd12466,17'd14048,17'd12622,17'd14423,17'd14970,17'd14971,17'd15476,17'd17904,17'd15476,17'd15476,17'd18500,17'd14051,17'd15856,17'd18972,17'd16373,17'd24153,17'd19851,17'd21456,17'd27698,17'd13171,17'd26955,17'd27816,17'd18137,17'd27817,17'd26332,17'd25637,17'd27818,17'd27819,17'd27820,17'd27821,17'd431,17'd1963,17'd1099,17'd5941,17'd27707,17'd27708,17'd27709,17'd2561,17'd24668,17'd26840,17'd27710,17'd27822,17'd27319,17'd27319,17'd26723,17'd26968,17'd26725,17'd26725,17'd26598,17'd23817,17'd24502,17'd26843,17'd26232,17'd26232,17'd5637,17'd5637,17'd26123,17'd24174,17'd27823,17'd27587,17'd16257,17'd15485,17'd4066,17'd27588,17'd27589,17'd4074,17'd3885,17'd20401,17'd3414,17'd409,17'd257,17'd265,17'd254,17'd27824
},
'{
17'd4243,17'd4733,17'd4887,17'd5508,17'd10535,17'd2594,17'd4247,17'd1127,17'd1127,17'd4247,17'd2594,17'd10535,17'd10535,17'd10535,17'd1831,17'd4247,17'd22965,17'd4089,17'd3905,17'd18,17'd1128,17'd1128,17'd1128,17'd1128,17'd18,17'd18,17'd652,17'd652,17'd980,17'd27,17'd20570,17'd20570,17'd7225,17'd6745,17'd6437,17'd6903,17'd10408,17'd7730,17'd6112,17'd6442,17'd27446,17'd27825,17'd27448,17'd27212,17'd26237,17'd27826,17'd4265,17'd27827,17'd27828,17'd2956,17'd27829,17'd27830,17'd27831,17'd26982,17'd18159,17'd15371,17'd26610,17'd15888,17'd27832,17'd26985,17'd26853,17'd23151,17'd14470,17'd13094,17'd12362,17'd12680,17'd12681,17'd19753,17'd16766,17'd16986,17'd17319,17'd18060,17'd16659,17'd16169,17'd16033,17'd15524,17'd17448,17'd17810,17'd17448,17'd27833,17'd27834,17'd20148,17'd17689,17'd18655,17'd18174,17'd17205,17'd16410,17'd17319,17'd19256,17'd16028,17'd13844,17'd9704,17'd7088,17'd6138,17'd8381,17'd8383,17'd27835,17'd12371,17'd27836,17'd10294,17'd27837,17'd26483,17'd15917,17'd25132,17'd27221,17'd27838,17'd27839,17'd27840,17'd27841,17'd27842,17'd25918,17'd27843,17'd27844,17'd27845,17'd27846,17'd27847,17'd27848,17'd27849,17'd10833,17'd27850,17'd27851,17'd11124,17'd27852,17'd11955,17'd27733,17'd11386,17'd10840,17'd10840,17'd27853,17'd10837,17'd10592,17'd27854,17'd27855,17'd27856,17'd9346,17'd10173,17'd9620,17'd9885,17'd11670,17'd14931,17'd11807,17'd11963,17'd12113,17'd12577,17'd12414,17'd14807,17'd13515,17'd14003,17'd16913,17'd26758,17'd26629,17'd26872,17'd24857,17'd25526,17'd24705,17'd24538,17'd25927,17'd26757,17'd27857,17'd27858,17'd23855,17'd14807,17'd18197,17'd16204,17'd13362,17'd11807,17'd13646,17'd13366,17'd13764,17'd11395,17'd27859,17'd27236,17'd10023,17'd10326,17'd15176,17'd14134,17'd11524,17'd13138,17'd14810,17'd14931,17'd14931,17'd25144,17'd14132,17'd10990,17'd12720,17'd13137,17'd13000,17'd13886,17'd9883,17'd10743,17'd12117,17'd9189,17'd9345,17'd9741,17'd12585,17'd12423,17'd17343,17'd27860,17'd27861,17'd23168,17'd19283,17'd19032,17'd15434,17'd15434,17'd19032,17'd19032,17'd16685,17'd18564,17'd27862,17'd14130,17'd11806,17'd11667,17'd14810,17'd16555,17'd11133,17'd14518,17'd10165,17'd27863,17'd27864,17'd12862,17'd18078,17'd13764,17'd11962,17'd20313,17'd13253,17'd13253,17'd12113,17'd12858,17'd11963,17'd10989,17'd10991,17'd10479,17'd11277,17'd10172,17'd27865,17'd27866,17'd27867,17'd27868,17'd27354,17'd27869,17'd27870,17'd27871,17'd27872,17'd27753,17'd27873,17'd27874,17'd27875,17'd27876,17'd27758,17'd27877,17'd27878,17'd25168,17'd24398,17'd24402,17'd25169,17'd25308,17'd26054,17'd25551,17'd24578,17'd25428,17'd26652,17'd26652,17'd25555,17'd25554,17'd25554,17'd26780,17'd26652,17'd26780,17'd25558,17'd25558,17'd26278,17'd27768,17'd26523,17'd25558,17'd25944,17'd26167,17'd25700,17'd27879,17'd24243,17'd27880,17'd27881,17'd24417,17'd25030,17'd27764,17'd27882,17'd25566,17'd26062,17'd27883,17'd25313,17'd25312,17'd25429,17'd26279,17'd26279,17'd26279,17'd26279,17'd26279,17'd25696,17'd26279,17'd26279,17'd26394,17'd25698,17'd27768,17'd27884,17'd26277,17'd27885,17'd27886,17'd27887,17'd27888,17'd27889,17'd27890,17'd27891,17'd27775,17'd27892,17'd27893,17'd26539,17'd27894,17'd27895,17'd24601,17'd27896,17'd27897,17'd27898,17'd25453,17'd27899,17'd25849,17'd26304,17'd27660,17'd27900,17'd27532,17'd27901,17'd27902,17'd27903,17'd27275,17'd27904,17'd27905,17'd24273,17'd25723,17'd27906,17'd27907,17'd27908,17'd27909,17'd18723,17'd27910,17'd27400,17'd27911,17'd27673,17'd25214,17'd18735,17'd18605,17'd27404,17'd27912,17'd19689,17'd27797,17'd27913,17'd27914,17'd27915,17'd27916,17'd27917,17'd27918,17'd27919,17'd27920,17'd27921,17'd27922,17'd27296,17'd27923,17'd27924,17'd20670,17'd27925,17'd27926,17'd27927,17'd23444,17'd22080,17'd27690,17'd25481,17'd27691,17'd27813,17'd27928,17'd12281,17'd11549,17'd27929,17'd7169,17'd6214,17'd27930,17'd5915,17'd5332,17'd9394,17'd10513,17'd10777,17'd10777,17'd10513,17'd9657,17'd27931,17'd27932,17'd27933,17'd27934,17'd10642,17'd8780,17'd6391,17'd27935,17'd5002,17'd5329,17'd5329,17'd5330,17'd5762,17'd5336,17'd6389,17'd6707,17'd9394,17'd25226,17'd14301,17'd16123,17'd13925,17'd14971,17'd15340,17'd17904,17'd15476,17'd15340,17'd18500,17'd14051,17'd27936,17'd18972,17'd27937,17'd25227,17'd25485,17'd25089,17'd27938,17'd27939,17'd27940,17'd27941,17'd18137,17'd27942,17'd27943,17'd27944,17'd27818,17'd27945,17'd27946,17'd27947,17'd27948,17'd641,17'd1668,17'd1383,17'd27949,17'd27708,17'd27709,17'd2561,17'd24668,17'd26840,17'd27319,17'd27822,17'd27319,17'd27319,17'd26723,17'd26968,17'd26725,17'd26725,17'd26598,17'd23992,17'd24670,17'd27096,17'd26232,17'd26232,17'd26232,17'd5637,17'd26123,17'd23481,17'd24167,17'd27950,17'd17418,17'd3229,17'd3403,17'd2106,17'd3580,17'd3885,17'd3730,17'd20401,17'd3239,17'd409,17'd257,17'd2255,17'd254,17'd27824
},
'{
17'd27951,17'd4733,17'd4246,17'd13428,17'd7372,17'd7214,17'd1688,17'd1127,17'd4247,17'd1688,17'd1831,17'd10535,17'd10535,17'd10535,17'd1831,17'd4247,17'd22965,17'd1416,17'd3905,17'd3905,17'd1128,17'd1128,17'd1128,17'd1128,17'd3905,17'd18,17'd652,17'd652,17'd7060,17'd7060,17'd20570,17'd20570,17'd7387,17'd7387,17'd7062,17'd6599,17'd10672,17'd7730,17'd6112,17'd6442,17'd5813,17'd27825,17'd27952,17'd11456,17'd26238,17'd27953,17'd27954,17'd27955,17'd27828,17'd2956,17'd27956,17'd27957,17'd27103,17'd26133,17'd27958,17'd25392,17'd27959,17'd27960,17'd27719,17'd27456,17'd27457,17'd22117,17'd14470,17'd13094,17'd11913,17'd12680,17'd12681,17'd19753,17'd16766,17'd16986,17'd17319,17'd19256,17'd16519,17'd17942,17'd17810,17'd18534,17'd17690,17'd17690,17'd19011,17'd19255,17'd27961,17'd20148,17'd17689,17'd18655,17'd18174,17'd17205,17'd17318,17'd17319,17'd16659,17'd16659,17'd13469,17'd9704,17'd4926,17'd6304,17'd8543,17'd8384,17'd27962,17'd8702,17'd27836,17'd10129,17'd16180,17'd26483,17'd15917,17'd15786,17'd14905,17'd27963,17'd27964,17'd27965,17'd27966,17'd27842,17'd27967,17'd27968,17'd27969,17'd27970,17'd27971,17'd27972,17'd27973,17'd27339,17'd27974,17'd27975,17'd27976,17'd27977,17'd27978,17'd27979,17'd27733,17'd27980,17'd10726,17'd10318,17'd27618,17'd27981,17'd9874,17'd27982,17'd27983,17'd13887,17'd10174,17'd15807,17'd9620,17'd16796,17'd11132,17'd14673,17'd11807,17'd13135,17'd12111,17'd12413,17'd12109,17'd17348,17'd19407,17'd23681,17'd27121,17'd26629,17'd27121,17'd27004,17'd25526,17'd24705,17'd24705,17'd26493,17'd26757,17'd27984,17'd27857,17'd27737,17'd12108,17'd11959,17'd18917,17'd12422,17'd11963,17'd12861,17'd20313,17'd13764,17'd11666,17'd10990,17'd26374,17'd15300,17'd10023,17'd10606,17'd14518,17'd11399,17'd11274,17'd16068,17'd17236,17'd16320,17'd10739,17'd16555,17'd25144,17'd10736,17'd13885,17'd13000,17'd13138,17'd11527,17'd9741,17'd9339,17'd8873,17'd16318,17'd16554,17'd17719,17'd12423,17'd24540,17'd27985,17'd26149,17'd24856,17'd23511,17'd18083,17'd16559,17'd12860,17'd16559,17'd16559,17'd17727,17'd16558,17'd18200,17'd25670,17'd27986,17'd13520,17'd11808,17'd16555,17'd27002,17'd17720,17'd10164,17'd27987,17'd16555,17'd11520,17'd15175,17'd11961,17'd13135,17'd12858,17'd13363,17'd13366,17'd11961,17'd12259,17'd14002,17'd18447,17'd18560,17'd10603,17'd15688,17'd15048,17'd22812,17'd27988,17'd27989,17'd27990,17'd27991,17'd27992,17'd27993,17'd27994,17'd27995,17'd27996,17'd27997,17'd27998,17'd27999,17'd28000,17'd28001,17'd28002,17'd28003,17'd28004,17'd25548,17'd24396,17'd24402,17'd25825,17'd25825,17'd27508,17'd25551,17'd24578,17'd24578,17'd26652,17'd26652,17'd26780,17'd25558,17'd25554,17'd25558,17'd26523,17'd26780,17'd26167,17'd26167,17'd25553,17'd26524,17'd25558,17'd26524,17'd25698,17'd26279,17'd25703,17'd28005,17'd26061,17'd28006,17'd28007,17'd28008,17'd24898,17'd27637,17'd25177,17'd25435,17'd26174,17'd28009,17'd25430,17'd25313,17'd25311,17'd26400,17'd26167,17'd26167,17'd26167,17'd26167,17'd25696,17'd26167,17'd25944,17'd26394,17'd26394,17'd26278,17'd28010,17'd27761,17'd27885,17'd28011,17'd28012,17'd28013,17'd28014,17'd28015,17'd26409,17'd28016,17'd28017,17'd27034,17'd28018,17'd27038,17'd28019,17'd25453,17'd28020,17'd28021,17'd28022,17'd27033,17'd25188,17'd25586,17'd28023,17'd26669,17'd28024,17'd26677,17'd28025,17'd28026,17'd28027,17'd27275,17'd28028,17'd28024,17'd25056,17'd24433,17'd28029,17'd25855,17'd26422,17'd28030,17'd28031,17'd28032,17'd28033,17'd28034,17'd27911,17'd27673,17'd18014,17'd19816,17'd25608,17'd28035,17'd28036,17'd28037,17'd28038,17'd28039,17'd28040,17'd28041,17'd28042,17'd28043,17'd28044,17'd28045,17'd28046,17'd28047,17'd28048,17'd28049,17'd28050,17'd28051,17'd28052,17'd28053,17'd28054,17'd23266,17'd28055,17'd22081,17'd21923,17'd25481,17'd24640,17'd27928,17'd26447,17'd27423,17'd22245,17'd8145,17'd6213,17'd6552,17'd6552,17'd28056,17'd8154,17'd10513,17'd10777,17'd10513,17'd9657,17'd10513,17'd10897,17'd27931,17'd27933,17'd28057,17'd11037,17'd10514,17'd28058,17'd5614,17'd5004,17'd5002,17'd5002,17'd5329,17'd5333,17'd5336,17'd27935,17'd5615,17'd9090,17'd12465,17'd12760,17'd12622,17'd13925,17'd14970,17'd17655,17'd15476,17'd15340,17'd15340,17'd28059,17'd14424,17'd15611,17'd16126,17'd16489,17'd25227,17'd23288,17'd26114,17'd20852,17'd25486,17'd27940,17'd25775,17'd22598,17'd25887,17'd28060,17'd28061,17'd28062,17'd28063,17'd26593,17'd28064,17'd28065,17'd772,17'd191,17'd2098,17'd28066,17'd27708,17'd27709,17'd2561,17'd24668,17'd26725,17'd27319,17'd27320,17'd27319,17'd27319,17'd26723,17'd26723,17'd26725,17'd26725,17'd26598,17'd23817,17'd28067,17'd28068,17'd5638,17'd5638,17'd23133,17'd23133,17'd23481,17'd24329,17'd27587,17'd28069,17'd15865,17'd14980,17'd4066,17'd12775,17'd28070,17'd3885,17'd3730,17'd3236,17'd3239,17'd409,17'd1242,17'd254,17'd27824,17'd182
},
'{
17'd27951,17'd4245,17'd14743,17'd15746,17'd13428,17'd7545,17'd3250,17'd2781,17'd3250,17'd3250,17'd2422,17'd3252,17'd3252,17'd1831,17'd1688,17'd4247,17'd1416,17'd1416,17'd3905,17'd3905,17'd1128,17'd1128,17'd1128,17'd1128,17'd3905,17'd3905,17'd652,17'd652,17'd7060,17'd7060,17'd20570,17'd20570,17'd7387,17'd7387,17'd7062,17'd6599,17'd10672,17'd10672,17'd6112,17'd6442,17'd5813,17'd28071,17'd26734,17'd28072,17'd28073,17'd5390,17'd28074,17'd28075,17'd28076,17'd2956,17'd28077,17'd14753,17'd21480,17'd20728,17'd26479,17'd25392,17'd28078,17'd27960,17'd28079,17'd26612,17'd26353,17'd22117,17'd14470,17'd12362,17'd11913,17'd11629,17'd17941,17'd17205,17'd16986,17'd21185,17'd16519,17'd17694,17'd18776,17'd17810,17'd17448,17'd18776,17'd17690,17'd17445,17'd24688,17'd19259,17'd20148,17'd20148,17'd17689,17'd18774,17'd17205,17'd17206,17'd16289,17'd20585,17'd16659,17'd13721,17'd9575,17'd4611,17'd5252,17'd8847,17'd28080,17'd8222,17'd7921,17'd8702,17'd27836,17'd9587,17'd16780,17'd16295,17'd25132,17'd28081,17'd28082,17'd28083,17'd28084,17'd28085,17'd27966,17'd28086,17'd28087,17'd28088,17'd28089,17'd28090,17'd28091,17'd9722,17'd28092,17'd28093,17'd28094,17'd28095,17'd28096,17'd28097,17'd28098,17'd28099,17'd28100,17'd10464,17'd10155,17'd28101,17'd10722,17'd9874,17'd27982,17'd28102,17'd25281,17'd13887,17'd10174,17'd9344,17'd10992,17'd10330,17'd11524,17'd13762,17'd13135,17'd11961,17'd12718,17'd12577,17'd16321,17'd17348,17'd20452,17'd24704,17'd28103,17'd28104,17'd26370,17'd24537,17'd24705,17'd24031,17'd26493,17'd28105,17'd27984,17'd28106,17'd28104,17'd28107,17'd19408,17'd13883,17'd16204,17'd16204,17'd11957,17'd12112,17'd20313,17'd16064,17'd14810,17'd19282,17'd17124,17'd10023,17'd10164,17'd14518,17'd13886,17'd14931,17'd16068,17'd14673,17'd11524,17'd10476,17'd10991,17'd10475,17'd10737,17'd11666,17'd28108,17'd16068,17'd14134,17'd11276,17'd9620,17'd9043,17'd8873,17'd15180,17'd10856,17'd24996,17'd12583,17'd28109,17'd28110,17'd26370,17'd27121,17'd26629,17'd26373,17'd17727,17'd17727,17'd17971,17'd17971,17'd17846,17'd26373,17'd18084,17'd28111,17'd28112,17'd11397,17'd10854,17'd10855,17'd25811,17'd10023,17'd10023,17'd16320,17'd12862,17'd13253,17'd13520,17'd13883,17'd11960,17'd12420,17'd12419,17'd13761,17'd11961,17'd11958,17'd14002,17'd18447,17'd18560,17'd10740,17'd15688,17'd11809,17'd16552,17'd28113,17'd28114,17'd28115,17'd28116,17'd28117,17'd28118,17'd28119,17'd28120,17'd28121,17'd28122,17'd27998,17'd28123,17'd28124,17'd28125,17'd28002,17'd27877,17'd28126,17'd24888,17'd24396,17'd24889,17'd26053,17'd25825,17'd25551,17'd25826,17'd24578,17'd24578,17'd26277,17'd26652,17'd25555,17'd26524,17'd25554,17'd25558,17'd26523,17'd25555,17'd26400,17'd25702,17'd25311,17'd26400,17'd25559,17'd25553,17'd25696,17'd25311,17'd25431,17'd28127,17'd28005,17'd24244,17'd28128,17'd28129,17'd24895,17'd25179,17'd27637,17'd28130,17'd25833,17'd28131,17'd28132,17'd25313,17'd25311,17'd26400,17'd26167,17'd26167,17'd26167,17'd26167,17'd25553,17'd25696,17'd25698,17'd25944,17'd25557,17'd26523,17'd28010,17'd28133,17'd28134,17'd28135,17'd28136,17'd28137,17'd28138,17'd28139,17'd28140,17'd28141,17'd28017,17'd27378,17'd28018,17'd26670,17'd28142,17'd25189,17'd28143,17'd28144,17'd28145,17'd28146,17'd25042,17'd28147,17'd28148,17'd28149,17'd27661,17'd26919,17'd28150,17'd28151,17'd26913,17'd26792,17'd28152,17'd27533,17'd25199,17'd28153,17'd24761,17'd28154,17'd28155,17'd28156,17'd28157,17'd28158,17'd28159,17'd27543,17'd27793,17'd28160,17'd19328,17'd19710,17'd26688,17'd28161,17'd28162,17'd28163,17'd28164,17'd28165,17'd28166,17'd28167,17'd28168,17'd28169,17'd28170,17'd28171,17'd28172,17'd28173,17'd28174,17'd28175,17'd28176,17'd28177,17'd28178,17'd21742,17'd28179,17'd28180,17'd23615,17'd28181,17'd24638,17'd25481,17'd24640,17'd24640,17'd27928,17'd12444,17'd10361,17'd7990,17'd6213,17'd7667,17'd5918,17'd28182,17'd26709,17'd9657,17'd10777,17'd10513,17'd9657,17'd10777,17'd10897,17'd27931,17'd27933,17'd28183,17'd11037,17'd10642,17'd28184,17'd6219,17'd28185,17'd5004,17'd5002,17'd5005,17'd5334,17'd5335,17'd27935,17'd5615,17'd8154,17'd12466,17'd11854,17'd14301,17'd13558,17'd13925,17'd15094,17'd15476,17'd15340,17'd15340,17'd28186,17'd13167,17'd13801,17'd16126,17'd16489,17'd22090,17'd23288,17'd25363,17'd24315,17'd24946,17'd16253,17'd14579,17'd14056,17'd20257,17'd23469,17'd28187,17'd28188,17'd28189,17'd28190,17'd575,17'd28191,17'd771,17'd4084,17'd6721,17'd28066,17'd27708,17'd27709,17'd2243,17'd26967,17'd26725,17'd27320,17'd27320,17'd27319,17'd27319,17'd27209,17'd26723,17'd26725,17'd26725,17'd26598,17'd23817,17'd28192,17'd23480,17'd5638,17'd5638,17'd5638,17'd23133,17'd23481,17'd23307,17'd24325,17'd27950,17'd17418,17'd3229,17'd3716,17'd1954,17'd12638,17'd3730,17'd3581,17'd3236,17'd3239,17'd189,17'd801,17'd804,17'd182,17'd639
},
'{
17'd27951,17'd4245,17'd6420,17'd15876,17'd14743,17'd7545,17'd7545,17'd7711,17'd3250,17'd2784,17'd2935,17'd14070,17'd3252,17'd10535,17'd1831,17'd4247,17'd1416,17'd1416,17'd3905,17'd3905,17'd1128,17'd1128,17'd1128,17'd1128,17'd653,17'd653,17'd652,17'd28,17'd7060,17'd7060,17'd20570,17'd20570,17'd28193,17'd7387,17'd6599,17'd6904,17'd6441,17'd6441,17'd6112,17'd6442,17'd5813,17'd28071,17'd26734,17'd26237,17'd27826,17'd28194,17'd28195,17'd28075,17'd28196,17'd27596,17'd28197,17'd27717,17'd26849,17'd25907,17'd28198,17'd28199,17'd28200,17'd28201,17'd28202,17'd28203,17'd23151,17'd23836,17'd14470,17'd12361,17'd11764,17'd18412,17'd19753,17'd18174,17'd18656,17'd17319,17'd18060,17'd18534,17'd17810,17'd17692,17'd18776,17'd17448,17'd19130,17'd19008,17'd28204,17'd27961,17'd28205,17'd19382,17'd18774,17'd17689,17'd21649,17'd17206,17'd16289,17'd16880,17'd16880,17'd13469,17'd9007,17'd4767,17'd6304,17'd8380,17'd28206,17'd8222,17'd7923,17'd9167,17'd9447,17'd16997,17'd16781,17'd16046,17'd15785,17'd28207,17'd28208,17'd28209,17'd28210,17'd28211,17'd28212,17'd28213,17'd28087,17'd28214,17'd28215,17'd28216,17'd27972,17'd28217,17'd28218,17'd28219,17'd28220,17'd10155,17'd27732,17'd28221,17'd28222,17'd28099,17'd28223,17'd28224,17'd27618,17'd28225,17'd10314,17'd9733,17'd28226,17'd9476,17'd17964,17'd9039,17'd10174,17'd9346,17'd9885,17'd19282,17'd14673,17'd13762,17'd13135,17'd12419,17'd12718,17'd12419,17'd18198,17'd22819,17'd24537,17'd27004,17'd28103,17'd27737,17'd25927,17'd23512,17'd23515,17'd24537,17'd26370,17'd28227,17'd28228,17'd28229,17'd28230,17'd24033,17'd17722,17'd15185,17'd16204,17'd16204,17'd12858,17'd12112,17'd12861,17'd11520,17'd10475,17'd10166,17'd17719,17'd10479,17'd22296,17'd14518,17'd10990,17'd14673,17'd11522,17'd11274,17'd11524,17'd10476,17'd11132,17'd10739,17'd11395,17'd17598,17'd13885,17'd14931,17'd10330,17'd9742,17'd9743,17'd9043,17'd10174,17'd9478,17'd10741,17'd11274,17'd14260,17'd28231,17'd26370,17'd28103,17'd28104,17'd27349,17'd28232,17'd28233,17'd28234,17'd28234,17'd27349,17'd17846,17'd18083,17'd28235,17'd14260,17'd12583,17'd13521,17'd11399,17'd10991,17'd10166,17'd26374,17'd19156,17'd28236,17'd13885,17'd12996,17'd15053,17'd12419,17'd12109,17'd12995,17'd12856,17'd12419,17'd12420,17'd11960,17'd11806,17'd11963,17'd18445,17'd10325,17'd18196,17'd14674,17'd28237,17'd26633,17'd28238,17'd28238,17'd28239,17'd28240,17'd28241,17'd28242,17'd28243,17'd28244,17'd28245,17'd28246,17'd28247,17'd28000,17'd28248,17'd28249,17'd27759,17'd28250,17'd24732,17'd24396,17'd24574,17'd24402,17'd28251,17'd25826,17'd25826,17'd25169,17'd24578,17'd26652,17'd25697,17'd25555,17'd26524,17'd25554,17'd25558,17'd26523,17'd25554,17'd25948,17'd25431,17'd26285,17'd25562,17'd25831,17'd25702,17'd26055,17'd25312,17'd27514,17'd25707,17'd28252,17'd28253,17'd25029,17'd23562,17'd24416,17'd25031,17'd28254,17'd25317,17'd26174,17'd28131,17'd25704,17'd25172,17'd25312,17'd26400,17'd26167,17'd26167,17'd25698,17'd25698,17'd25558,17'd26524,17'd25554,17'd25558,17'd25555,17'd26780,17'd28255,17'd28256,17'd28257,17'd28258,17'd28259,17'd28260,17'd28261,17'd28262,17'd28263,17'd28264,17'd27035,17'd27379,17'd28265,17'd27663,17'd28266,17'd28267,17'd28268,17'd28269,17'd28270,17'd28022,17'd24910,17'd28271,17'd28272,17'd28023,17'd27162,17'd28273,17'd28274,17'd28275,17'd28276,17'd28277,17'd28278,17'd28152,17'd26542,17'd28279,17'd24437,17'd24912,17'd24273,17'd28280,17'd28281,17'd28282,17'd25612,17'd27793,17'd28283,17'd28284,17'd17517,17'd19569,17'd18014,17'd28285,17'd19465,17'd28286,17'd28287,17'd28288,17'd28289,17'd28290,17'd28291,17'd28292,17'd28293,17'd28294,17'd28295,17'd28296,17'd28297,17'd28298,17'd28299,17'd28300,17'd28301,17'd28302,17'd28303,17'd22576,17'd22407,17'd24139,17'd22241,17'd24638,17'd21923,17'd24640,17'd25622,17'd26582,17'd10766,17'd8913,17'd6845,17'd6214,17'd5918,17'd28304,17'd26709,17'd9090,17'd10777,17'd10777,17'd10777,17'd10513,17'd10897,17'd10897,17'd28305,17'd28306,17'd11709,17'd11709,17'd10777,17'd9090,17'd8303,17'd28307,17'd4842,17'd4686,17'd5330,17'd5334,17'd5335,17'd5614,17'd8303,17'd26219,17'd11853,17'd12467,17'd14301,17'd14301,17'd14971,17'd15340,17'd17655,17'd15094,17'd15727,17'd17535,17'd15611,17'd16126,17'd14426,17'd16251,17'd23981,17'd23804,17'd21005,17'd24946,17'd15099,17'd14579,17'd14056,17'd26116,17'd26715,17'd28308,17'd28309,17'd28310,17'd28311,17'd28312,17'd28313,17'd404,17'd410,17'd14178,17'd28314,17'd28315,17'd27581,17'd2243,17'd27095,17'd26722,17'd27320,17'd27320,17'd27319,17'd27319,17'd27319,17'd27320,17'd26968,17'd26968,17'd28316,17'd23817,17'd28192,17'd23480,17'd28317,17'd5638,17'd5638,17'd23133,17'd23133,17'd5945,17'd27587,17'd28069,17'd15865,17'd3229,17'd3716,17'd1675,17'd28318,17'd3728,17'd3581,17'd10389,17'd23301,17'd189,17'd255,17'd1123,17'd1683,17'd15492
},
'{
17'd25384,17'd4245,17'd6420,17'd27951,17'd6420,17'd4246,17'd4887,17'd4887,17'd2784,17'd2935,17'd3101,17'd3101,17'd14070,17'd3252,17'd1831,17'd4247,17'd1416,17'd1416,17'd3905,17'd3905,17'd1128,17'd1128,17'd1128,17'd1128,17'd653,17'd653,17'd652,17'd28,17'd7060,17'd7060,17'd20570,17'd20570,17'd28193,17'd7386,17'd6904,17'd6904,17'd6441,17'd28319,17'd6442,17'd5814,17'd5386,17'd5387,17'd6603,17'd28320,17'd4902,17'd28321,17'd28195,17'd27828,17'd28322,17'd2622,17'd27830,17'd28323,17'd28324,17'd4108,17'd18525,17'd15125,17'd28325,17'd28079,17'd26612,17'd28326,17'd22117,17'd25123,17'd16287,17'd16658,17'd11629,17'd18533,17'd17205,17'd17206,17'd17207,17'd16519,17'd17694,17'd18776,17'd18175,17'd18413,17'd18534,17'd17445,17'd19385,17'd18656,17'd27834,17'd23155,17'd20886,17'd19382,17'd18774,17'd19893,17'd21964,17'd16410,17'd16880,17'd15766,17'd13469,17'd9575,17'd4611,17'd5253,17'd8847,17'd8382,17'd8222,17'd8077,17'd7590,17'd9587,17'd16997,17'd16997,17'd16781,17'd16046,17'd15785,17'd28327,17'd28328,17'd28329,17'd28210,17'd28211,17'd28212,17'd28330,17'd27968,17'd28331,17'd28332,17'd28333,17'd28334,17'd28092,17'd28335,17'd28336,17'd28337,17'd11128,17'd27852,17'd28222,17'd28222,17'd27979,17'd11128,17'd28338,17'd28339,17'd28340,17'd28341,17'd9736,17'd28342,17'd18194,17'd16318,17'd9039,17'd8874,17'd15295,17'd10024,17'd10476,17'd16069,17'd12996,17'd12719,17'd12419,17'd12110,17'd11958,17'd19408,17'd24030,17'd25927,17'd26872,17'd26629,17'd27737,17'd24537,17'd23514,17'd23512,17'd24856,17'd28343,17'd28344,17'd28345,17'd27857,17'd28107,17'd22818,17'd16442,17'd15185,17'd16204,17'd16204,17'd12858,17'd12112,17'd16797,17'd11519,17'd19532,17'd16796,17'd9884,17'd17599,17'd26037,17'd10476,17'd11808,17'd11395,17'd16068,17'd11808,17'd11399,17'd12721,17'd21206,17'd10990,17'd11666,17'd13764,17'd11520,17'd10476,17'd12116,17'd22812,17'd9481,17'd8874,17'd15187,17'd12116,17'd11399,17'd23171,17'd28346,17'd25927,17'd28347,17'd28103,17'd28348,17'd27235,17'd28349,17'd28350,17'd28351,17'd28351,17'd28234,17'd26758,17'd16685,17'd16443,17'd11274,17'd11399,17'd11669,17'd28352,17'd24996,17'd11132,17'd17121,17'd21986,17'd11666,17'd16323,17'd13364,17'd11960,17'd12580,17'd12580,17'd12417,17'd12859,17'd12995,17'd12419,17'd15299,17'd13366,17'd11520,17'd10852,17'd10163,17'd9618,17'd24361,17'd28353,17'd24367,17'd8878,17'd9195,17'd8878,17'd26499,17'd28354,17'd28355,17'd28356,17'd28357,17'd28358,17'd28359,17'd28360,17'd28361,17'd28362,17'd28002,17'd28363,17'd27024,17'd24732,17'd28364,17'd24396,17'd24399,17'd25170,17'd25308,17'd25308,17'd24578,17'd25021,17'd26523,17'd25556,17'd25828,17'd25558,17'd25554,17'd25558,17'd26523,17'd26167,17'd25562,17'd24242,17'd23554,17'd23554,17'd24583,17'd25431,17'd28365,17'd25948,17'd27514,17'd26903,17'd25833,17'd28366,17'd25177,17'd28367,17'd24252,17'd28368,17'd25030,17'd28369,17'd26174,17'd27883,17'd24735,17'd25172,17'd25312,17'd26400,17'd26167,17'd26167,17'd25698,17'd25698,17'd25554,17'd26525,17'd25558,17'd26278,17'd26523,17'd25697,17'd28370,17'd28371,17'd28372,17'd28373,17'd28374,17'd28375,17'd28376,17'd28262,17'd28377,17'd27651,17'd27035,17'd28378,17'd28265,17'd26793,17'd28379,17'd26196,17'd28380,17'd28381,17'd28144,17'd28145,17'd28382,17'd28383,17'd28272,17'd28384,17'd27660,17'd28385,17'd25195,17'd25195,17'd28386,17'd28387,17'd28388,17'd28389,17'd26671,17'd25449,17'd24432,17'd28390,17'd28279,17'd23759,17'd28391,17'd28392,17'd28393,17'd28394,17'd28395,17'd18010,17'd17395,17'd28396,17'd18012,17'd28397,17'd19470,17'd28398,17'd28399,17'd28400,17'd28401,17'd28402,17'd28403,17'd28404,17'd28405,17'd28406,17'd28407,17'd28408,17'd28409,17'd28410,17'd28411,17'd28412,17'd28413,17'd28414,17'd28415,17'd22574,17'd28416,17'd22582,17'd24299,17'd24638,17'd24638,17'd21923,17'd25994,17'd21766,17'd11421,17'd28417,17'd7167,17'd6213,17'd8931,17'd5918,17'd6553,17'd8154,17'd10777,17'd11576,17'd10641,17'd27931,17'd27931,17'd27932,17'd28305,17'd28306,17'd11709,17'd11577,17'd10777,17'd10777,17'd9657,17'd28307,17'd28418,17'd4841,17'd5329,17'd5330,17'd5335,17'd5614,17'd26709,17'd9394,17'd11576,17'd12760,17'd12467,17'd14301,17'd14970,17'd17655,17'd15094,17'd15094,17'd15727,17'd28186,17'd13801,17'd16248,17'd14426,17'd15228,17'd28419,17'd23288,17'd28420,17'd12311,17'd16377,17'd16490,17'd28421,17'd24807,17'd23293,17'd28422,17'd28423,17'd28424,17'd28425,17'd28426,17'd28427,17'd933,17'd1240,17'd6868,17'd28428,17'd28315,17'd28429,17'd27581,17'd27095,17'd26967,17'd27320,17'd27319,17'd27319,17'd27319,17'd27319,17'd27320,17'd26968,17'd26968,17'd28316,17'd23817,17'd28192,17'd23480,17'd28317,17'd5638,17'd5638,17'd23133,17'd23133,17'd5638,17'd24325,17'd28430,17'd28431,17'd3229,17'd3716,17'd1954,17'd12638,17'd3728,17'd3730,17'd3236,17'd8642,17'd935,17'd595,17'd1683,17'd15492,17'd17185
},
'{
17'd4428,17'd4892,17'd4892,17'd25384,17'd4245,17'd4733,17'd4733,17'd4733,17'd2934,17'd2593,17'd2935,17'd3101,17'd3252,17'd1831,17'd4247,17'd4247,17'd1416,17'd1416,17'd3905,17'd3905,17'd18,17'd18,17'd1128,17'd20404,17'd653,17'd652,17'd4430,17'd6744,17'd7060,17'd7060,17'd7387,17'd7387,17'd28432,17'd7226,17'd6599,17'd6904,17'd6441,17'd28319,17'd6442,17'd5813,17'd5386,17'd5387,17'd6603,17'd26015,17'd28433,17'd28321,17'd28195,17'd28075,17'd28196,17'd27596,17'd28434,17'd13956,17'd28435,17'd20137,17'd17926,17'd28436,17'd27832,17'd28202,17'd28203,17'd23500,17'd22117,17'd21963,17'd16027,17'd16765,17'd17941,17'd18174,17'd18174,17'd17572,17'd17207,17'd16519,17'd18534,17'd17942,17'd17810,17'd17694,17'd19011,17'd28437,17'd27460,17'd19007,17'd20148,17'd20886,17'd28438,17'd19006,17'd19893,17'd17689,17'd16986,17'd21185,17'd16289,17'd16880,17'd13601,17'd9575,17'd4767,17'd9303,17'd8381,17'd8383,17'd8222,17'd7264,17'd8855,17'd9709,17'd16997,17'd28439,17'd24844,17'd16419,17'd9450,17'd11921,17'd28440,17'd28441,17'd9025,17'd28442,17'd28443,17'd28444,17'd28445,17'd28446,17'd28447,17'd28448,17'd28449,17'd28450,17'd28451,17'd28452,17'd28453,17'd16905,17'd15678,17'd28222,17'd28454,17'd28455,17'd28456,17'd10014,17'd28457,17'd28458,17'd9614,17'd18196,17'd9478,17'd15180,17'd9039,17'd8873,17'd9192,17'd9341,17'd10479,17'd14931,17'd13762,17'd12996,17'd12419,17'd12110,17'd12420,17'd12106,17'd22819,17'd24856,17'd26370,17'd26872,17'd26873,17'd24856,17'd28459,17'd23514,17'd23511,17'd27121,17'd28460,17'd28461,17'd28462,17'd27737,17'd23168,17'd17722,17'd19158,17'd16326,17'd16204,17'd15053,17'd12111,17'd12112,17'd15810,17'd24708,17'd10327,17'd9883,17'd19642,17'd15943,17'd10476,17'd10854,17'd10989,17'd11520,17'd10737,17'd14931,17'd11399,17'd28352,17'd28463,17'd16069,17'd13764,17'd13885,17'd10990,17'd9883,17'd15187,17'd9043,17'd15682,17'd15807,17'd9741,17'd15176,17'd28464,17'd27986,17'd25670,17'd27123,17'd27737,17'd27737,17'd27348,17'd27235,17'd28465,17'd28466,17'd28467,17'd28460,17'd27737,17'd28468,17'd18450,17'd11667,17'd16320,17'd10991,17'd24996,17'd28352,17'd11808,17'd16069,17'd13764,17'd15299,17'd14808,17'd13363,17'd12420,17'd12419,17'd12575,17'd12256,17'd12418,17'd12995,17'd13519,17'd12857,17'd13764,17'd28469,17'd14803,17'd10477,17'd17839,17'd9478,17'd9039,17'd15297,17'd8567,17'd8567,17'd8567,17'd12263,17'd28470,17'd28471,17'd28472,17'd27008,17'd28473,17'd28474,17'd28475,17'd28476,17'd28361,17'd28248,17'd28477,17'd27759,17'd28478,17'd24572,17'd28479,17'd23905,17'd25023,17'd25169,17'd25308,17'd26523,17'd25558,17'd25558,17'd26523,17'd25555,17'd25698,17'd25558,17'd25554,17'd25558,17'd25554,17'd26400,17'd27766,17'd28130,17'd28480,17'd25709,17'd25566,17'd27767,17'd28481,17'd27260,17'd28482,17'd27639,17'd25833,17'd28483,17'd28484,17'd28485,17'd28008,17'd24252,17'd24898,17'd27882,17'd27766,17'd27514,17'd27883,17'd27640,17'd27371,17'd26782,17'd28486,17'd28486,17'd25944,17'd25554,17'd25558,17'd27368,17'd26523,17'd26780,17'd26278,17'd26652,17'd26897,17'd28487,17'd28488,17'd28371,17'd28489,17'd28490,17'd28491,17'd28492,17'd28493,17'd28494,17'd28495,17'd28495,17'd26539,17'd28496,17'd28379,17'd25576,17'd28497,17'd28498,17'd28499,17'd28500,17'd28501,17'd28271,17'd28502,17'd28503,17'd26920,17'd27391,17'd25195,17'd26082,17'd28504,17'd28505,17'd28506,17'd28507,17'd26081,17'd25592,17'd28390,17'd24432,17'd28508,17'd28509,17'd28510,17'd28511,17'd18723,17'd28512,17'd28395,17'd18607,17'd17767,17'd17395,17'd18366,17'd17518,17'd25614,17'd28513,17'd28514,17'd28515,17'd28516,17'd28517,17'd28518,17'd28519,17'd28520,17'd28521,17'd28522,17'd28172,17'd28523,17'd28524,17'd28525,17'd28526,17'd28527,17'd28528,17'd28529,17'd22383,17'd28530,17'd22738,17'd24139,17'd22241,17'd22081,17'd22081,17'd28531,17'd25994,17'd12444,17'd10499,17'd9219,17'd28532,17'd8931,17'd6704,17'd6553,17'd6707,17'd9090,17'd10777,17'd10641,17'd27932,17'd10897,17'd28533,17'd28306,17'd28534,17'd11431,17'd11431,17'd11431,17'd11576,17'd9657,17'd28535,17'd28536,17'd5327,17'd5002,17'd5330,17'd5335,17'd5615,17'd6390,17'd6391,17'd10641,17'd11854,17'd12467,17'd12467,17'd13558,17'd15094,17'd17655,17'd14971,17'd15610,17'd27198,17'd17408,17'd16248,17'd16850,17'd15228,17'd16128,17'd26586,17'd26114,17'd19852,17'd27939,17'd28537,17'd14056,17'd18265,17'd19595,17'd28538,17'd28539,17'd28540,17'd28541,17'd28542,17'd28543,17'd455,17'd2924,17'd2409,17'd28428,17'd28544,17'd27581,17'd28545,17'd28546,17'd27583,17'd27320,17'd27319,17'd27319,17'd27710,17'd27319,17'd27320,17'd26723,17'd26723,17'd27582,17'd28547,17'd28067,17'd23480,17'd28317,17'd28317,17'd28317,17'd28317,17'd5638,17'd26970,17'd27587,17'd28548,17'd15865,17'd3229,17'd3716,17'd2106,17'd3580,17'd3580,17'd3581,17'd10389,17'd23301,17'd21161,17'd804,17'd1683,17'd15492,17'd1543
},
'{
17'd4244,17'd4892,17'd4892,17'd4892,17'd4088,17'd4733,17'd4733,17'd6584,17'd2934,17'd2934,17'd2935,17'd3101,17'd3252,17'd1831,17'd4247,17'd4247,17'd1416,17'd1416,17'd3905,17'd3905,17'd18,17'd18,17'd1128,17'd20404,17'd653,17'd652,17'd6744,17'd6744,17'd7060,17'd7060,17'd7387,17'd7387,17'd7226,17'd7226,17'd6904,17'd6441,17'd28319,17'd28319,17'd6442,17'd5813,17'd5386,17'd27098,17'd5226,17'd12040,17'd4902,17'd5667,17'd3444,17'd27828,17'd28322,17'd28549,17'd28550,17'd28551,17'd28552,17'd19885,17'd18161,17'd28436,17'd28553,17'd28202,17'd27457,17'd22460,17'd21963,17'd16287,17'd16027,17'd20292,17'd18774,17'd17318,17'd17572,17'd17207,17'd17320,17'd16519,17'd18534,17'd17810,17'd17448,17'd18060,17'd27833,17'd19385,17'd25512,17'd19893,17'd18884,17'd20886,17'd28554,17'd19006,17'd19893,17'd27834,17'd21650,17'd16289,17'd16880,17'd13470,17'd12959,17'd8066,17'd5253,17'd9842,17'd8694,17'd28555,17'd8077,17'd8702,17'd16044,17'd16996,17'd17945,17'd28439,17'd24844,17'd16419,17'd9450,17'd28556,17'd28440,17'd28441,17'd27965,17'd28442,17'd28557,17'd9175,17'd28558,17'd28559,17'd28560,17'd28561,17'd28562,17'd28563,17'd28564,17'd28565,17'd10595,17'd25277,17'd21819,17'd28566,17'd28567,17'd10980,17'd10728,17'd9876,17'd28568,17'd9868,17'd28569,17'd9619,17'd15187,17'd15430,17'd9038,17'd8720,17'd16793,17'd10992,17'd12863,17'd14931,17'd11807,17'd13135,17'd12419,17'd12580,17'd16321,17'd12107,17'd24859,17'd27004,17'd26370,17'd26757,17'd28570,17'd24859,17'd23514,17'd24859,17'd26629,17'd28460,17'd28571,17'd28571,17'd27857,17'd24856,17'd19408,17'd18917,17'd19158,17'd19158,17'd18917,17'd13883,17'd11961,17'd11962,17'd11965,17'd10474,17'd10327,17'd11134,17'd17599,17'd11527,17'd11399,17'd25280,17'd11522,17'd11395,17'd10737,17'd10739,17'd14263,17'd13521,17'd12583,17'd17125,17'd23338,17'd15182,17'd11133,17'd9740,17'd21984,17'd17600,17'd10335,17'd9742,17'd11526,17'd17343,17'd27986,17'd24538,17'd25927,17'd27123,17'd27737,17'd27858,17'd27349,17'd28348,17'd28572,17'd28462,17'd28462,17'd28573,17'd28574,17'd28235,17'd13135,17'd10736,17'd10603,17'd10023,17'd27487,17'd10854,17'd11521,17'd13520,17'd18565,17'd28575,17'd14130,17'd12419,17'd12419,17'd12110,17'd12257,17'd12575,17'd12856,17'd12995,17'd12257,17'd13363,17'd13137,17'd24035,17'd15940,17'd28576,17'd28577,17'd28578,17'd9038,17'd8722,17'd28579,17'd28580,17'd28581,17'd28582,17'd28583,17'd28584,17'd26632,17'd28585,17'd28586,17'd28587,17'd28588,17'd28589,17'd28590,17'd28591,17'd28592,17'd28593,17'd25167,17'd24395,17'd23904,17'd24579,17'd24890,17'd24403,17'd26780,17'd26780,17'd25554,17'd25554,17'd26780,17'd25555,17'd25698,17'd25558,17'd26524,17'd26525,17'd25558,17'd25702,17'd28594,17'd25177,17'd28595,17'd28596,17'd28597,17'd28598,17'd28599,17'd28253,17'd26062,17'd28482,17'd27766,17'd28253,17'd28600,17'd27764,17'd28601,17'd24090,17'd24896,17'd25438,17'd28602,17'd27514,17'd27514,17'd27259,17'd27371,17'd26782,17'd28486,17'd28486,17'd25944,17'd25554,17'd25558,17'd27368,17'd26278,17'd26523,17'd26276,17'd26897,17'd26522,17'd28371,17'd28488,17'd28372,17'd28603,17'd28604,17'd28605,17'd28606,17'd27383,17'd26182,17'd28495,17'd28607,17'd26668,17'd28608,17'd28609,17'd25576,17'd28610,17'd28611,17'd28612,17'd28613,17'd28614,17'd26188,17'd28615,17'd25586,17'd28616,17'd28617,17'd27388,17'd28618,17'd28619,17'd28620,17'd28621,17'd28622,17'd28623,17'd25718,17'd28624,17'd28625,17'd26412,17'd28625,17'd22885,17'd28626,17'd28627,17'd28628,17'd27542,17'd16941,17'd17889,17'd17397,17'd28629,17'd28630,17'd25981,17'd19578,17'd28631,17'd28632,17'd28633,17'd22176,17'd28634,17'd28635,17'd28636,17'd28637,17'd28638,17'd28639,17'd28640,17'd28641,17'd28642,17'd28643,17'd28644,17'd28645,17'd20673,17'd28646,17'd22057,17'd28647,17'd22582,17'd24140,17'd22241,17'd22081,17'd28531,17'd25622,17'd28648,17'd20993,17'd28649,17'd7825,17'd6214,17'd7176,17'd9523,17'd6553,17'd9090,17'd10777,17'd27932,17'd27932,17'd28650,17'd28533,17'd28650,17'd28305,17'd11181,17'd11181,17'd11431,17'd11431,17'd27931,17'd26708,17'd4842,17'd5152,17'd5005,17'd5329,17'd5160,17'd5336,17'd5614,17'd6391,17'd10641,17'd14049,17'd12467,17'd12467,17'd13558,17'd14971,17'd17655,17'd14971,17'd15610,17'd12761,17'd14050,17'd16125,17'd16249,17'd15228,17'd14854,17'd17781,17'd20699,17'd19852,17'd12477,17'd19351,17'd14056,17'd18265,17'd19353,17'd28651,17'd28652,17'd28653,17'd26961,17'd28654,17'd28655,17'd28656,17'd1957,17'd5957,17'd28657,17'd28544,17'd27581,17'd28545,17'd28546,17'd27583,17'd27320,17'd27319,17'd27319,17'd27710,17'd27319,17'd27319,17'd26723,17'd26723,17'd27582,17'd28547,17'd28067,17'd23480,17'd28317,17'd28317,17'd28317,17'd5638,17'd5638,17'd28317,17'd24325,17'd28658,17'd28431,17'd3876,17'd2401,17'd2106,17'd3580,17'd3580,17'd3581,17'd3414,17'd23301,17'd2112,17'd1682,17'd180,17'd280,17'd1543
},
'{
17'd3902,17'd3902,17'd3902,17'd4892,17'd4088,17'd3904,17'd4733,17'd4733,17'd6420,17'd4245,17'd3101,17'd3101,17'd3252,17'd1688,17'd4247,17'd4247,17'd1416,17'd1416,17'd1416,17'd17,17'd18,17'd18,17'd3905,17'd3905,17'd653,17'd652,17'd6744,17'd6744,17'd7060,17'd7060,17'd7387,17'd7386,17'd6599,17'd6599,17'd6441,17'd6441,17'd28319,17'd28659,17'd27446,17'd10410,17'd9818,17'd26734,17'd28660,17'd5666,17'd28661,17'd5667,17'd28662,17'd28076,17'd27596,17'd23661,17'd28663,17'd28664,17'd28665,17'd19115,17'd17562,17'd28666,17'd15755,17'd28202,17'd27457,17'd22117,17'd16287,17'd20885,17'd28667,17'd19892,17'd18656,17'd17319,17'd17207,17'd16034,17'd24348,17'd16769,17'd15524,17'd15902,17'd16519,17'd16519,17'd19385,17'd28668,17'd19128,17'd18884,17'd28667,17'd16765,17'd22630,17'd22630,17'd19006,17'd17689,17'd16986,17'd16289,17'd16659,17'd16880,17'd13469,17'd8538,17'd5689,17'd28669,17'd8848,17'd28670,17'd14359,17'd8702,17'd9314,17'd16996,17'd17945,17'd16668,17'd17214,17'd9993,17'd9319,17'd28671,17'd28440,17'd28329,17'd28672,17'd28442,17'd28442,17'd28673,17'd28674,17'd28675,17'd28676,17'd28677,17'd28678,17'd27229,17'd28452,17'd28679,17'd11516,17'd28680,17'd11805,17'd28566,17'd28681,17'd26868,17'd28682,17'd28683,17'd28684,17'd28685,17'd25407,17'd15569,17'd15180,17'd9039,17'd8873,17'd17600,17'd15295,17'd10024,17'd10476,17'd14673,17'd11807,17'd11806,17'd12420,17'd16321,17'd17348,17'd12108,17'd25927,17'd26370,17'd26757,17'd26873,17'd25927,17'd23515,17'd23682,17'd26370,17'd27857,17'd28571,17'd28686,17'd28571,17'd26872,17'd23168,17'd15053,17'd16326,17'd13362,17'd11963,17'd11806,17'd13761,17'd11806,17'd14262,17'd14263,17'd27487,17'd10167,17'd10479,17'd11527,17'd15176,17'd11399,17'd16068,17'd11807,17'd14262,17'd16320,17'd10475,17'd14263,17'd11808,17'd17125,17'd14669,17'd13137,17'd10605,17'd9739,17'd27856,17'd28687,17'd9043,17'd17965,17'd28688,17'd23337,17'd27860,17'd26149,17'd24856,17'd26758,17'd27736,17'd27736,17'd28689,17'd28234,17'd28690,17'd28691,17'd28462,17'd28462,17'd28692,17'd28693,17'd18565,17'd10989,17'd10740,17'd28694,17'd25811,17'd10739,17'd11807,17'd18565,17'd15184,17'd16203,17'd12579,17'd14807,17'd12995,17'd13763,17'd13763,17'd13763,17'd13763,17'd12110,17'd12110,17'd28695,17'd17598,17'd28696,17'd28697,17'd28698,17'd28699,17'd28700,17'd28701,17'd9335,17'd28702,17'd28703,17'd28704,17'd28705,17'd28706,17'd28707,17'd23860,17'd17480,17'd28708,17'd28709,17'd28710,17'd28711,17'd28712,17'd28713,17'd28714,17'd28715,17'd28593,17'd25167,17'd28716,17'd24580,17'd23904,17'd24238,17'd24403,17'd26780,17'd25558,17'd25696,17'd25696,17'd25558,17'd25555,17'd25698,17'd25558,17'd25554,17'd25558,17'd25696,17'd25562,17'd28717,17'd24897,17'd28008,17'd28718,17'd28719,17'd28717,17'd27512,17'd28369,17'd28720,17'd28602,17'd28720,17'd28721,17'd28721,17'd25438,17'd24742,17'd28722,17'd23561,17'd25177,17'd28723,17'd25949,17'd27515,17'd28724,17'd28725,17'd26782,17'd26901,17'd26901,17'd28726,17'd28727,17'd26780,17'd27768,17'd27768,17'd27768,17'd27761,17'd26522,17'd26522,17'd28257,17'd28728,17'd28728,17'd28729,17'd28730,17'd28731,17'd27382,17'd27383,17'd28732,17'd28495,17'd28607,17'd27156,17'd26670,17'd26541,17'd25960,17'd28733,17'd28734,17'd28735,17'd28736,17'd28737,17'd28738,17'd25042,17'd28739,17'd28740,17'd27168,17'd26919,17'd25195,17'd28741,17'd28742,17'd28743,17'd28744,17'd28623,17'd28745,17'd28746,17'd28747,17'd26080,17'd27159,17'd26307,17'd28748,17'd28749,17'd28750,17'd28751,17'd18120,17'd18119,17'd28752,17'd28753,17'd16942,17'd18606,17'd19207,17'd28754,17'd28755,17'd28756,17'd28757,17'd28758,17'd28759,17'd28760,17'd28761,17'd28762,17'd28763,17'd28764,17'd28765,17'd28766,17'd28767,17'd28768,17'd28769,17'd28770,17'd21117,17'd28771,17'd28772,17'd22564,17'd28773,17'd28774,17'd28775,17'd28776,17'd28531,17'd11985,17'd12884,17'd8913,17'd28777,17'd6213,17'd6068,17'd6388,17'd6553,17'd9090,17'd26219,17'd11576,17'd11181,17'd28306,17'd28650,17'd27931,17'd10897,17'd27932,17'd11181,17'd11037,17'd11037,17'd10515,17'd7499,17'd5163,17'd28778,17'd28536,17'd5329,17'd25627,17'd5335,17'd5615,17'd6221,17'd26219,17'd14048,17'd12760,17'd12760,17'd14301,17'd27198,17'd28186,17'd12761,17'd17173,17'd27198,17'd17408,17'd16125,17'd13561,17'd28779,17'd28780,17'd16374,17'd26454,17'd25881,17'd25486,17'd28781,17'd14056,17'd19093,17'd28782,17'd28783,17'd28784,17'd28785,17'd28786,17'd28787,17'd28788,17'd28789,17'd3100,17'd604,17'd15233,17'd28314,17'd26228,17'd27709,17'd28790,17'd28791,17'd27319,17'd27710,17'd28792,17'd28793,17'd27710,17'd27319,17'd26723,17'd26723,17'd27582,17'd28316,17'd28067,17'd23480,17'd28317,17'd28317,17'd28317,17'd5638,17'd5638,17'd28317,17'd24325,17'd2745,17'd3077,17'd3229,17'd1817,17'd2106,17'd3580,17'd3580,17'd3412,17'd3414,17'd23301,17'd26343,17'd1682,17'd15626,17'd770,17'd1116
},
'{
17'd4087,17'd4087,17'd4087,17'd4244,17'd4428,17'd4088,17'd4733,17'd4245,17'd6420,17'd4245,17'd3101,17'd14070,17'd10535,17'd1688,17'd4247,17'd4247,17'd1416,17'd1416,17'd1416,17'd17,17'd3905,17'd3905,17'd3905,17'd3905,17'd653,17'd652,17'd6744,17'd6744,17'd7060,17'd7060,17'd7386,17'd7386,17'd6599,17'd6599,17'd6441,17'd6441,17'd6113,17'd28794,17'd27446,17'd10410,17'd6751,17'd26734,17'd28320,17'd5666,17'd28795,17'd3270,17'd3271,17'd28076,17'd27596,17'd27830,17'd28796,17'd28797,17'd27598,17'd28798,17'd28799,17'd14201,17'd28800,17'd26740,17'd23669,17'd24344,17'd20885,17'd20886,17'd20148,17'd27461,17'd18657,17'd17320,17'd16034,17'd16033,17'd15524,17'd15524,17'd15902,17'd15524,17'd18060,17'd17207,17'd20149,17'd18655,17'd18884,17'd20886,17'd16765,17'd16658,17'd22630,17'd12681,17'd17204,17'd21649,17'd16164,17'd16289,17'd16659,17'd13470,17'd9301,17'd4927,17'd10695,17'd9012,17'd9162,17'd8700,17'd14359,17'd8703,17'd28801,17'd17583,17'd17946,17'd17945,17'd17214,17'd9589,17'd9171,17'd28802,17'd28803,17'd28329,17'd27840,17'd28085,17'd28804,17'd28805,17'd28806,17'd28807,17'd28808,17'd28809,17'd28810,17'd10717,17'd10834,17'd28811,17'd10847,17'd23164,17'd12114,17'd28812,17'd28813,17'd10158,17'd9735,17'd10012,17'd28814,17'd28702,17'd28815,17'd14674,17'd15430,17'd9039,17'd9041,17'd15682,17'd9620,17'd12585,17'd17236,17'd11964,17'd11962,17'd11961,17'd12420,17'd17474,17'd12107,17'd12255,17'd26872,17'd28816,17'd26873,17'd28570,17'd24859,17'd28817,17'd24537,17'd28343,17'd28818,17'd28571,17'd28461,17'd28460,17'd24537,17'd20314,17'd19158,17'd11964,17'd11963,17'd11806,17'd13363,17'd15299,17'd11807,17'd11130,17'd19281,17'd28819,17'd9883,17'd12863,17'd14134,17'd12584,17'd25280,17'd16068,17'd16068,17'd10989,17'd10739,17'd16555,17'd11130,17'd11522,17'd14669,17'd23338,17'd13138,17'd12863,17'd17011,17'd21984,17'd28820,17'd9345,17'd13522,17'd28821,17'd28822,17'd26149,17'd25927,17'd26872,17'd27737,17'd28689,17'd27736,17'd27858,17'd27485,17'd28823,17'd28824,17'd28825,17'd28826,17'd28570,17'd21362,17'd11397,17'd10739,17'd27987,17'd27987,17'd10738,17'd13885,17'd13364,17'd15184,17'd12253,17'd12254,17'd13515,17'd12418,17'd12418,17'd12575,17'd13763,17'd12258,17'd12718,17'd12718,17'd16322,17'd17598,17'd28696,17'd28827,17'd28828,17'd28829,17'd28830,17'd28831,17'd28832,17'd28833,17'd28834,17'd28835,17'd28836,17'd28837,17'd28838,17'd28839,17'd28840,17'd17716,17'd28841,17'd28243,17'd28842,17'd28843,17'd28844,17'd28845,17'd28714,17'd28715,17'd28846,17'd28847,17'd28848,17'd24580,17'd24580,17'd24579,17'd24890,17'd26524,17'd26524,17'd25553,17'd25696,17'd25558,17'd25555,17'd25698,17'd25558,17'd25698,17'd25696,17'd25560,17'd24583,17'd28719,17'd24743,17'd28849,17'd24090,17'd24897,17'd28254,17'd24896,17'd25030,17'd25709,17'd27765,17'd28130,17'd27765,17'd25435,17'd28850,17'd28851,17'd28852,17'd28367,17'd27637,17'd28130,17'd28602,17'd25833,17'd28724,17'd28853,17'd26782,17'd26901,17'd26901,17'd28726,17'd28727,17'd25555,17'd26278,17'd27768,17'd27761,17'd28370,17'd28854,17'd28855,17'd28856,17'd28857,17'd28728,17'd28858,17'd28859,17'd28860,17'd28861,17'd28862,17'd27899,17'd27035,17'd28863,17'd26790,17'd27038,17'd28864,17'd28019,17'd28865,17'd28866,17'd28867,17'd28868,17'd28869,17'd28870,17'd25583,17'd28871,17'd26676,17'd28872,17'd27531,17'd27388,17'd28618,17'd28873,17'd28874,17'd28875,17'd28623,17'd26297,17'd25454,17'd28876,17'd26301,17'd26412,17'd24271,17'd28877,17'd28878,17'd28879,17'd28880,17'd18603,17'd28881,17'd28882,17'd28882,17'd28883,17'd28034,17'd28884,17'd28885,17'd26097,17'd28886,17'd28887,17'd28888,17'd28889,17'd28890,17'd28891,17'd28892,17'd28893,17'd28894,17'd28895,17'd28896,17'd28767,17'd28897,17'd28898,17'd28899,17'd20820,17'd28900,17'd28901,17'd28902,17'd23787,17'd28181,17'd28775,17'd28776,17'd22242,17'd25996,17'd28903,17'd28904,17'd9219,17'd6846,17'd6216,17'd5918,17'd6387,17'd6852,17'd26219,17'd11576,17'd11181,17'd28306,17'd28306,17'd27931,17'd10897,17'd27932,17'd27932,17'd11037,17'd27934,17'd28183,17'd28184,17'd5167,17'd28778,17'd28905,17'd5002,17'd5004,17'd5160,17'd5615,17'd5919,17'd9394,17'd25226,17'd12760,17'd12760,17'd12467,17'd14423,17'd28186,17'd12761,17'd17173,17'd14423,17'd17408,17'd16617,17'd13561,17'd28906,17'd28907,17'd7015,17'd23288,17'd20548,17'd20118,17'd28908,17'd18028,17'd19093,17'd21937,17'd28909,17'd28910,17'd28911,17'd28912,17'd28913,17'd28914,17'd28915,17'd610,17'd411,17'd1383,17'd28916,17'd26228,17'd27580,17'd28790,17'd28917,17'd28791,17'd27710,17'd28792,17'd28793,17'd27710,17'd27319,17'd26723,17'd26723,17'd26722,17'd28316,17'd28192,17'd23480,17'd28317,17'd28317,17'd28317,17'd5638,17'd5638,17'd28317,17'd28430,17'd2564,17'd3079,17'd3876,17'd2401,17'd2106,17'd3580,17'd3580,17'd3237,17'd3414,17'd4421,17'd22100,17'd186,17'd251,17'd433,17'd20001
},
'{
17'd5201,17'd4426,17'd4087,17'd4244,17'd4428,17'd4428,17'd4245,17'd6420,17'd15746,17'd14743,17'd13428,17'd13428,17'd10535,17'd1688,17'd1127,17'd4247,17'd1414,17'd1414,17'd17,17'd17,17'd3905,17'd3905,17'd3905,17'd3905,17'd653,17'd652,17'd6744,17'd6744,17'd6745,17'd6745,17'd7386,17'd7386,17'd6599,17'd6904,17'd6441,17'd6441,17'd28319,17'd28659,17'd27446,17'd10410,17'd6751,17'd6603,17'd12040,17'd3922,17'd28795,17'd28918,17'd28662,17'd28076,17'd28919,17'd28920,17'd28921,17'd28435,17'd20137,17'd19745,17'd18048,17'd28922,17'd28923,17'd28924,17'd23669,17'd24519,17'd28925,17'd19621,17'd19007,17'd19255,17'd17942,17'd15902,17'd16033,17'd16033,17'd15524,17'd15902,17'd16034,17'd15899,17'd16289,17'd19385,17'd28926,17'd17689,17'd20886,17'd20885,17'd14622,17'd15764,17'd13969,17'd16658,17'd19006,17'd17689,17'd16986,17'd16289,17'd16659,17'd16880,17'd9703,17'd5409,17'd10431,17'd8695,17'd8851,17'd16042,17'd12370,17'd11920,17'd18064,17'd28927,17'd17946,17'd16997,17'd9709,17'd9170,17'd28928,17'd28802,17'd28803,17'd28929,17'd27840,17'd28085,17'd28930,17'd28931,17'd28932,17'd28933,17'd28934,17'd28935,17'd28810,17'd28936,17'd28937,17'd10462,17'd28567,17'd28938,17'd11957,17'd28812,17'd28939,17'd28940,17'd9872,17'd9606,17'd28941,17'd28942,17'd24211,17'd24361,17'd9039,17'd9194,17'd9044,17'd9481,17'd17965,17'd15176,17'd16068,17'd13762,17'd11962,17'd12857,17'd12420,17'd17474,17'd23512,17'd24856,17'd26872,17'd28227,17'd26873,17'd24856,17'd26756,17'd25526,17'd28816,17'd28943,17'd28571,17'd28944,17'd28945,17'd26758,17'd16203,17'd18917,17'd11964,17'd11964,17'd11957,17'd12857,17'd13363,17'd13646,17'd11274,17'd27623,17'd10327,17'd21503,17'd11528,17'd11527,17'd11399,17'd25280,17'd14673,17'd14673,17'd11274,17'd10990,17'd16555,17'd10475,17'd10989,17'd13253,17'd15175,17'd15182,17'd11527,17'd12116,17'd9191,17'd28946,17'd9339,17'd18556,17'd13647,17'd28947,17'd28948,17'd24856,17'd26872,17'd27737,17'd27858,17'd27858,17'd27349,17'd28234,17'd28351,17'd28823,17'd28825,17'd28949,17'd28574,17'd28950,17'd18444,17'd14381,17'd27739,17'd27987,17'd10736,17'd19157,17'd11961,17'd12577,17'd12414,17'd13517,17'd14003,17'd14672,17'd13643,17'd13760,17'd13763,17'd13763,17'd12718,17'd23854,17'd21204,17'd18805,17'd17121,17'd28951,17'd28952,17'd28953,17'd28954,17'd28955,17'd28956,17'd28957,17'd28958,17'd28959,17'd28960,17'd28961,17'd28962,17'd28963,17'd23684,17'd28964,17'd28815,17'd28965,17'd28966,17'd28967,17'd28968,17'd28969,17'd28845,17'd28970,17'd28971,17'd28972,17'd25824,17'd28973,17'd28848,17'd24395,17'd24579,17'd23905,17'd26524,17'd26524,17'd25553,17'd25553,17'd26524,17'd26780,17'd25554,17'd26524,17'd25558,17'd25553,17'd26055,17'd23553,17'd28974,17'd28975,17'd28976,17'd23732,17'd24416,17'd24744,17'd24252,17'd24252,17'd24897,17'd25178,17'd28484,17'd28369,17'd25317,17'd27511,17'd28977,17'd28975,17'd23562,17'd24897,17'd28850,17'd28594,17'd26174,17'd28978,17'd28853,17'd28725,17'd26902,17'd26901,17'd28979,17'd28727,17'd28980,17'd27642,17'd26276,17'd27761,17'd28370,17'd28370,17'd28981,17'd28981,17'd28372,17'd28728,17'd28982,17'd28983,17'd28984,17'd28985,17'd27897,17'd26188,17'd28986,17'd28607,17'd28987,17'd27894,17'd28988,17'd28989,17'd28502,17'd28990,17'd28991,17'd28992,17'd28993,17'd24102,17'd25192,17'd25043,17'd26414,17'd28994,17'd27045,17'd28275,17'd28618,17'd28995,17'd28996,17'd28997,17'd28623,17'd25960,17'd25853,17'd27160,17'd26413,17'd26301,17'd24755,17'd22702,17'd28998,17'd28999,17'd29000,17'd17264,17'd20084,17'd20084,17'd29001,17'd19324,17'd27400,17'd29002,17'd18102,17'd23772,17'd29003,17'd29004,17'd29005,17'd29006,17'd29007,17'd29008,17'd29009,17'd29010,17'd29011,17'd29012,17'd29013,17'd29014,17'd29015,17'd29016,17'd29017,17'd29018,17'd29019,17'd29020,17'd29021,17'd23787,17'd28181,17'd28774,17'd28776,17'd22242,17'd24942,17'd12741,17'd29022,17'd9219,17'd6846,17'd24150,17'd26451,17'd6388,17'd6707,17'd9394,17'd10641,17'd11576,17'd27932,17'd27932,17'd27931,17'd10897,17'd27815,17'd10515,17'd28057,17'd27934,17'd28057,17'd10515,17'd5168,17'd28778,17'd29023,17'd29024,17'd25627,17'd5160,17'd5615,17'd5919,17'd9394,17'd25226,17'd11854,17'd11854,17'd11710,17'd12906,17'd12761,17'd16615,17'd13406,17'd16123,17'd17408,17'd16617,17'd29025,17'd29026,17'd29027,17'd29028,17'd23288,17'd25089,17'd29029,17'd29030,17'd16853,17'd19093,17'd21937,17'd29031,17'd29032,17'd29033,17'd29034,17'd29035,17'd1083,17'd29036,17'd403,17'd1111,17'd413,17'd1671,17'd29037,17'd2741,17'd5031,17'd29038,17'd28791,17'd27710,17'd28792,17'd28793,17'd29039,17'd29040,17'd27209,17'd26723,17'd27208,17'd29041,17'd28192,17'd28067,17'd28317,17'd28317,17'd28317,17'd5638,17'd5638,17'd28317,17'd29042,17'd2564,17'd3079,17'd3229,17'd1817,17'd2106,17'd3580,17'd12638,17'd3237,17'd3414,17'd4421,17'd22100,17'd639,17'd770,17'd1116,17'd15742
},
'{
17'd4735,17'd4735,17'd4426,17'd4087,17'd4244,17'd4428,17'd6420,17'd25384,17'd14743,17'd14743,17'd13428,17'd13428,17'd10535,17'd1688,17'd1127,17'd4247,17'd1414,17'd1414,17'd17,17'd17,17'd3905,17'd3905,17'd3905,17'd3905,17'd653,17'd652,17'd6744,17'd6744,17'd6745,17'd6745,17'd7386,17'd7386,17'd6904,17'd6904,17'd6441,17'd6441,17'd28319,17'd6442,17'd5813,17'd5386,17'd5387,17'd6603,17'd12040,17'd3922,17'd29043,17'd3270,17'd3271,17'd28322,17'd27956,17'd13582,17'd29044,17'd26133,17'd29045,17'd17193,17'd29046,17'd28922,17'd26851,17'd29047,17'd23835,17'd29048,17'd19621,17'd19754,17'd21185,17'd17445,17'd16768,17'd16987,17'd16987,17'd16987,17'd15902,17'd15902,17'd16034,17'd15899,17'd17319,17'd29049,17'd19891,17'd17204,17'd12531,17'd20885,17'd14622,17'd29050,17'd13969,17'd12532,17'd17204,17'd21649,17'd16164,17'd16289,17'd16659,17'd13470,17'd7582,17'd6140,17'd9441,17'd8695,17'd8851,17'd16042,17'd12370,17'd10127,17'd18180,17'd28927,17'd17946,17'd18064,17'd9587,17'd9169,17'd28928,17'd28802,17'd29051,17'd28929,17'd29052,17'd29053,17'd29054,17'd29055,17'd29056,17'd29057,17'd29058,17'd29059,17'd28810,17'd29060,17'd29061,17'd29062,17'd11956,17'd12858,17'd13135,17'd16198,17'd10848,17'd9875,17'd9730,17'd9608,17'd29063,17'd29064,17'd16553,17'd9038,17'd9040,17'd9045,17'd17600,17'd9191,17'd11671,17'd14134,17'd16069,17'd11807,17'd12861,17'd12857,17'd11958,17'd14807,17'd24707,17'd26370,17'd26872,17'd26873,17'd28570,17'd23856,17'd26756,17'd29065,17'd28943,17'd29066,17'd29067,17'd28944,17'd27349,17'd23855,17'd18198,17'd16326,17'd11396,17'd11964,17'd12113,17'd12857,17'd11961,17'd11522,17'd11669,17'd26369,17'd17719,17'd9739,17'd29068,17'd10478,17'd11524,17'd11523,17'd11396,17'd11274,17'd10854,17'd10854,17'd29069,17'd10854,17'd11520,17'd13253,17'd16064,17'd10604,17'd11134,17'd9345,17'd16550,17'd17600,17'd9480,17'd19278,17'd13367,17'd29070,17'd24856,17'd28343,17'd28104,17'd27857,17'd27858,17'd29071,17'd28234,17'd28465,17'd28467,17'd28466,17'd28691,17'd28949,17'd24207,17'd16442,17'd24029,17'd29072,17'd10327,17'd10604,17'd13764,17'd11960,17'd12419,17'd12109,17'd12256,17'd12997,17'd14523,17'd14809,17'd15942,17'd14526,17'd12995,17'd13763,17'd12718,17'd12112,17'd16797,17'd16435,17'd29073,17'd29074,17'd29075,17'd29076,17'd29077,17'd29078,17'd29079,17'd29080,17'd29081,17'd29082,17'd29083,17'd29084,17'd29085,17'd29086,17'd29087,17'd29088,17'd29089,17'd29090,17'd29091,17'd29092,17'd29093,17'd29094,17'd29095,17'd29096,17'd29097,17'd28972,17'd26651,17'd29098,17'd28848,17'd24069,17'd24404,17'd23905,17'd25554,17'd25553,17'd26055,17'd25553,17'd26524,17'd26780,17'd25558,17'd26525,17'd26524,17'd25553,17'd26055,17'd24242,17'd28595,17'd23564,17'd23386,17'd29099,17'd24415,17'd24743,17'd23917,17'd28722,17'd29100,17'd24417,17'd29101,17'd28369,17'd25709,17'd25320,17'd25032,17'd24090,17'd29102,17'd28718,17'd29103,17'd27765,17'd25949,17'd28978,17'd27258,17'd26902,17'd26901,17'd28486,17'd28979,17'd28727,17'd28980,17'd27642,17'd26276,17'd27884,17'd28133,17'd28133,17'd29104,17'd29105,17'd29106,17'd28857,17'd29107,17'd29108,17'd29109,17'd29110,17'd29111,17'd24754,17'd28378,17'd29112,17'd26910,17'd29113,17'd27523,17'd26539,17'd27377,17'd29114,17'd29115,17'd29116,17'd29117,17'd29118,17'd29119,17'd25189,17'd26414,17'd27657,17'd25454,17'd29120,17'd27164,17'd27392,17'd29121,17'd29122,17'd28623,17'd29123,17'd27162,17'd29124,17'd29125,17'd29126,17'd29127,17'd29128,17'd22880,17'd29129,17'd29130,17'd29131,17'd29132,17'd29133,17'd29134,17'd17160,17'd28033,17'd29135,17'd20804,17'd29136,17'd29137,17'd29138,17'd29139,17'd29140,17'd29141,17'd29142,17'd29143,17'd29144,17'd29145,17'd29146,17'd29147,17'd29148,17'd29149,17'd29150,17'd29151,17'd29152,17'd20973,17'd29153,17'd29154,17'd22390,17'd29155,17'd24140,17'd29156,17'd28531,17'd25220,17'd29157,17'd10628,17'd8913,17'd7661,17'd6703,17'd5917,17'd26451,17'd6387,17'd9090,17'd10513,17'd10641,17'd27932,17'd27932,17'd10897,17'd10897,17'd27815,17'd10515,17'd28183,17'd28057,17'd29158,17'd10642,17'd29159,17'd4684,17'd29160,17'd4685,17'd25627,17'd5160,17'd5614,17'd5615,17'd9090,17'd12465,17'd11854,17'd11854,17'd29161,17'd12906,17'd12761,17'd16615,17'd13406,17'd12622,17'd17408,17'd15855,17'd13169,17'd29162,17'd29163,17'd7014,17'd29164,17'd25089,17'd29029,17'd25230,17'd16853,17'd18265,17'd21937,17'd29165,17'd29166,17'd29167,17'd29034,17'd29168,17'd1375,17'd21160,17'd403,17'd605,17'd2589,17'd1671,17'd29169,17'd2741,17'd5031,17'd29038,17'd28791,17'd27710,17'd28793,17'd29170,17'd29039,17'd29040,17'd27209,17'd26723,17'd27208,17'd29171,17'd29172,17'd28067,17'd28317,17'd28317,17'd28317,17'd28317,17'd28317,17'd28317,17'd29042,17'd2564,17'd3079,17'd3395,17'd2401,17'd1954,17'd12638,17'd12638,17'd3237,17'd3414,17'd4421,17'd8950,17'd592,17'd1543,17'd20001,17'd29173
},
'{
17'd5197,17'd4734,17'd5646,17'd3902,17'd4892,17'd4428,17'd6420,17'd15876,17'd14743,17'd14743,17'd13428,17'd13428,17'd10535,17'd1688,17'd1127,17'd4247,17'd1414,17'd1415,17'd17,17'd17,17'd3905,17'd3905,17'd3905,17'd3905,17'd653,17'd652,17'd6744,17'd6744,17'd6745,17'd6745,17'd7386,17'd7386,17'd6904,17'd6904,17'd6441,17'd28319,17'd28659,17'd27593,17'd29174,17'd9818,17'd29175,17'd5226,17'd5666,17'd29176,17'd29043,17'd3270,17'd3271,17'd28322,17'd29177,17'd16012,17'd29178,17'd4107,17'd25508,17'd17193,17'd29046,17'd29179,17'd29180,17'd29047,17'd25658,17'd29048,17'd17317,17'd10945,17'd17207,17'd16033,17'd16768,17'd14892,17'd14346,17'd14765,17'd14347,17'd14347,17'd24348,17'd15899,17'd17207,17'd19383,17'd17689,17'd20886,17'd16765,17'd12361,17'd14764,17'd14891,17'd12361,17'd16658,17'd19006,17'd27834,17'd21650,17'd18060,17'd16659,17'd15766,17'd13846,17'd6625,17'd29181,17'd9013,17'd29182,17'd13611,17'd19521,17'd10701,17'd18180,17'd18180,17'd17947,17'd18064,17'd9314,17'd9169,17'd12539,17'd29183,17'd29184,17'd27722,17'd29185,17'd29186,17'd29187,17'd29188,17'd29189,17'd29190,17'd29191,17'd29192,17'd28810,17'd10585,17'd29193,17'd27979,17'd16434,17'd12260,17'd13135,17'd21982,17'd10986,17'd9735,17'd29194,17'd29195,17'd9335,17'd17472,17'd15430,17'd8873,17'd9348,17'd8881,17'd16910,17'd9344,17'd19642,17'd11524,17'd13000,17'd11963,17'd12999,17'd12113,17'd11958,17'd12579,17'd25927,17'd26370,17'd27737,17'd27858,17'd24856,17'd23682,17'd29196,17'd29197,17'd29066,17'd28686,17'd29198,17'd28945,17'd27486,17'd15570,17'd17843,17'd12262,17'd11395,17'd11666,17'd18077,17'd15809,17'd11962,17'd11275,17'd19281,17'd16796,17'd9618,17'd27482,17'd29199,17'd10477,17'd14810,17'd11396,17'd11396,17'd11808,17'd11399,17'd11669,17'd11669,17'd14673,17'd13253,17'd17598,17'd11519,17'd10740,17'd10742,17'd9043,17'd16066,17'd10336,17'd15566,17'd12584,17'd28822,17'd29200,17'd26872,17'd28229,17'd28348,17'd28348,17'd28234,17'd27485,17'd28351,17'd28823,17'd29201,17'd29201,17'd28825,17'd18083,17'd18197,17'd29202,17'd29203,17'd27739,17'd10991,17'd15805,17'd13883,17'd12253,17'd12997,17'd12575,17'd13512,17'd29204,17'd29205,17'd29206,17'd29207,17'd29208,17'd13518,17'd13136,17'd12113,17'd12114,17'd15186,17'd18915,17'd29209,17'd29210,17'd29211,17'd29212,17'd29213,17'd29214,17'd29215,17'd29216,17'd29217,17'd29218,17'd29219,17'd29220,17'd29221,17'd29222,17'd29223,17'd29224,17'd29225,17'd29226,17'd29227,17'd29228,17'd29229,17'd29230,17'd29231,17'd29232,17'd29233,17'd29234,17'd29235,17'd29236,17'd29237,17'd29238,17'd29239,17'd24238,17'd25554,17'd25696,17'd25560,17'd26055,17'd25553,17'd25554,17'd25698,17'd25558,17'd25554,17'd26167,17'd25702,17'd25316,17'd29240,17'd23384,17'd23923,17'd23736,17'd23732,17'd23917,17'd29241,17'd29242,17'd23565,17'd28852,17'd27637,17'd28369,17'd25438,17'd28254,17'd25032,17'd24742,17'd29243,17'd29100,17'd29244,17'd28369,17'd28602,17'd28724,17'd27258,17'd28853,17'd27027,17'd28486,17'd28727,17'd29245,17'd29246,17'd27642,17'd27761,17'd27884,17'd28133,17'd28256,17'd28257,17'd29247,17'd29248,17'd29249,17'd29107,17'd29250,17'd29251,17'd29252,17'd24102,17'd27033,17'd27036,17'd29253,17'd28017,17'd26790,17'd27156,17'd26668,17'd29254,17'd29255,17'd29256,17'd25319,17'd29257,17'd29258,17'd29259,17'd27528,17'd24909,17'd27899,17'd26086,17'd25845,17'd25195,17'd27392,17'd29260,17'd29261,17'd28623,17'd27167,17'd28389,17'd29262,17'd26676,17'd26189,17'd29263,17'd29264,17'd23059,17'd29265,17'd29266,17'd29267,17'd27791,17'd29268,17'd29269,17'd29270,17'd29271,17'd29272,17'd29273,17'd24932,17'd29274,17'd29275,17'd29276,17'd29277,17'd29278,17'd29279,17'd29280,17'd29281,17'd29282,17'd29283,17'd29284,17'd29285,17'd29286,17'd29287,17'd29288,17'd29289,17'd29290,17'd21124,17'd22226,17'd29291,17'd22409,17'd22410,17'd23968,17'd28531,17'd25482,17'd11830,17'd10359,17'd29292,17'd7328,17'd7328,17'd24150,17'd5917,17'd5918,17'd7999,17'd9090,17'd10777,17'd27932,17'd27932,17'd27932,17'd10897,17'd27815,17'd10515,17'd28183,17'd28183,17'd29158,17'd28057,17'd29293,17'd27697,17'd29294,17'd29295,17'd5004,17'd5160,17'd5614,17'd5615,17'd6220,17'd29296,17'd11854,17'd14049,17'd11577,17'd13046,17'd16615,17'd16615,17'd13406,17'd29297,17'd29298,17'd16617,17'd12165,17'd29299,17'd29300,17'd7014,17'd29164,17'd22091,17'd29029,17'd19853,17'd29301,17'd15100,17'd18506,17'd29302,17'd29303,17'd29304,17'd29305,17'd26593,17'd25893,17'd18632,17'd404,17'd644,17'd193,17'd776,17'd29169,17'd2741,17'd5360,17'd3224,17'd27319,17'd27710,17'd28793,17'd29170,17'd29039,17'd29040,17'd27209,17'd26723,17'd27208,17'd29171,17'd29172,17'd28067,17'd23989,17'd23989,17'd28317,17'd28317,17'd23306,17'd23989,17'd29042,17'd2564,17'd3079,17'd3080,17'd1817,17'd1954,17'd12638,17'd3235,17'd3237,17'd3414,17'd4421,17'd22100,17'd1683,17'd589,17'd281,17'd16746
},
'{
17'd5374,17'd6263,17'd4734,17'd4426,17'd4892,17'd6420,17'd6420,17'd6420,17'd4245,17'd14743,17'd13428,17'd13428,17'd1831,17'd1689,17'd1127,17'd4247,17'd1414,17'd1415,17'd17,17'd17,17'd3905,17'd3905,17'd3905,17'd3905,17'd653,17'd652,17'd6744,17'd6744,17'd6745,17'd6745,17'd7386,17'd7386,17'd6904,17'd6904,17'd6441,17'd28319,17'd28659,17'd27446,17'd10410,17'd5387,17'd5388,17'd5665,17'd5666,17'd3921,17'd29043,17'd3270,17'd29306,17'd2798,17'd29307,17'd29308,17'd29309,17'd4107,17'd25508,17'd18161,17'd18526,17'd29310,17'd29180,17'd28203,17'd25511,17'd28925,17'd19754,17'd17318,17'd16034,17'd16411,17'd14346,17'd14893,17'd14346,17'd16032,17'd14347,17'd14347,17'd24348,17'd17319,17'd29049,17'd19891,17'd17317,17'd20424,17'd12361,17'd12361,17'd14621,17'd15764,17'd12361,17'd12532,17'd17317,17'd21649,17'd16164,17'd16659,17'd16659,17'd13469,17'd6143,17'd7249,17'd9578,17'd9443,17'd9014,17'd13611,17'd10818,17'd10701,17'd17947,17'd18180,17'd18180,17'd18064,17'd9314,17'd9169,17'd14490,17'd28802,17'd28440,17'd27722,17'd29311,17'd29312,17'd29313,17'd29314,17'd29315,17'd29316,17'd29317,17'd29318,17'd29319,17'd29320,17'd29321,17'd11956,17'd12114,17'd12996,17'd13135,17'd16435,17'd29322,17'd29323,17'd29324,17'd29325,17'd9039,17'd17472,17'd17123,17'd16067,17'd8723,17'd8881,17'd19033,17'd9479,17'd26037,17'd13138,17'd11666,17'd11962,17'd12861,17'd12113,17'd12106,17'd12254,17'd27123,17'd26370,17'd27858,17'd26873,17'd24859,17'd29326,17'd29327,17'd29328,17'd29329,17'd29067,17'd29330,17'd28572,17'd12255,17'd17967,17'd17604,17'd12262,17'd11667,17'd18679,17'd12258,17'd12112,17'd11395,17'd11669,17'd10167,17'd10169,17'd14928,17'd25676,17'd17720,17'd10604,17'd16068,17'd11397,17'd11274,17'd11274,17'd11399,17'd28352,17'd11275,17'd11520,17'd13885,17'd29331,17'd29332,17'd17839,17'd9743,17'd29333,17'd29334,17'd10334,17'd29335,17'd28464,17'd28948,17'd26872,17'd28228,17'd28818,17'd28460,17'd29336,17'd28350,17'd28351,17'd28823,17'd29337,17'd29337,17'd28691,17'd28570,17'd21363,17'd18444,17'd29203,17'd29338,17'd10475,17'd15432,17'd13253,17'd16203,17'd18564,17'd13884,17'd12997,17'd13760,17'd14521,17'd29339,17'd29340,17'd29340,17'd29340,17'd13881,17'd12259,17'd18447,17'd29341,17'd29342,17'd29343,17'd29344,17'd29076,17'd29345,17'd29346,17'd29347,17'd29348,17'd29349,17'd29350,17'd29351,17'd29352,17'd29353,17'd29354,17'd29355,17'd29356,17'd29357,17'd29358,17'd29359,17'd29360,17'd29361,17'd29362,17'd29363,17'd29364,17'd29365,17'd29366,17'd29367,17'd29368,17'd29369,17'd29370,17'd29371,17'd29372,17'd29373,17'd24404,17'd26055,17'd26055,17'd25560,17'd25560,17'd26167,17'd25944,17'd26394,17'd25698,17'd25554,17'd26279,17'd25703,17'd25176,17'd28367,17'd28976,17'd29374,17'd23387,17'd23918,17'd29375,17'd29241,17'd23386,17'd29376,17'd29377,17'd28718,17'd29244,17'd27511,17'd28596,17'd25032,17'd28851,17'd29378,17'd28722,17'd25179,17'd28369,17'd26064,17'd28724,17'd27258,17'd26902,17'd26901,17'd28486,17'd28727,17'd29245,17'd29379,17'd27642,17'd27761,17'd27884,17'd28133,17'd28371,17'd28371,17'd29380,17'd28857,17'd29249,17'd29381,17'd29382,17'd29383,17'd29384,17'd24263,17'd29385,17'd27036,17'd29112,17'd27035,17'd27379,17'd27034,17'd27652,17'd26296,17'd29252,17'd26403,17'd29386,17'd29387,17'd29388,17'd29389,17'd25191,17'd29390,17'd27899,17'd27043,17'd25731,17'd27163,17'd29391,17'd29392,17'd29393,17'd29394,17'd27167,17'd29395,17'd27386,17'd29396,17'd26302,17'd29397,17'd29398,17'd29399,17'd22030,17'd29400,17'd29401,17'd29267,17'd29402,17'd29403,17'd29404,17'd18234,17'd26091,17'd29405,17'd29406,17'd23959,17'd29407,17'd29408,17'd29409,17'd29410,17'd29411,17'd29412,17'd29413,17'd29414,17'd29415,17'd29416,17'd29417,17'd29418,17'd29149,17'd29419,17'd29420,17'd29421,17'd29422,17'd29423,17'd29424,17'd23617,17'd22583,17'd29425,17'd28531,17'd25482,17'd29426,17'd29427,17'd29292,17'd7660,17'd7166,17'd24150,17'd5917,17'd5918,17'd9523,17'd8154,17'd10513,17'd10897,17'd27932,17'd27932,17'd10897,17'd27815,17'd27815,17'd27933,17'd28183,17'd29158,17'd27934,17'd29428,17'd29429,17'd29430,17'd29431,17'd5005,17'd25627,17'd5336,17'd5919,17'd6220,17'd10514,17'd14049,17'd14049,17'd11854,17'd13046,17'd16615,17'd16615,17'd13406,17'd12622,17'd17408,17'd15855,17'd29432,17'd29299,17'd29026,17'd7502,17'd29433,17'd8158,17'd19852,17'd29434,17'd29435,17'd15100,17'd21937,17'd29436,17'd22951,17'd29437,17'd29438,17'd29439,17'd26008,17'd1236,17'd1960,17'd970,17'd11445,17'd29440,17'd1950,17'd29037,17'd2741,17'd29038,17'd28792,17'd27822,17'd28793,17'd29170,17'd29441,17'd29040,17'd27209,17'd26723,17'd27208,17'd29171,17'd29172,17'd28067,17'd23989,17'd23989,17'd23989,17'd28317,17'd23306,17'd5363,17'd2910,17'd2564,17'd3079,17'd3395,17'd2401,17'd1954,17'd12638,17'd3235,17'd3412,17'd3414,17'd4421,17'd8950,17'd592,17'd589,17'd281,17'd29442
},
'{
17'd7046,17'd6262,17'd5053,17'd10533,17'd4428,17'd6420,17'd25384,17'd27951,17'd3427,17'd2934,17'd2935,17'd2422,17'd1831,17'd4247,17'd4247,17'd4247,17'd1416,17'd17,17'd17,17'd17,17'd17,17'd17,17'd17,17'd17,17'd653,17'd652,17'd6744,17'd6744,17'd7225,17'd7225,17'd7386,17'd7386,17'd6904,17'd6904,17'd29443,17'd29444,17'd28659,17'd27446,17'd5523,17'd27098,17'd29445,17'd29446,17'd29447,17'd28661,17'd29448,17'd29449,17'd3111,17'd29450,17'd16012,17'd29451,17'd29452,17'd29453,17'd29045,17'd18285,17'd24187,17'd27455,17'd29454,17'd24011,17'd24684,17'd29455,17'd27834,17'd17207,17'd16169,17'd16411,17'd16987,17'd16768,17'd14346,17'd14768,17'd24192,17'd15902,17'd18060,17'd17207,17'd19620,17'd19382,17'd20424,17'd12362,17'd12362,17'd14622,17'd14622,17'd14622,17'd12815,17'd12532,17'd17941,17'd21649,17'd16164,17'd16880,17'd15766,17'd9300,17'd6769,17'd10117,17'd9579,17'd9581,17'd14109,17'd9165,17'd9312,17'd9708,17'd17947,17'd17947,17'd29456,17'd28801,17'd7428,17'd29457,17'd11240,17'd29458,17'd29459,17'd29460,17'd29461,17'd29462,17'd29463,17'd29464,17'd29465,17'd29466,17'd29467,17'd10834,17'd29468,17'd29469,17'd10729,17'd28938,17'd19157,17'd11520,17'd11520,17'd24860,17'd29470,17'd9870,17'd29471,17'd29472,17'd25531,17'd28353,17'd29473,17'd9046,17'd8727,17'd29474,17'd26626,17'd9739,17'd10739,17'd11666,17'd11807,17'd12861,17'd13135,17'd18197,17'd23168,17'd24856,17'd26872,17'd28227,17'd29475,17'd27347,17'd23856,17'd28105,17'd29476,17'd29328,17'd28944,17'd29198,17'd28466,17'd27121,17'd20314,17'd18681,17'd18444,17'd11963,17'd12111,17'd15809,17'd18077,17'd15186,17'd11132,17'd10024,17'd9742,17'd15566,17'd19642,17'd19532,17'd10990,17'd11965,17'd16068,17'd16068,17'd11399,17'd11399,17'd11399,17'd14263,17'd13362,17'd12861,17'd29477,17'd28697,17'd11277,17'd10173,17'd17607,17'd16202,17'd29478,17'd29479,17'd23513,17'd23855,17'd27348,17'd28945,17'd28691,17'd28345,17'd29480,17'd29481,17'd29482,17'd29483,17'd29484,17'd29485,17'd29486,17'd29487,17'd29488,17'd23337,17'd28352,17'd19281,17'd11131,17'd11520,17'd21204,17'd12577,17'd15434,17'd16685,17'd12997,17'd12575,17'd13881,17'd13881,17'd29489,17'd29490,17'd29489,17'd29490,17'd29491,17'd29492,17'd29493,17'd24360,17'd29494,17'd29495,17'd29496,17'd29497,17'd29498,17'd29499,17'd29347,17'd29500,17'd29501,17'd29216,17'd28959,17'd29502,17'd29503,17'd29504,17'd29505,17'd29506,17'd29507,17'd29508,17'd10323,17'd29509,17'd29510,17'd29511,17'd29512,17'd29513,17'd29514,17'd29515,17'd29516,17'd29517,17'd29369,17'd29518,17'd29519,17'd29520,17'd29521,17'd29522,17'd29523,17'd29524,17'd29525,17'd26055,17'd26055,17'd26167,17'd25429,17'd26279,17'd25554,17'd25311,17'd28252,17'd25317,17'd24743,17'd29526,17'd23923,17'd29374,17'd23565,17'd29527,17'd29528,17'd29529,17'd29530,17'd29531,17'd29532,17'd29533,17'd25568,17'd27512,17'd24744,17'd29534,17'd29528,17'd29378,17'd24898,17'd27765,17'd27513,17'd26174,17'd29535,17'd27258,17'd27027,17'd28486,17'd28727,17'd28980,17'd29246,17'd29379,17'd27884,17'd28256,17'd28257,17'd28728,17'd29536,17'd29106,17'd28372,17'd29537,17'd29538,17'd29539,17'd29540,17'd29541,17'd28731,17'd29542,17'd29543,17'd29544,17'd27266,17'd29545,17'd26910,17'd27265,17'd27265,17'd29546,17'd29547,17'd29548,17'd29549,17'd29550,17'd29551,17'd29552,17'd27528,17'd26797,17'd26086,17'd26084,17'd27900,17'd27163,17'd29553,17'd29554,17'd29555,17'd29556,17'd29557,17'd29558,17'd29559,17'd29560,17'd29561,17'd29562,17'd27888,17'd29563,17'd29564,17'd29400,17'd29565,17'd26804,17'd29566,17'd26310,17'd28750,17'd29567,17'd29568,17'd29569,17'd29570,17'd29571,17'd29572,17'd29573,17'd29574,17'd29575,17'd29279,17'd29576,17'd29577,17'd29578,17'd29579,17'd29580,17'd29581,17'd29582,17'd29583,17'd29584,17'd29585,17'd29586,17'd21584,17'd29587,17'd29588,17'd22753,17'd23788,17'd29589,17'd22412,17'd25996,17'd29590,17'd10627,17'd7327,17'd7166,17'd5916,17'd5918,17'd9523,17'd7999,17'd29591,17'd9931,17'd10513,17'd10777,17'd27932,17'd27932,17'd29592,17'd29593,17'd29592,17'd27933,17'd28183,17'd11037,17'd11316,17'd6392,17'd29594,17'd29595,17'd4841,17'd5329,17'd5334,17'd5762,17'd7499,17'd29592,17'd11037,17'd13678,17'd11854,17'd12467,17'd12622,17'd27198,17'd12467,17'd14301,17'd12161,17'd29596,17'd29597,17'd29025,17'd28906,17'd29598,17'd10898,17'd29599,17'd12474,17'd29600,17'd20854,17'd29601,17'd21937,17'd29602,17'd29603,17'd29604,17'd29605,17'd29606,17'd29607,17'd29608,17'd933,17'd259,17'd11445,17'd29440,17'd29609,17'd26966,17'd29610,17'd29611,17'd29612,17'd2743,17'd28793,17'd29170,17'd29039,17'd29039,17'd27710,17'd27319,17'd27320,17'd27320,17'd29613,17'd28067,17'd28192,17'd23480,17'd23479,17'd23306,17'd23479,17'd29614,17'd28658,17'd14737,17'd3079,17'd3080,17'd1816,17'd19495,17'd12916,17'd28318,17'd3581,17'd3414,17'd4421,17'd2112,17'd1683,17'd17423,17'd16746,17'd16263
},
'{
17'd7883,17'd7369,17'd10532,17'd10533,17'd4892,17'd25384,17'd4243,17'd4243,17'd3901,17'd2934,17'd2935,17'd2422,17'd1831,17'd4247,17'd4247,17'd4247,17'd1416,17'd17,17'd17,17'd17,17'd17,17'd17,17'd17,17'd17,17'd653,17'd652,17'd6744,17'd6744,17'd7225,17'd7225,17'd7386,17'd7388,17'd6904,17'd6904,17'd29443,17'd29444,17'd28659,17'd27446,17'd5524,17'd5062,17'd5665,17'd5666,17'd4902,17'd28795,17'd29448,17'd29449,17'd29615,17'd29616,17'd29308,17'd29617,17'd29618,17'd29453,17'd20017,17'd18285,17'd29619,17'd26851,17'd29620,17'd24343,17'd29621,17'd29622,17'd19259,17'd17445,17'd16411,17'd16411,17'd16987,17'd16768,17'd14346,17'd14346,17'd16411,17'd24348,17'd16289,17'd19383,17'd19511,17'd19006,17'd20885,17'd12815,17'd14470,17'd14622,17'd14622,17'd12361,17'd20424,17'd17317,17'd16766,17'd10945,17'd29623,17'd16880,17'd9703,17'd8537,17'd6770,17'd10432,17'd9579,17'd9581,17'd14109,17'd9165,17'd9312,17'd9708,17'd18787,17'd17947,17'd29456,17'd28801,17'd7428,17'd29457,17'd11767,17'd29624,17'd29625,17'd29460,17'd28211,17'd29626,17'd29627,17'd29628,17'd29190,17'd29629,17'd29630,17'd29631,17'd29632,17'd29633,17'd29634,17'd11963,17'd11395,17'd11395,17'd12720,17'd29332,17'd24028,17'd9608,17'd29635,17'd29636,17'd29637,17'd29638,17'd29639,17'd24368,17'd12723,17'd8405,17'd23165,17'd10022,17'd14931,17'd11667,17'd11962,17'd13135,17'd15053,17'd20314,17'd24859,17'd26370,17'd28343,17'd27984,17'd26873,17'd25527,17'd29640,17'd29641,17'd27984,17'd28462,17'd29642,17'd29201,17'd27857,17'd24859,17'd22472,17'd18327,17'd11964,17'd11806,17'd13763,17'd13763,17'd12999,17'd10737,17'd10479,17'd18556,17'd17232,17'd29643,17'd19155,17'd21206,17'd13516,17'd11964,17'd14673,17'd14673,17'd11524,17'd21206,17'd21206,17'd11808,17'd11962,17'd12112,17'd29331,17'd10606,17'd16065,17'd24212,17'd8411,17'd10337,17'd27744,17'd23166,17'd22819,17'd27234,17'd29644,17'd28572,17'd28229,17'd28943,17'd29645,17'd29646,17'd29647,17'd29648,17'd29484,17'd29649,17'd29650,17'd15184,17'd12583,17'd12423,17'd19280,17'd15176,17'd14673,17'd20313,17'd13763,17'd18684,17'd12859,17'd12997,17'd16799,17'd18684,17'd13760,17'd29489,17'd29651,17'd29652,17'd29653,17'd29654,17'd29492,17'd29655,17'd10987,17'd29656,17'd29657,17'd29658,17'd29659,17'd29660,17'd27480,17'd29497,17'd29661,17'd29501,17'd29662,17'd29663,17'd29664,17'd29664,17'd29664,17'd29665,17'd29666,17'd29667,17'd29668,17'd29669,17'd29670,17'd10850,17'd29671,17'd29672,17'd29673,17'd29513,17'd29674,17'd29675,17'd29676,17'd29677,17'd29678,17'd29519,17'd29679,17'd29680,17'd29681,17'd29682,17'd29683,17'd29684,17'd28365,17'd25560,17'd25559,17'd26055,17'd26167,17'd26167,17'd25698,17'd25312,17'd25707,17'd28484,17'd24252,17'd29685,17'd29686,17'd29374,17'd29242,17'd29241,17'd24087,17'd29687,17'd23923,17'd29374,17'd23385,17'd29688,17'd25177,17'd25568,17'd24745,17'd29534,17'd29528,17'd29689,17'd24897,17'd25567,17'd27513,17'd27514,17'd27258,17'd27027,17'd26901,17'd28727,17'd29246,17'd29246,17'd29246,17'd29379,17'd27884,17'd28256,17'd28257,17'd28857,17'd29690,17'd29691,17'd29692,17'd29536,17'd29538,17'd29693,17'd29694,17'd29695,17'd29696,17'd29697,17'd29698,17'd29699,17'd29700,17'd29700,17'd26910,17'd27265,17'd27037,17'd27653,17'd29701,17'd29702,17'd29703,17'd29704,17'd27890,17'd29705,17'd25191,17'd27042,17'd25337,17'd26084,17'd27387,17'd27273,17'd29706,17'd26548,17'd29707,17'd28506,17'd29708,17'd29558,17'd29709,17'd26414,17'd29384,17'd29710,17'd29711,17'd29712,17'd23058,17'd29713,17'd29714,17'd29715,17'd29716,17'd29717,17'd26686,17'd20957,17'd29718,17'd29719,17'd29720,17'd29721,17'd29722,17'd29723,17'd29724,17'd29725,17'd29726,17'd29727,17'd29728,17'd29729,17'd29730,17'd29731,17'd29581,17'd29732,17'd29733,17'd29734,17'd28898,17'd29735,17'd21430,17'd29736,17'd22396,17'd22565,17'd22583,17'd29737,17'd24303,17'd24942,17'd11830,17'd10882,17'd29022,17'd7166,17'd5916,17'd6552,17'd9523,17'd7999,17'd29591,17'd9931,17'd10513,17'd10777,17'd11181,17'd27932,17'd29592,17'd29592,17'd29592,17'd27933,17'd10642,17'd10642,17'd28057,17'd10514,17'd5328,17'd29738,17'd4841,17'd5002,17'd29739,17'd5762,17'd29740,17'd29593,17'd10642,17'd13678,17'd25085,17'd24653,17'd12622,17'd14423,17'd12467,17'd14301,17'd12161,17'd29596,17'd29597,17'd29025,17'd16850,17'd14303,17'd29741,17'd7182,17'd12474,17'd26115,17'd20854,17'd29601,17'd21937,17'd29742,17'd29743,17'd29744,17'd29745,17'd29746,17'd29747,17'd29748,17'd29749,17'd954,17'd11600,17'd29750,17'd29609,17'd29751,17'd29170,17'd29611,17'd29611,17'd29752,17'd29170,17'd29170,17'd29039,17'd29039,17'd27710,17'd27319,17'd27320,17'd27320,17'd29613,17'd28192,17'd28192,17'd23480,17'd23479,17'd23306,17'd23479,17'd23479,17'd29613,17'd14737,17'd3079,17'd3080,17'd1816,17'd19495,17'd12916,17'd28318,17'd3581,17'd3414,17'd4421,17'd1239,17'd592,17'd214,17'd29753,17'd16263
},
'{
17'd7882,17'd29754,17'd29755,17'd29756,17'd4892,17'd27951,17'd27713,17'd4892,17'd3901,17'd2934,17'd2935,17'd1831,17'd4247,17'd4247,17'd4247,17'd4247,17'd1416,17'd17,17'd17,17'd17,17'd17,17'd17,17'd17,17'd17,17'd653,17'd652,17'd7060,17'd7061,17'd7225,17'd7225,17'd7386,17'd7388,17'd6904,17'd6904,17'd29443,17'd29444,17'd28659,17'd10410,17'd5387,17'd6603,17'd12040,17'd5666,17'd29176,17'd29757,17'd29758,17'd3111,17'd2954,17'd29759,17'd29760,17'd29761,17'd26982,17'd29762,17'd25508,17'd17087,17'd18049,17'd24189,17'd29047,17'd24518,17'd29763,17'd29764,17'd21185,17'd17690,17'd24192,17'd14767,17'd16987,17'd16768,17'd16768,17'd16987,17'd16033,17'd24348,17'd17319,17'd20149,17'd18774,17'd12532,17'd12815,17'd17940,17'd14621,17'd14621,17'd14470,17'd14622,17'd16658,17'd19006,17'd17689,17'd17205,17'd17318,17'd29623,17'd9159,17'd6143,17'd7249,17'd10118,17'd9580,17'd9582,17'd9309,17'd9311,17'd9446,17'd9708,17'd18787,17'd18787,17'd18420,17'd28801,17'd16294,17'd7764,17'd11767,17'd29624,17'd29765,17'd29766,17'd29767,17'd29768,17'd29769,17'd29770,17'd29771,17'd29772,17'd29773,17'd27340,17'd29774,17'd28339,17'd29775,17'd11962,17'd11395,17'd14262,17'd11274,17'd10739,17'd23852,17'd29776,17'd29777,17'd29636,17'd29637,17'd16317,17'd8570,17'd8412,17'd8409,17'd8722,17'd16554,17'd10606,17'd12720,17'd11807,17'd11806,17'd16204,17'd17722,17'd23168,17'd24856,17'd29778,17'd28227,17'd28106,17'd26872,17'd29326,17'd29778,17'd29328,17'd28571,17'd29779,17'd29780,17'd28572,17'd28107,17'd29781,17'd20609,17'd16326,17'd11963,17'd11961,17'd13763,17'd13365,17'd11963,17'd16555,17'd16796,17'd9885,17'd15566,17'd17469,17'd14134,17'd11399,17'd13516,17'd13762,17'd11274,17'd11808,17'd11524,17'd21206,17'd11131,17'd11520,17'd12861,17'd20313,17'd16320,17'd9739,17'd15944,17'd8882,17'd10338,17'd26153,17'd29782,17'd29783,17'd25925,17'd28234,17'd29784,17'd28465,17'd28229,17'd28345,17'd29482,17'd29785,17'd29786,17'd29484,17'd29787,17'd29788,17'd18564,17'd18681,17'd29789,17'd29790,17'd11669,17'd17236,17'd13253,17'd12718,17'd12257,17'd13512,17'd29205,17'd29791,17'd29205,17'd29340,17'd29792,17'd29651,17'd29651,17'd29653,17'd29793,17'd21819,17'd29794,17'd29795,17'd10986,17'd26147,17'd29796,17'd29797,17'd10461,17'd10016,17'd27232,17'd29798,17'd29799,17'd29800,17'd29801,17'd29802,17'd29803,17'd29803,17'd29804,17'd29805,17'd29806,17'd29807,17'd29808,17'd29809,17'd29810,17'd29811,17'd28699,17'd29812,17'd29813,17'd29814,17'd29815,17'd29816,17'd29817,17'd29818,17'd29819,17'd29820,17'd29821,17'd29680,17'd29822,17'd29823,17'd29824,17'd29683,17'd25830,17'd25702,17'd26055,17'd25559,17'd26055,17'd25696,17'd25698,17'd25313,17'd25707,17'd29825,17'd23916,17'd29685,17'd29826,17'd23923,17'd23385,17'd24086,17'd29241,17'd29827,17'd29828,17'd29829,17'd29830,17'd23731,17'd25320,17'd25177,17'd24895,17'd23916,17'd29527,17'd29689,17'd24896,17'd28369,17'd27513,17'd26174,17'd28978,17'd27027,17'd26901,17'd28727,17'd29246,17'd29246,17'd29379,17'd27642,17'd27884,17'd28256,17'd28257,17'd29537,17'd29831,17'd29690,17'd29832,17'd29831,17'd29833,17'd29693,17'd29834,17'd29835,17'd28860,17'd29836,17'd29837,17'd29838,17'd29700,17'd29700,17'd29839,17'd26909,17'd27034,17'd29840,17'd29841,17'd29842,17'd29843,17'd29844,17'd29712,17'd29845,17'd25965,17'd25336,17'd25337,17'd29846,17'd29847,17'd26919,17'd28873,17'd29554,17'd28505,17'd29848,17'd29849,17'd26791,17'd26410,17'd28140,17'd29850,17'd29851,17'd29852,17'd27772,17'd29853,17'd29854,17'd29855,17'd29856,17'd29857,17'd29858,17'd22198,17'd29859,17'd29860,17'd29861,17'd29862,17'd29863,17'd29864,17'd29865,17'd29866,17'd29867,17'd29868,17'd29869,17'd29870,17'd29871,17'd29872,17'd29873,17'd29874,17'd29875,17'd29876,17'd29877,17'd29878,17'd29879,17'd29880,17'd29881,17'd29882,17'd22568,17'd23618,17'd29883,17'd23969,17'd22412,17'd22413,17'd26826,17'd7824,17'd7166,17'd6384,17'd5916,17'd5918,17'd5918,17'd7999,17'd8629,17'd10513,17'd10777,17'd11181,17'd27932,17'd10515,17'd27815,17'd29592,17'd29592,17'd27933,17'd28183,17'd28183,17'd12160,17'd5334,17'd29884,17'd5327,17'd4686,17'd5330,17'd5336,17'd9091,17'd9933,17'd10515,17'd12160,17'd14048,17'd25085,17'd14301,17'd12906,17'd12467,17'd14301,17'd14301,17'd13800,17'd13169,17'd12165,17'd16850,17'd14303,17'd6561,17'd7182,17'd12167,17'd26115,17'd13172,17'd29601,17'd18860,17'd29885,17'd29886,17'd29887,17'd29888,17'd29889,17'd29890,17'd1235,17'd29891,17'd1679,17'd11337,17'd12644,17'd29609,17'd26966,17'd29892,17'd29611,17'd29892,17'd29038,17'd29170,17'd29170,17'd27708,17'd29170,17'd28793,17'd28792,17'd27583,17'd27583,17'd29893,17'd23651,17'd23651,17'd29894,17'd29895,17'd23306,17'd23479,17'd29614,17'd28658,17'd14737,17'd3079,17'd3230,17'd1535,17'd1536,17'd12916,17'd28318,17'd3581,17'd10389,17'd9662,17'd26343,17'd1683,17'd17423,17'd29896,17'd16140
},
'{
17'd8336,17'd8508,17'd10397,17'd10533,17'd4892,17'd29897,17'd27713,17'd4892,17'd3901,17'd2934,17'd2935,17'd2422,17'd1688,17'd4247,17'd1127,17'd4247,17'd1416,17'd17,17'd17,17'd17,17'd17,17'd1416,17'd17,17'd17,17'd653,17'd652,17'd7060,17'd7061,17'd7225,17'd7225,17'd7386,17'd7388,17'd6904,17'd6441,17'd28319,17'd28659,17'd27446,17'd29898,17'd5225,17'd5062,17'd6116,17'd5064,17'd25502,17'd29757,17'd29758,17'd3111,17'd2797,17'd29899,17'd22110,17'd29900,17'd29901,17'd29762,17'd25508,17'd18400,17'd24188,17'd29902,17'd23834,17'd25912,17'd29903,17'd28204,17'd16519,17'd16411,17'd14767,17'd14767,17'd16987,17'd16768,17'd16768,17'd16987,17'd15902,17'd17320,17'd19008,17'd19620,17'd19006,17'd20885,17'd29904,17'd17940,17'd14621,17'd14621,17'd14470,17'd16765,17'd18884,17'd17204,17'd16766,17'd20023,17'd29905,17'd10565,17'd8537,17'd6770,17'd10117,17'd10118,17'd9706,17'd9582,17'd9310,17'd9311,17'd9446,17'd9708,17'd18787,17'd9586,17'd18420,17'd16044,17'd7266,17'd13613,17'd29906,17'd29907,17'd29908,17'd29909,17'd29910,17'd29911,17'd29912,17'd29913,17'd29914,17'd29915,17'd29773,17'd29631,17'd29916,17'd29917,17'd15939,17'd11806,17'd11807,17'd14673,17'd11274,17'd10476,17'd16319,17'd29918,17'd29474,17'd29919,17'd29920,17'd29921,17'd16562,17'd9886,17'd8726,17'd9188,17'd17011,17'd14518,17'd16068,17'd11964,17'd13135,17'd18917,17'd19408,17'd24707,17'd27004,17'd28343,17'd28106,17'd27984,17'd25672,17'd29922,17'd29923,17'd29924,17'd29067,17'd29925,17'd29926,17'd28104,17'd20452,17'd19409,17'd18806,17'd13762,17'd12861,17'd13363,17'd12110,17'd12113,17'd14262,17'd10166,17'd18916,17'd9741,17'd11277,17'd19642,17'd10476,17'd11275,17'd14673,17'd11396,17'd11808,17'd11808,17'd11524,17'd11275,17'd10989,17'd13764,17'd13253,17'd16069,17'd10329,17'd9479,17'd8566,17'd15178,17'd9194,17'd10172,17'd29927,17'd29928,17'd27736,17'd27485,17'd29929,17'd29784,17'd28465,17'd29337,17'd29198,17'd29930,17'd29926,17'd29931,17'd29486,17'd18083,17'd18198,17'd29932,17'd22816,17'd22647,17'd11808,17'd13000,17'd13364,17'd12110,17'd18684,17'd29205,17'd29791,17'd29933,17'd29934,17'd29935,17'd29935,17'd29936,17'd29653,17'd29937,17'd17837,17'd29938,17'd10598,17'd29939,17'd29670,17'd29940,17'd10019,17'd29797,17'd29941,17'd10016,17'd29659,17'd29942,17'd29943,17'd29944,17'd29945,17'd29946,17'd29947,17'd29948,17'd29949,17'd29950,17'd29951,17'd29952,17'd29953,17'd29347,17'd29498,17'd29954,17'd29955,17'd29956,17'd29957,17'd29958,17'd29959,17'd29960,17'd29961,17'd29962,17'd29963,17'd29964,17'd29679,17'd29965,17'd29966,17'd29967,17'd29968,17'd29969,17'd25830,17'd25702,17'd26400,17'd25560,17'd26055,17'd25696,17'd25698,17'd25313,17'd25833,17'd29970,17'd28851,17'd29971,17'd23386,17'd29376,17'd29972,17'd24086,17'd29241,17'd23387,17'd29973,17'd29974,17'd29975,17'd29378,17'd29976,17'd25438,17'd25032,17'd23916,17'd29375,17'd23384,17'd24417,17'd28369,17'd27513,17'd27514,17'd28853,17'd27027,17'd26901,17'd28727,17'd29379,17'd29379,17'd29379,17'd29977,17'd28370,17'd29247,17'd29380,17'd29536,17'd29978,17'd29979,17'd29980,17'd29979,17'd29981,17'd29982,17'd29983,17'd29984,17'd29985,17'd29986,17'd29987,17'd29988,17'd29989,17'd29989,17'd29988,17'd29990,17'd26911,17'd29991,17'd29992,17'd29993,17'd29994,17'd29995,17'd29117,17'd28145,17'd29996,17'd25336,17'd28876,17'd29846,17'd29997,17'd27531,17'd29998,17'd28742,17'd29261,17'd28387,17'd26912,17'd26791,17'd26304,17'd28384,17'd29999,17'd30000,17'd30001,17'd30002,17'd30003,17'd30004,17'd24927,17'd30005,17'd30006,17'd30007,17'd19305,17'd30008,17'd30009,17'd30010,17'd30011,17'd30012,17'd30013,17'd30014,17'd30015,17'd30016,17'd30017,17'd30018,17'd30019,17'd30020,17'd30021,17'd29579,17'd30022,17'd30023,17'd29015,17'd28897,17'd30024,17'd30025,17'd30026,17'd21281,17'd30027,17'd22395,17'd23268,17'd23619,17'd30028,17'd24303,17'd25221,17'd11692,17'd10627,17'd7166,17'd6384,17'd5916,17'd5918,17'd5918,17'd7999,17'd8000,17'd9090,17'd10513,17'd27932,17'd27932,17'd10515,17'd27815,17'd29592,17'd29592,17'd27933,17'd27933,17'd28183,17'd11316,17'd6392,17'd30029,17'd30030,17'd4686,17'd5330,17'd5335,17'd6219,17'd7668,17'd10514,17'd12160,17'd11853,17'd11854,17'd11710,17'd13046,17'd12467,17'd12467,17'd12467,17'd13800,17'd13169,17'd12165,17'd30031,17'd14303,17'd30032,17'd7503,17'd12907,17'd30033,17'd22255,17'd18860,17'd29601,17'd30034,17'd30035,17'd30036,17'd30037,17'd30038,17'd30039,17'd30040,17'd30041,17'd1957,17'd5050,17'd14178,17'd2560,17'd26966,17'd29610,17'd29611,17'd29892,17'd29038,17'd29170,17'd29170,17'd27708,17'd29170,17'd28793,17'd28792,17'd27583,17'd27583,17'd30042,17'd30043,17'd30043,17'd30044,17'd29895,17'd23306,17'd23479,17'd23479,17'd29613,17'd14737,17'd2911,17'd3081,17'd1388,17'd1536,17'd30045,17'd12916,17'd3582,17'd3414,17'd4420,17'd2111,17'd592,17'd214,17'd30046,17'd16264
},
'{
17'd8335,17'd8508,17'd5198,17'd30047,17'd4244,17'd27713,17'd27713,17'd4428,17'd3901,17'd2934,17'd2935,17'd1831,17'd4247,17'd4247,17'd4247,17'd4247,17'd1416,17'd17,17'd17,17'd17,17'd1416,17'd1416,17'd4089,17'd3905,17'd653,17'd652,17'd7060,17'd7061,17'd7386,17'd7386,17'd7388,17'd7388,17'd6904,17'd6441,17'd28319,17'd28659,17'd27446,17'd5523,17'd6114,17'd12039,17'd6116,17'd30048,17'd25502,17'd30049,17'd29449,17'd29615,17'd30050,17'd30051,17'd30052,17'd29900,17'd30053,17'd25655,17'd30054,17'd24681,17'd24010,17'd30055,17'd30056,17'd30057,17'd29764,17'd21650,17'd24348,17'd16168,17'd14767,17'd14893,17'd16768,17'd16768,17'd16411,17'd16033,17'd17320,17'd17207,17'd19383,17'd19511,17'd20886,17'd30058,17'd29904,17'd13211,17'd14621,17'd14621,17'd14470,17'd12361,17'd12681,17'd17204,17'd16766,17'd18174,17'd20023,17'd10428,17'd8369,17'd6770,17'd30059,17'd24198,17'd9706,17'd9707,17'd9445,17'd9311,17'd9446,17'd9586,17'd18307,17'd9586,17'd9313,17'd8856,17'd29457,17'd7926,17'd28671,17'd29459,17'd30060,17'd30061,17'd30062,17'd30063,17'd30064,17'd29465,17'd30065,17'd30066,17'd30067,17'd10834,17'd30068,17'd10980,17'd11805,17'd13883,17'd11807,17'd14673,17'd14931,17'd10991,17'd25529,17'd30069,17'd8405,17'd29919,17'd25677,17'd30070,17'd8411,17'd9482,17'd15297,17'd13887,17'd11277,17'd13886,17'd16069,17'd11964,17'd12996,17'd17722,17'd23168,17'd24537,17'd27346,17'd28344,17'd28106,17'd28816,17'd29640,17'd28816,17'd30071,17'd30072,17'd30073,17'd30074,17'd28345,17'd27121,17'd30075,17'd12582,17'd13362,17'd11962,17'd20313,17'd13364,17'd11960,17'd16204,17'd10475,17'd21503,17'd11136,17'd12116,17'd11135,17'd11527,17'd11524,17'd11808,17'd16068,17'd11808,17'd10990,17'd11524,17'd11275,17'd11808,17'd11667,17'd13764,17'd14133,17'd12584,17'd9885,17'd9043,17'd11403,17'd11403,17'd8874,17'd24709,17'd28947,17'd30076,17'd30077,17'd27485,17'd29784,17'd29784,17'd30078,17'd29485,17'd30079,17'd29930,17'd30080,17'd30081,17'd30082,17'd21363,17'd30083,17'd14671,17'd14671,17'd13645,17'd11807,17'd13364,17'd12413,17'd12575,17'd18684,17'd29791,17'd29933,17'd30084,17'd30085,17'd30085,17'd30086,17'd30087,17'd30088,17'd30089,17'd30090,17'd30091,17'd30092,17'd10984,17'd30093,17'd10018,17'd10018,17'd10017,17'd10017,17'd30094,17'd30095,17'd30096,17'd30097,17'd30098,17'd30099,17'd30100,17'd30101,17'd30102,17'd30103,17'd30104,17'd30105,17'd30106,17'd29661,17'd30107,17'd30108,17'd30109,17'd30110,17'd30111,17'd30112,17'd30113,17'd30114,17'd30115,17'd30116,17'd29962,17'd30117,17'd30118,17'd30119,17'd30120,17'd30121,17'd30122,17'd30123,17'd30124,17'd30125,17'd29523,17'd25699,17'd25699,17'd26055,17'd25559,17'd25696,17'd25312,17'd26174,17'd28484,17'd30126,17'd29377,17'd29376,17'd30127,17'd23384,17'd24087,17'd23734,17'd30128,17'd30129,17'd22503,17'd23215,17'd29529,17'd24898,17'd25320,17'd25180,17'd23916,17'd29375,17'd23384,17'd24743,17'd28850,17'd27638,17'd26174,17'd28978,17'd27027,17'd26901,17'd28727,17'd29379,17'd29379,17'd29977,17'd29977,17'd28370,17'd28133,17'd28257,17'd29831,17'd30130,17'd30131,17'd30132,17'd29978,17'd29981,17'd29982,17'd29539,17'd30133,17'd30134,17'd30135,17'd30136,17'd29545,17'd29989,17'd29989,17'd29988,17'd29990,17'd27380,17'd30137,17'd30138,17'd30139,17'd29994,17'd30140,17'd30141,17'd28500,17'd27898,17'd30142,17'd28876,17'd29846,17'd25342,17'd28024,17'd27900,17'd26919,17'd28620,17'd30143,17'd27534,17'd27265,17'd30144,17'd30145,17'd30146,17'd30147,17'd30148,17'd30149,17'd30150,17'd30151,17'd30152,17'd30153,17'd30154,17'd30155,17'd30156,17'd19552,17'd30157,17'd30158,17'd30159,17'd19176,17'd30160,17'd30161,17'd30162,17'd30163,17'd30164,17'd30165,17'd30166,17'd30167,17'd30168,17'd30169,17'd30170,17'd30171,17'd30172,17'd30173,17'd30174,17'd30175,17'd30176,17'd30177,17'd30178,17'd21908,17'd22394,17'd23621,17'd23619,17'd30028,17'd25360,17'd11692,17'd10359,17'd7009,17'd5914,17'd6384,17'd5916,17'd5917,17'd5918,17'd7999,17'd8154,17'd9394,17'd10641,17'd10641,17'd10515,17'd10515,17'd27815,17'd27815,17'd29592,17'd27933,17'd28183,17'd11316,17'd30179,17'd30180,17'd30181,17'd4840,17'd5329,17'd5160,17'd6219,17'd7668,17'd10514,17'd12160,17'd11853,17'd11709,17'd11710,17'd13046,17'd13407,17'd13407,17'd12467,17'd13800,17'd30182,17'd12165,17'd12165,17'd7179,17'd30032,17'd7503,17'd12907,17'd30033,17'd30183,17'd24807,17'd29601,17'd30184,17'd30035,17'd30185,17'd30186,17'd29305,17'd30187,17'd30188,17'd30189,17'd1958,17'd2559,17'd2097,17'd2394,17'd2560,17'd27707,17'd29892,17'd28545,17'd28791,17'd29170,17'd27708,17'd27708,17'd27708,17'd29170,17'd28793,17'd28791,17'd28791,17'd30190,17'd30043,17'd29893,17'd23651,17'd30191,17'd5363,17'd23479,17'd29614,17'd30192,17'd2565,17'd2911,17'd3081,17'd1388,17'd13058,17'd30045,17'd12916,17'd3411,17'd10389,17'd23301,17'd26343,17'd180,17'd649,17'd30193,17'd30194
},
'{
17'd30195,17'd8508,17'd5375,17'd30047,17'd3902,17'd27713,17'd4243,17'd4428,17'd3901,17'd2934,17'd2935,17'd1831,17'd4247,17'd4247,17'd4247,17'd4247,17'd1416,17'd1416,17'd17,17'd17,17'd1416,17'd1416,17'd4089,17'd4089,17'd653,17'd652,17'd7060,17'd7061,17'd7386,17'd7386,17'd7388,17'd7556,17'd10408,17'd10672,17'd28319,17'd6442,17'd30196,17'd26974,17'd5525,17'd30197,17'd30198,17'd4097,17'd29757,17'd30049,17'd29449,17'd2954,17'd30199,17'd30200,17'd30201,17'd30202,17'd20728,17'd25655,17'd17800,17'd28436,17'd30203,17'd30204,17'd25911,17'd29622,17'd27834,17'd16289,17'd14219,17'd14768,17'd15384,17'd15641,17'd14768,17'd16987,17'd16033,17'd15902,17'd17320,17'd19008,17'd25512,17'd19382,17'd20885,17'd12815,17'd17096,17'd13211,17'd14621,17'd14621,17'd14622,17'd16658,17'd19006,17'd17204,17'd16766,17'd20023,17'd30205,17'd9574,17'd6142,17'd7412,17'd10118,17'd9580,17'd9582,17'd12822,17'd9445,17'd9446,17'd10701,17'd9708,17'd9446,17'd9312,17'd27836,17'd8855,17'd9021,17'd14490,17'd30206,17'd29051,17'd30207,17'd30208,17'd30209,17'd30210,17'd30211,17'd30212,17'd30213,17'd30066,17'd30214,17'd10586,17'd30215,17'd30216,17'd12999,17'd16325,17'd11521,17'd14810,17'd17236,17'd11670,17'd9338,17'd17230,17'd12722,17'd12424,17'd26259,17'd16562,17'd30217,17'd11672,17'd9045,17'd9345,17'd11135,17'd13001,17'd16069,17'd15185,17'd12582,17'd21671,17'd25925,17'd27004,17'd30218,17'd30071,17'd28344,17'd27346,17'd30219,17'd29328,17'd29067,17'd30220,17'd30221,17'd29198,17'd30222,17'd24537,17'd18197,17'd12422,17'd13362,17'd18805,17'd15564,17'd15564,17'd13646,17'd24029,17'd26152,17'd11136,17'd10992,17'd11671,17'd12863,17'd10476,17'd14931,17'd11274,17'd14673,17'd11130,17'd11399,17'd11524,17'd11275,17'd14673,17'd13253,17'd11667,17'd27350,17'd19779,17'd10173,17'd15941,17'd14675,17'd16067,17'd25145,17'd28821,17'd30223,17'd26873,17'd28228,17'd28465,17'd29784,17'd29784,17'd30224,17'd30225,17'd30226,17'd29926,17'd30227,17'd30228,17'd30229,17'd30230,17'd29789,17'd19533,17'd14671,17'd16204,17'd13363,17'd12413,17'd12855,17'd16799,17'd30231,17'd30232,17'd30233,17'd30234,17'd30085,17'd30235,17'd30236,17'd30088,17'd30237,17'd30238,17'd30239,17'd30240,17'd24701,17'd10984,17'd10728,17'd10727,17'd30094,17'd10013,17'd29496,17'd30241,17'd30242,17'd30243,17'd30244,17'd30245,17'd30246,17'd30247,17'd30248,17'd30249,17'd30250,17'd30251,17'd30252,17'd30253,17'd30254,17'd30255,17'd30256,17'd29222,17'd30257,17'd30258,17'd30259,17'd30260,17'd30261,17'd30115,17'd30262,17'd30263,17'd30264,17'd30265,17'd30266,17'd30267,17'd30268,17'd30269,17'd30270,17'd30271,17'd30272,17'd30273,17'd29523,17'd25701,17'd29524,17'd30274,17'd25553,17'd25429,17'd27515,17'd28130,17'd25032,17'd29243,17'd23918,17'd29241,17'd30275,17'd29375,17'd30127,17'd23217,17'd22859,17'd30276,17'd30277,17'd30278,17'd24743,17'd27637,17'd29976,17'd24742,17'd29534,17'd23384,17'd29100,17'd29103,17'd28598,17'd25949,17'd28978,17'd27027,17'd26901,17'd28727,17'd29379,17'd29379,17'd30279,17'd30279,17'd28370,17'd29247,17'd29380,17'd29831,17'd30130,17'd30280,17'd30132,17'd30131,17'd29981,17'd30281,17'd30282,17'd30283,17'd30284,17'd30285,17'd30286,17'd30287,17'd29989,17'd29989,17'd30288,17'd30289,17'd30290,17'd30137,17'd30291,17'd30292,17'd24251,17'd30293,17'd30294,17'd28736,17'd28614,17'd30295,17'd25448,17'd28876,17'd29846,17'd25342,17'd28024,17'd27531,17'd28620,17'd30296,17'd28027,17'd26296,17'd27270,17'd30297,17'd30146,17'd30298,17'd30299,17'd30300,17'd30301,17'd30302,17'd21716,17'd30303,17'd30304,17'd30305,17'd30306,17'd30307,17'd25742,17'd24451,17'd30308,17'd30309,17'd30310,17'd30311,17'd30312,17'd30313,17'd30314,17'd30315,17'd30316,17'd30317,17'd30318,17'd30319,17'd30320,17'd30321,17'd30023,17'd30322,17'd30323,17'd30324,17'd30325,17'd30326,17'd30327,17'd30328,17'd23271,17'd23097,17'd30329,17'd29883,17'd24474,17'd22413,17'd30330,17'd30331,17'd6844,17'd5914,17'd5916,17'd5916,17'd5918,17'd5918,17'd6707,17'd9090,17'd10777,17'd10641,17'd10515,17'd10515,17'd27815,17'd27815,17'd29592,17'd27933,17'd28183,17'd11037,17'd30332,17'd5615,17'd30181,17'd4995,17'd5329,17'd30333,17'd5614,17'd6391,17'd10514,17'd30332,17'd11431,17'd11709,17'd29161,17'd12905,17'd13407,17'd13166,17'd12760,17'd13800,17'd30182,17'd29597,17'd29597,17'd8155,17'd14303,17'd7330,17'd16739,17'd30334,17'd30335,17'd20855,17'd29601,17'd30184,17'd30336,17'd30337,17'd30338,17'd29305,17'd30339,17'd30340,17'd30341,17'd30342,17'd2739,17'd7210,17'd1383,17'd1672,17'd29037,17'd29610,17'd28545,17'd28791,17'd29170,17'd27708,17'd27708,17'd27708,17'd29170,17'd28793,17'd28791,17'd28791,17'd30190,17'd29893,17'd30042,17'd23651,17'd30343,17'd23479,17'd29895,17'd29895,17'd24166,17'd24500,17'd2747,17'd1387,17'd1389,17'd13421,17'd13057,17'd30045,17'd3411,17'd3239,17'd4421,17'd8950,17'd213,17'd20001,17'd30344,17'd30345
},
'{
17'd30346,17'd8508,17'd6422,17'd5199,17'd4426,17'd4891,17'd3902,17'd4244,17'd3901,17'd2934,17'd3252,17'd1831,17'd4247,17'd4247,17'd1688,17'd4247,17'd1416,17'd1416,17'd17,17'd17,17'd1416,17'd1416,17'd2938,17'd2938,17'd1278,17'd980,17'd20570,17'd7385,17'd7386,17'd7386,17'd7388,17'd6600,17'd6441,17'd6112,17'd6442,17'd27446,17'd29898,17'd5664,17'd6115,17'd30347,17'd30048,17'd4097,17'd30348,17'd3269,17'd30349,17'd30350,17'd30351,17'd30352,17'd30353,17'd26982,17'd20728,17'd5071,17'd30354,17'd18402,17'd30355,17'd24683,17'd25912,17'd29764,17'd16986,17'd17319,17'd14347,17'd14626,17'd15384,17'd14892,17'd17321,17'd16033,17'd15902,17'd15902,17'd17320,17'd19383,17'd18655,17'd18884,17'd30058,17'd17940,17'd19005,17'd15383,17'd14621,17'd14621,17'd14622,17'd16658,17'd17204,17'd16766,17'd17205,17'd18174,17'd30356,17'd9573,17'd7412,17'd7412,17'd24198,17'd9706,17'd9707,17'd9444,17'd10126,17'd10292,17'd18897,17'd17947,17'd9446,17'd10701,17'd9313,17'd7266,17'd13613,17'd30357,17'd30358,17'd30359,17'd30207,17'd30360,17'd30361,17'd30362,17'd28933,17'd30363,17'd30364,17'd30365,17'd30366,17'd30367,17'd30368,17'd28566,17'd12113,17'd18917,17'd11395,17'd14931,17'd10605,17'd9739,17'd11529,17'd19159,17'd12722,17'd23517,17'd24368,17'd8412,17'd15296,17'd20176,17'd9189,17'd9885,17'd11527,17'd13138,17'd16068,17'd15185,17'd15053,17'd16324,17'd25927,17'd28816,17'd28344,17'd29328,17'd28343,17'd27346,17'd30369,17'd30370,17'd29785,17'd30371,17'd30372,17'd30373,17'd27121,17'd22819,17'd12582,17'd12262,17'd11962,17'd21204,17'd15564,17'd13764,17'd11396,17'd11669,17'd10992,17'd9341,17'd9741,17'd11135,17'd11527,17'd13886,17'd14810,17'd14673,17'd11808,17'd11808,17'd11399,17'd11399,17'd11274,17'd11666,17'd11962,17'd16068,17'd11401,17'd10334,17'd9348,17'd15568,17'd8727,17'd9189,17'd17842,17'd30374,17'd28570,17'd27857,17'd28465,17'd28465,17'd28465,17'd30224,17'd30226,17'd30375,17'd30226,17'd30376,17'd30377,17'd25670,17'd23513,17'd22816,17'd11130,17'd11129,17'd12262,17'd12857,17'd12256,17'd14523,17'd14523,17'd30378,17'd30231,17'd30379,17'd29934,17'd29936,17'd30236,17'd30380,17'd30381,17'd30382,17'd30383,17'd30384,17'd30385,17'd10982,17'd24990,17'd30386,17'd29917,17'd30387,17'd30388,17'd30389,17'd30242,17'd30390,17'd30391,17'd30392,17'd30393,17'd30394,17'd30394,17'd30395,17'd30396,17'd30397,17'd30398,17'd30399,17'd30400,17'd30401,17'd30402,17'd30403,17'd30404,17'd30405,17'd30406,17'd30407,17'd30408,17'd30409,17'd30410,17'd30411,17'd30412,17'd30413,17'd30414,17'd30415,17'd30416,17'd30417,17'd30418,17'd30419,17'd30420,17'd30421,17'd30271,17'd30272,17'd30125,17'd30273,17'd30422,17'd30423,17'd27369,17'd26167,17'd27515,17'd28130,17'd25031,17'd24902,17'd23733,17'd23920,17'd30275,17'd30424,17'd23736,17'd30425,17'd30426,17'd30427,17'd30428,17'd30429,17'd30430,17'd29548,17'd29976,17'd24742,17'd30431,17'd29972,17'd29102,17'd30432,17'd28597,17'd25949,17'd28978,17'd27027,17'd26901,17'd28727,17'd29379,17'd29379,17'd30279,17'd30279,17'd28370,17'd29247,17'd29380,17'd29536,17'd30130,17'd30280,17'd30433,17'd30280,17'd29981,17'd30434,17'd30435,17'd30436,17'd30437,17'd30438,17'd30286,17'd30439,17'd29989,17'd30440,17'd30441,17'd30442,17'd30290,17'd30443,17'd30444,17'd30445,17'd30446,17'd29102,17'd29994,17'd30447,17'd30448,17'd30449,17'd27159,17'd27042,17'd26075,17'd25853,17'd30450,17'd27387,17'd30451,17'd28386,17'd26793,17'd30452,17'd29698,17'd30453,17'd30136,17'd30454,17'd30455,17'd30456,17'd25952,17'd30457,17'd30458,17'd30459,17'd30460,17'd25063,17'd30461,17'd29129,17'd30462,17'd30463,17'd24452,17'd30464,17'd30465,17'd30466,17'd30467,17'd30468,17'd30469,17'd21529,17'd30470,17'd30471,17'd30472,17'd30473,17'd29873,17'd30474,17'd30475,17'd30476,17'd30477,17'd30478,17'd30479,17'd30480,17'd30481,17'd30482,17'd22068,17'd22065,17'd22567,17'd30483,17'd30484,17'd25877,17'd26448,17'd7165,17'd6212,17'd6383,17'd6384,17'd23630,17'd5760,17'd5332,17'd6553,17'd8154,17'd10513,17'd10777,17'd27932,17'd27932,17'd10515,17'd27815,17'd29592,17'd27933,17'd27933,17'd28183,17'd11037,17'd30179,17'd30485,17'd30486,17'd5005,17'd30333,17'd27935,17'd5919,17'd30487,17'd30332,17'd11181,17'd28534,17'd30488,17'd11710,17'd13166,17'd13166,17'd12760,17'd13800,17'd11038,17'd10779,17'd29432,17'd8155,17'd14303,17'd7330,17'd30489,17'd30490,17'd30491,17'd17072,17'd29601,17'd30492,17'd30493,17'd30494,17'd30495,17'd29305,17'd30496,17'd30497,17'd30498,17'd29749,17'd627,17'd2559,17'd2575,17'd2394,17'd29037,17'd29610,17'd28545,17'd27710,17'd29170,17'd27708,17'd27708,17'd27708,17'd29170,17'd28793,17'd28793,17'd28793,17'd30190,17'd29893,17'd30042,17'd30043,17'd30343,17'd23479,17'd30191,17'd2910,17'd30499,17'd24499,17'd2744,17'd1387,17'd1389,17'd13421,17'd13057,17'd30045,17'd27712,17'd19732,17'd30500,17'd20867,17'd280,17'd29173,17'd30344,17'd398
},
'{
17'd30501,17'd8336,17'd6422,17'd6421,17'd5646,17'd4891,17'd3902,17'd3902,17'd3901,17'd2934,17'd3252,17'd1831,17'd4247,17'd4247,17'd1688,17'd1831,17'd1414,17'd1416,17'd17,17'd17,17'd1416,17'd1416,17'd2938,17'd2938,17'd1278,17'd980,17'd20570,17'd7385,17'd7386,17'd7386,17'd7388,17'd6600,17'd10672,17'd6112,17'd6442,17'd30196,17'd5523,17'd5664,17'd6115,17'd30502,17'd30048,17'd30348,17'd30503,17'd12790,17'd30504,17'd30505,17'd22790,17'd30506,17'd29044,17'd28435,17'd20415,17'd30507,17'd30508,17'd18288,17'd24342,17'd30509,17'd30057,17'd30510,17'd21185,17'd24348,17'd16168,17'd15384,17'd16029,17'd14766,17'd17321,17'd16033,17'd15902,17'd17445,17'd19008,17'd28668,17'd30511,17'd20885,17'd17940,17'd17940,17'd19005,17'd15383,17'd14764,17'd14621,17'd14622,17'd16658,17'd19893,17'd16766,17'd18174,17'd20023,17'd12682,17'd9701,17'd7412,17'd7581,17'd9579,17'd9581,17'd9309,17'd9445,17'd10292,17'd10292,17'd18897,17'd17947,17'd10701,17'd10701,17'd9167,17'd13222,17'd9022,17'd29906,17'd29907,17'd30512,17'd30513,17'd30514,17'd30515,17'd30516,17'd30517,17'd30518,17'd30519,17'd30365,17'd30520,17'd30521,17'd30092,17'd12999,17'd13883,17'd19158,17'd14673,17'd10605,17'd26037,17'd17011,17'd16910,17'd30522,17'd22473,17'd8730,17'd15429,17'd9744,17'd30523,17'd9348,17'd10335,17'd10024,17'd15176,17'd11274,17'd11964,17'd15185,17'd11959,17'd25670,17'd26370,17'd28943,17'd30370,17'd29066,17'd30524,17'd30525,17'd30526,17'd30527,17'd30221,17'd30528,17'd29648,17'd28572,17'd24856,17'd20314,17'd19158,17'd13762,17'd12861,17'd23854,17'd18679,17'd11666,17'd11399,17'd26152,17'd9480,17'd9480,17'd11277,17'd20756,17'd11132,17'd11399,17'd11274,17'd11274,17'd11130,17'd11274,17'd11399,17'd21206,17'd16068,17'd13137,17'd11520,17'd14931,17'd15566,17'd17480,17'd30523,17'd11137,17'd8881,17'd17470,17'd13367,17'd30529,17'd27485,17'd28572,17'd28465,17'd28351,17'd28945,17'd29642,17'd30530,17'd30531,17'd29485,17'd29486,17'd28693,17'd22472,17'd30532,17'd11398,17'd10990,17'd20451,17'd12861,17'd12257,17'd16799,17'd30231,17'd30533,17'd30534,17'd30379,17'd29792,17'd29339,17'd29653,17'd30535,17'd30381,17'd30536,17'd30537,17'd30538,17'd30539,17'd10979,17'd24990,17'd10984,17'd10158,17'd30094,17'd30540,17'd30541,17'd30542,17'd29802,17'd30543,17'd30544,17'd30545,17'd30546,17'd30547,17'd30548,17'd30549,17'd30550,17'd30398,17'd30551,17'd30400,17'd30552,17'd30553,17'd30402,17'd30554,17'd30555,17'd30556,17'd30557,17'd30558,17'd30559,17'd30560,17'd30561,17'd30562,17'd30563,17'd30564,17'd30414,17'd30565,17'd30566,17'd30567,17'd30568,17'd30569,17'd30570,17'd30571,17'd30572,17'd30573,17'd30574,17'd30575,17'd30576,17'd30423,17'd30577,17'd25696,17'd26903,17'd28594,17'd25179,17'd29100,17'd23732,17'd30275,17'd28849,17'd30578,17'd30579,17'd30129,17'd22159,17'd30580,17'd30581,17'd30582,17'd30583,17'd30584,17'd25031,17'd24742,17'd24249,17'd29377,17'd30585,17'd25031,17'd27882,17'd26062,17'd28724,17'd27258,17'd30586,17'd28727,17'd29379,17'd29246,17'd27885,17'd30279,17'd28370,17'd29247,17'd30587,17'd29690,17'd30280,17'd30280,17'd30433,17'd30280,17'd29981,17'd30434,17'd30588,17'd30589,17'd30590,17'd30591,17'd30286,17'd30592,17'd29700,17'd30440,17'd30593,17'd30442,17'd30297,17'd30443,17'd30594,17'd30595,17'd30446,17'd30596,17'd30597,17'd30598,17'd28268,17'd24601,17'd30599,17'd25189,17'd30600,17'd27044,17'd27530,17'd27391,17'd30601,17'd30602,17'd29394,17'd26669,17'd30290,17'd30603,17'd30136,17'd30604,17'd30605,17'd30606,17'd25436,17'd30598,17'd30607,17'd30608,17'd30609,17'd19942,17'd30610,17'd30611,17'd30612,17'd30613,17'd30614,17'd30615,17'd30616,17'd30617,17'd30618,17'd30619,17'd30620,17'd30621,17'd30622,17'd30623,17'd30624,17'd30625,17'd30626,17'd30627,17'd30628,17'd30629,17'd30475,17'd30477,17'd30630,17'd30631,17'd30632,17'd30633,17'd30634,17'd22064,17'd22740,17'd22567,17'd30635,17'd24642,17'd30636,17'd10197,17'd6842,17'd6382,17'd6384,17'd23630,17'd5760,17'd5760,17'd6387,17'd6707,17'd9394,17'd10777,17'd27932,17'd11181,17'd10515,17'd27815,17'd27933,17'd27933,17'd27933,17'd28183,17'd27934,17'd30332,17'd5328,17'd29595,17'd30637,17'd30638,17'd5336,17'd5615,17'd28058,17'd10515,17'd28306,17'd28305,17'd30639,17'd29161,17'd13166,17'd14166,17'd11854,17'd13800,17'd10642,17'd10516,17'd29432,17'd8155,17'd7179,17'd7330,17'd30640,17'd30641,17'd30642,17'd13567,17'd29601,17'd30643,17'd9528,17'd27574,17'd30644,17'd30645,17'd30646,17'd30647,17'd30648,17'd26338,17'd234,17'd1680,17'd412,17'd779,17'd3223,17'd29892,17'd27581,17'd30649,17'd29170,17'd29170,17'd27708,17'd27708,17'd29170,17'd29170,17'd28793,17'd28793,17'd30650,17'd30042,17'd30042,17'd30043,17'd30651,17'd29895,17'd30191,17'd30043,17'd27582,17'd24499,17'd2744,17'd2752,17'd1252,17'd13421,17'd13178,17'd13057,17'd27712,17'd8642,17'd30652,17'd30653,17'd280,17'd20266,17'd586,17'd398
},
'{
17'd30346,17'd7882,17'd6422,17'd6421,17'd5201,17'd4426,17'd4891,17'd4244,17'd3901,17'd3101,17'd1831,17'd4247,17'd15745,17'd2594,17'd1831,17'd4247,17'd1416,17'd1416,17'd1416,17'd1416,17'd4089,17'd4089,17'd2938,17'd653,17'd980,17'd27,17'd7385,17'd7555,17'd7388,17'd7388,17'd7389,17'd6600,17'd27592,17'd6280,17'd5812,17'd30196,17'd26974,17'd5525,17'd5665,17'd26014,17'd25903,17'd30654,17'd3920,17'd3269,17'd30504,17'd23660,17'd16267,17'd29308,17'd30655,17'd28435,17'd20282,17'd14878,17'd18048,17'd14998,17'd24682,17'd30656,17'd29903,17'd27834,17'd16289,17'd16169,17'd16881,17'd14767,17'd14892,17'd14893,17'd16987,17'd16033,17'd17320,17'd16519,17'd19255,17'd19620,17'd19382,17'd30058,17'd30657,17'd15383,17'd19890,17'd13599,17'd13211,17'd14621,17'd12362,17'd19006,17'd21649,17'd16410,17'd20023,17'd10944,17'd9701,17'd8536,17'd30658,17'd30659,17'd9705,17'd9581,17'd9583,17'd9584,17'd10292,17'd10292,17'd18897,17'd17947,17'd30660,17'd18420,17'd8855,17'd7925,17'd8081,17'd28671,17'd28208,17'd30661,17'd30662,17'd30663,17'd30664,17'd30665,17'd30666,17'd30667,17'd28564,17'd30520,17'd30668,17'd30669,17'd30670,17'd14002,17'd12113,17'd11807,17'd14931,17'd10477,17'd19642,17'd15187,17'd15179,17'd30671,17'd30672,17'd8574,17'd8413,17'd18201,17'd14675,17'd9348,17'd15807,17'd11135,17'd13886,17'd11808,17'd11964,17'd13883,17'd16324,17'd26036,17'd26757,17'd30673,17'd30370,17'd30674,17'd30524,17'd30370,17'd30675,17'd30676,17'd30677,17'd30678,17'd28467,17'd27234,17'd23168,17'd16442,17'd18444,17'd11806,17'd12718,17'd12857,17'd11962,17'd16068,17'd12863,17'd10992,17'd9620,17'd9479,17'd11277,17'd11528,17'd13886,17'd14810,17'd11274,17'd22647,17'd21206,17'd11524,17'd21206,17'd17236,17'd15182,17'd12862,17'd14810,17'd10326,17'd22814,17'd8726,17'd14135,17'd19535,17'd15682,17'd14668,17'd27861,17'd27858,17'd30078,17'd30679,17'd28690,17'd28351,17'd29780,17'd30372,17'd30680,17'd30681,17'd29787,17'd17971,17'd20314,17'd30083,17'd24029,17'd11399,17'd10990,17'd11520,17'd30682,17'd12576,17'd30378,17'd30683,17'd30232,17'd30232,17'd29792,17'd29792,17'd30684,17'd30685,17'd30686,17'd30687,17'd30537,17'd30688,17'd30689,17'd11516,17'd30690,17'd30691,17'd11271,17'd29658,17'd30692,17'd29349,17'd29800,17'd30693,17'd30694,17'd30695,17'd30696,17'd30697,17'd30698,17'd30699,17'd30700,17'd30551,17'd30701,17'd30702,17'd30703,17'd30704,17'd30552,17'd29349,17'd30705,17'd30706,17'd30707,17'd30708,17'd30709,17'd30710,17'd30711,17'd30712,17'd30713,17'd30714,17'd30715,17'd30716,17'd30716,17'd30717,17'd30718,17'd30719,17'd30720,17'd30721,17'd30722,17'd30723,17'd30724,17'd30572,17'd30725,17'd30575,17'd30726,17'd30423,17'd27369,17'd25696,17'd28978,17'd28720,17'd25030,17'd24415,17'd24086,17'd30275,17'd24902,17'd29528,17'd23215,17'd22680,17'd22162,17'd30727,17'd30728,17'd30729,17'd30730,17'd30731,17'd28851,17'd24416,17'd29534,17'd30275,17'd30732,17'd30733,17'd25317,17'd30734,17'd25707,17'd27258,17'd27027,17'd30735,17'd29245,17'd27642,17'd30279,17'd29977,17'd28370,17'd29247,17'd30587,17'd28857,17'd30130,17'd30736,17'd30737,17'd30737,17'd30738,17'd30739,17'd30740,17'd30741,17'd30742,17'd30743,17'd30744,17'd30745,17'd30746,17'd29700,17'd30288,17'd30747,17'd29698,17'd30748,17'd30749,17'd30750,17'd30446,17'd30596,17'd30751,17'd30752,17'd30753,17'd28985,17'd24910,17'd29390,17'd30754,17'd26183,17'd27782,17'd27391,17'd30601,17'd28273,17'd30143,17'd30755,17'd30756,17'd30757,17'd30758,17'd30604,17'd30759,17'd28481,17'd28597,17'd29256,17'd30760,17'd30761,17'd30762,17'd30763,17'd30764,17'd30765,17'd30766,17'd30767,17'd30768,17'd30769,17'd30770,17'd30771,17'd30772,17'd30773,17'd30774,17'd30775,17'd30776,17'd30777,17'd30778,17'd30779,17'd30780,17'd30781,17'd30782,17'd30476,17'd30783,17'd30784,17'd30785,17'd30786,17'd30787,17'd30788,17'd30789,17'd21747,17'd30790,17'd30791,17'd30792,17'd30793,17'd25768,17'd26449,17'd6212,17'd6212,17'd5759,17'd26328,17'd5482,17'd5482,17'd6387,17'd6707,17'd9090,17'd9394,17'd10641,17'd11576,17'd10642,17'd27815,17'd29592,17'd27933,17'd28057,17'd29592,17'd29158,17'd11316,17'd30794,17'd30795,17'd30796,17'd30333,17'd5336,17'd26949,17'd28058,17'd10514,17'd11431,17'd28305,17'd11431,17'd11710,17'd13166,17'd14166,17'd11577,17'd11316,17'd10515,17'd10516,17'd10779,17'd8155,17'd7179,17'd6712,17'd7183,17'd17410,17'd30797,17'd30798,17'd24807,17'd30799,17'd4044,17'd30800,17'd30801,17'd30802,17'd30803,17'd30804,17'd30805,17'd30806,17'd245,17'd232,17'd7210,17'd2098,17'd5777,17'd29037,17'd27581,17'd27710,17'd27708,17'd29610,17'd27708,17'd27708,17'd27708,17'd29170,17'd29170,17'd28793,17'd30807,17'd5499,17'd30650,17'd30043,17'd30042,17'd23651,17'd30191,17'd28431,17'd24500,17'd24499,17'd14738,17'd1386,17'd1390,17'd1391,17'd30045,17'd13057,17'd20401,17'd30808,17'd30500,17'd30653,17'd280,17'd15742,17'd30809,17'd30810
},
'{
17'd30346,17'd7882,17'd6422,17'd6421,17'd5201,17'd4426,17'd4891,17'd4892,17'd3427,17'd3101,17'd1831,17'd4247,17'd15745,17'd2594,17'd1688,17'd1688,17'd1414,17'd1416,17'd1416,17'd1416,17'd4089,17'd4089,17'd653,17'd653,17'd980,17'd27,17'd7385,17'd7555,17'd7388,17'd7388,17'd7389,17'd6600,17'd27592,17'd6280,17'd5812,17'd5385,17'd5664,17'd5525,17'd5665,17'd30198,17'd4261,17'd30811,17'd30812,17'd30813,17'd2954,17'd22970,17'd30814,17'd1991,17'd30815,17'd30816,17'd25796,17'd30817,17'd18526,17'd15374,17'd24517,17'd30818,17'd30819,17'd21650,17'd15899,17'd16411,17'd14767,17'd14892,17'd14892,17'd14892,17'd16987,17'd15902,17'd17320,17'd17319,17'd18656,17'd18655,17'd19006,17'd12815,17'd23325,17'd19005,17'd13210,17'd19005,17'd14764,17'd12361,17'd16658,17'd19006,17'd21649,17'd16164,17'd15765,17'd21967,17'd7250,17'd7086,17'd8685,17'd9705,17'd30820,17'd9582,17'd9583,17'd9584,17'd10292,17'd10292,17'd18897,17'd17947,17'd29456,17'd15537,17'd7266,17'd9021,17'd7594,17'd28671,17'd28208,17'd28209,17'd28210,17'd30821,17'd30822,17'd30823,17'd30824,17'd30825,17'd28564,17'd30366,17'd30826,17'd30827,17'd30216,17'd12858,17'd13135,17'd11964,17'd10990,17'd10478,17'd15431,17'd15944,17'd30522,17'd8409,17'd8575,17'd8573,17'd25147,17'd12724,17'd8409,17'd8721,17'd9479,17'd12585,17'd11524,17'd11397,17'd19158,17'd11959,17'd30828,17'd28570,17'd28106,17'd30829,17'd30370,17'd30830,17'd30831,17'd30832,17'd30833,17'd30834,17'd30677,17'd29930,17'd28350,17'd18200,17'd11959,17'd16442,17'd19158,17'd11961,17'd13882,17'd11961,17'd11807,17'd10990,17'd9883,17'd9620,17'd9479,17'd16549,17'd11135,17'd10991,17'd10990,17'd14931,17'd11808,17'd11130,17'd11399,17'd11399,17'd11399,17'd17838,17'd15182,17'd24860,17'd13886,17'd12116,17'd9041,17'd18201,17'd12865,17'd30671,17'd10025,17'd30835,17'd28570,17'd28467,17'd30836,17'd30836,17'd28465,17'd28466,17'd29930,17'd29785,17'd29647,17'd30225,17'd27484,17'd15434,17'd18681,17'd30532,17'd11274,17'd10990,17'd14810,17'd30837,17'd15686,17'd18684,17'd30838,17'd30838,17'd30839,17'd30840,17'd29934,17'd29651,17'd30685,17'd30841,17'd30842,17'd30843,17'd30844,17'd30845,17'd30846,17'd26146,17'd30847,17'd30848,17'd30849,17'd30692,17'd29350,17'd30850,17'd30851,17'd30852,17'd30696,17'd30696,17'd30853,17'd30854,17'd30855,17'd30856,17'd30857,17'd30551,17'd30702,17'd30858,17'd30859,17'd30860,17'd29662,17'd30104,17'd30861,17'd30862,17'd30863,17'd30864,17'd30865,17'd30866,17'd30867,17'd30868,17'd30869,17'd30870,17'd30871,17'd30872,17'd30873,17'd30874,17'd30875,17'd30719,17'd30720,17'd30876,17'd30877,17'd30878,17'd30123,17'd30572,17'd30573,17'd30574,17'd30726,17'd30423,17'd27369,17'd26167,17'd28724,17'd28720,17'd25030,17'd24743,17'd30879,17'd23564,17'd24086,17'd29528,17'd29973,17'd22856,17'd22861,17'd30880,17'd23220,17'd30881,17'd30882,17'd30883,17'd23916,17'd23916,17'd24249,17'd30275,17'd29529,17'd29688,17'd28850,17'd30734,17'd25707,17'd27258,17'd27027,17'd28727,17'd29246,17'd27642,17'd30279,17'd30279,17'd28370,17'd29247,17'd30587,17'd30884,17'd30280,17'd30736,17'd30737,17'd30736,17'd30885,17'd30739,17'd30434,17'd29983,17'd30886,17'd30887,17'd30888,17'd30888,17'd30889,17'd30889,17'd30890,17'd30747,17'd30891,17'd27377,17'd30892,17'd30893,17'd24250,17'd30894,17'd30596,17'd30895,17'd30002,17'd30896,17'd30897,17'd26080,17'd28739,17'd25730,17'd26547,17'd27661,17'd30451,17'd30451,17'd29555,17'd30898,17'd30899,17'd30900,17'd30901,17'd30604,17'd30902,17'd26062,17'd28599,17'd30903,17'd30904,17'd30905,17'd22700,17'd30906,17'd30907,17'd30908,17'd30909,17'd20201,17'd30910,17'd30911,17'd30912,17'd30913,17'd30914,17'd30915,17'd30916,17'd30917,17'd30918,17'd30919,17'd30920,17'd30921,17'd30922,17'd30923,17'd30924,17'd30925,17'd30926,17'd30927,17'd30928,17'd30929,17'd30930,17'd30931,17'd30932,17'd30634,17'd22063,17'd22064,17'd22222,17'd22932,17'd25878,17'd10196,17'd23799,17'd6382,17'd5759,17'd26328,17'd5482,17'd5481,17'd5332,17'd6218,17'd9090,17'd9394,17'd10641,17'd11576,17'd10642,17'd27815,17'd29592,17'd27933,17'd27933,17'd30933,17'd30934,17'd28057,17'd30935,17'd28905,17'd30936,17'd25627,17'd5333,17'd26949,17'd6391,17'd27815,17'd28305,17'd28305,17'd11181,17'd29161,17'd13166,17'd14049,17'd11316,17'd11316,17'd10515,17'd27815,17'd10516,17'd10517,17'd7179,17'd30937,17'd7841,17'd30489,17'd26001,17'd23983,17'd19352,17'd30799,17'd4548,17'd30938,17'd30939,17'd30940,17'd30803,17'd30941,17'd30805,17'd30806,17'd239,17'd233,17'd2905,17'd7027,17'd7682,17'd30942,17'd27708,17'd27710,17'd27708,17'd29610,17'd27708,17'd27708,17'd27708,17'd27708,17'd29170,17'd29170,17'd27711,17'd30807,17'd30650,17'd29893,17'd30042,17'd30043,17'd30343,17'd30043,17'd26722,17'd24499,17'd24667,17'd2568,17'd1390,17'd18272,17'd1392,17'd13178,17'd20401,17'd30943,17'd30944,17'd594,17'd1543,17'd29753,17'd30945,17'd30946
},
'{
17'd30947,17'd7883,17'd6422,17'd5053,17'd4735,17'd4426,17'd4891,17'd4892,17'd3427,17'd14070,17'd1831,17'd4247,17'd2595,17'd2594,17'd1688,17'd1688,17'd1414,17'd1414,17'd1416,17'd1416,17'd1416,17'd1416,17'd653,17'd653,17'd27444,17'd7060,17'd7385,17'd7555,17'd7388,17'd7388,17'd6600,17'd6441,17'd30948,17'd5812,17'd30196,17'd26974,17'd5225,17'd6284,17'd6116,17'd30198,17'd4261,17'd30811,17'd30812,17'd30949,17'd2798,17'd29899,17'd30950,17'd21796,17'd30951,17'd30952,17'd4910,17'd14757,17'd18402,17'd30953,17'd30954,17'd30955,17'd30956,17'd19255,17'd16034,17'd16168,17'd14767,17'd14892,17'd17208,17'd16987,17'd17448,17'd17320,17'd17319,17'd17319,17'd18656,17'd17941,17'd12531,17'd17940,17'd17809,17'd13210,17'd19005,17'd15383,17'd14891,17'd13969,17'd12532,17'd17689,17'd16164,17'd30957,17'd14222,17'd13847,17'd30958,17'd7580,17'd30659,17'd9705,17'd9846,17'd9707,17'd9444,17'd9584,17'd10292,17'd10292,17'd18897,17'd17947,17'd30959,17'd17581,17'd29457,17'd13613,17'd7594,17'd8082,17'd28328,17'd30960,17'd30961,17'd30962,17'd30963,17'd30964,17'd29190,17'd30364,17'd30965,17'd28336,17'd30966,17'd30967,17'd30968,17'd12858,17'd11963,17'd10989,17'd10739,17'd20756,17'd28578,17'd8873,17'd30969,17'd8572,17'd8575,17'd8413,17'd14135,17'd30970,17'd20453,17'd9188,17'd16549,17'd12863,17'd11524,17'd13516,17'd18917,17'd16324,17'd27736,17'd28229,17'd30829,17'd30971,17'd30071,17'd29066,17'd29067,17'd30972,17'd30834,17'd30973,17'd30974,17'd29201,17'd26373,17'd12108,17'd15053,17'd16204,17'd13135,17'd11961,17'd13761,17'd11806,17'd11274,17'd19532,17'd9885,17'd9620,17'd16549,17'd22131,17'd11528,17'd10477,17'd10990,17'd11275,17'd11399,17'd11399,17'd11399,17'd21206,17'd10990,17'd15182,17'd14803,17'd10477,17'd10479,17'd9344,17'd8410,17'd18808,17'd12723,17'd8720,17'd14668,17'd30975,17'd27857,17'd30976,17'd30977,17'd30978,17'd30836,17'd29926,17'd29785,17'd29785,17'd29647,17'd30979,17'd16685,17'd18917,17'd30980,17'd19533,17'd11275,17'd14931,17'd18805,17'd30981,17'd30982,17'd30983,17'd30232,17'd30839,17'd30233,17'd30234,17'd30087,17'd30984,17'd30985,17'd30986,17'd30987,17'd30988,17'd30989,17'd30990,17'd26146,17'd30991,17'd30992,17'd30552,17'd30993,17'd30994,17'd29804,17'd30995,17'd30996,17'd30997,17'd30853,17'd30697,17'd30548,17'd30699,17'd30700,17'd30551,17'd30701,17'd30998,17'd30999,17'd31000,17'd31001,17'd29804,17'd31002,17'd31003,17'd31004,17'd31005,17'd31006,17'd31007,17'd31008,17'd31009,17'd31010,17'd31011,17'd31012,17'd31013,17'd31014,17'd31015,17'd31016,17'd31017,17'd31018,17'd31019,17'd31020,17'd31021,17'd31022,17'd31023,17'd31024,17'd31025,17'd30572,17'd31026,17'd30574,17'd31027,17'd31028,17'd25553,17'd29535,17'd25566,17'd25320,17'd24416,17'd23917,17'd23732,17'd24086,17'd31029,17'd23740,17'd22506,17'd21847,17'd31030,17'd21846,17'd31031,17'd30582,17'd31032,17'd31033,17'd24249,17'd31033,17'd23732,17'd29685,17'd30431,17'd31034,17'd28598,17'd25565,17'd28978,17'd27027,17'd31035,17'd29245,17'd29379,17'd30279,17'd30279,17'd28370,17'd29247,17'd28856,17'd29106,17'd30130,17'd31036,17'd30736,17'd30736,17'd31037,17'd30739,17'd31038,17'd31039,17'd31040,17'd30887,17'd30888,17'd31041,17'd29545,17'd30287,17'd27036,17'd31042,17'd31043,17'd31044,17'd28271,17'd31045,17'd31046,17'd31047,17'd31048,17'd23916,17'd30447,17'd31049,17'd31050,17'd24430,17'd31051,17'd27899,17'd25843,17'd27533,17'd28386,17'd28620,17'd28505,17'd31052,17'd29849,17'd27380,17'd30901,17'd31053,17'd31054,17'd26287,17'd31055,17'd25835,17'd31056,17'd31057,17'd31058,17'd31059,17'd31060,17'd31061,17'd29265,17'd31062,17'd31063,17'd31064,17'd31065,17'd31066,17'd31067,17'd31068,17'd31069,17'd31070,17'd31071,17'd31072,17'd31073,17'd31074,17'd31075,17'd31076,17'd31077,17'd30478,17'd31078,17'd31079,17'd31080,17'd31081,17'd31082,17'd31083,17'd31084,17'd31085,17'd31086,17'd31087,17'd22393,17'd24142,17'd23109,17'd11158,17'd23975,17'd31088,17'd5759,17'd24799,17'd5760,17'd5481,17'd5158,17'd5332,17'd6707,17'd9090,17'd10777,17'd11576,17'd27932,17'd10897,17'd10897,17'd27932,17'd29593,17'd28183,17'd30933,17'd28183,17'd30179,17'd25627,17'd31089,17'd30637,17'd5334,17'd26949,17'd6220,17'd8780,17'd27932,17'd28305,17'd11181,17'd11577,17'd14049,17'd11853,17'd11316,17'd11316,17'd10515,17'd27815,17'd10516,17'd10517,17'd7179,17'd6711,17'd7331,17'd31090,17'd31091,17'd31092,17'd20855,17'd31093,17'd4548,17'd31094,17'd31095,17'd31096,17'd31097,17'd31098,17'd30805,17'd31099,17'd240,17'd31100,17'd4084,17'd2575,17'd7682,17'd3223,17'd28429,17'd30649,17'd29170,17'd31101,17'd31101,17'd31101,17'd31101,17'd31101,17'd29170,17'd29170,17'd28792,17'd30807,17'd27711,17'd31102,17'd30190,17'd29893,17'd30042,17'd29613,17'd24668,17'd24499,17'd24667,17'd14859,17'd18145,17'd18272,17'd1392,17'd13178,17'd3236,17'd23815,17'd3415,17'd404,17'd589,17'd615,17'd31103,17'd31104
},
'{
17'd31105,17'd7883,17'd6422,17'd5053,17'd4735,17'd4426,17'd4891,17'd4892,17'd3427,17'd14070,17'd1831,17'd4247,17'd2595,17'd2594,17'd1688,17'd3250,17'd2596,17'd2257,17'd22965,17'd22965,17'd1416,17'd1416,17'd653,17'd653,17'd27444,17'd7060,17'd7385,17'd7555,17'd7388,17'd7388,17'd6600,17'd6904,17'd27592,17'd6280,17'd5811,17'd26974,17'd5525,17'd6115,17'd26014,17'd30198,17'd4261,17'd30811,17'd30812,17'd24969,17'd31106,17'd14875,17'd29760,17'd21796,17'd30951,17'd31107,17'd31108,17'd17193,17'd14997,17'd31109,17'd31110,17'd31111,17'd19131,17'd17320,17'd14347,17'd14767,17'd14893,17'd14892,17'd17208,17'd16987,17'd17448,17'd16519,17'd17319,17'd19383,17'd19511,17'd19006,17'd30058,17'd17940,17'd15383,17'd19890,17'd15383,17'd14764,17'd13969,17'd12532,17'd17204,17'd16766,17'd15898,17'd16412,17'd14348,17'd31112,17'd31113,17'd12816,17'd20435,17'd9705,17'd18666,17'd12822,17'd9445,17'd9584,17'd10292,17'd10292,17'd18897,17'd30660,17'd30959,17'd31114,17'd29457,17'd9022,17'd31115,17'd8082,17'd28440,17'd28329,17'd31116,17'd31117,17'd31118,17'd31119,17'd31120,17'd31121,17'd28564,17'd31122,17'd31123,17'd31124,17'd16313,17'd11806,17'd13762,17'd10990,17'd11132,17'd29199,17'd31125,17'd9348,17'd30969,17'd8571,17'd8575,17'd17481,17'd17126,17'd31126,17'd8567,17'd26626,17'd11277,17'd11400,17'd11398,17'd16326,17'd18198,17'd24207,17'd27858,17'd28345,17'd30971,17'd29924,17'd30831,17'd29329,17'd30972,17'd30834,17'd31127,17'd31128,17'd31129,17'd28345,17'd18200,17'd19408,17'd18917,17'd16204,17'd11806,17'd11806,17'd11961,17'd11667,17'd11399,17'd26152,17'd10992,17'd9479,17'd19279,17'd14928,17'd14518,17'd10605,17'd14931,17'd11130,17'd21206,17'd11399,17'd11399,17'd11399,17'd12720,17'd15432,17'd31130,17'd15943,17'd16549,17'd19033,17'd31131,17'd17481,17'd15941,17'd17965,17'd31132,17'd31133,17'd28467,17'd31134,17'd31135,17'd31136,17'd29337,17'd29780,17'd29785,17'd30073,17'd29926,17'd28234,17'd14130,17'd14671,17'd22816,17'd11275,17'd31137,17'd14262,17'd30981,17'd15686,17'd30983,17'd31138,17'd30839,17'd30233,17'd31139,17'd30087,17'd31140,17'd31141,17'd31142,17'd31143,17'd30988,17'd31144,17'd31145,17'd24990,17'd31146,17'd31147,17'd29349,17'd31148,17'd31149,17'd30693,17'd31150,17'd30996,17'd31151,17'd31152,17'd31153,17'd31154,17'd31155,17'd31156,17'd30702,17'd31157,17'd31158,17'd31159,17'd31160,17'd31161,17'd31162,17'd31163,17'd31164,17'd31165,17'd31166,17'd31167,17'd31168,17'd31169,17'd31170,17'd31171,17'd31172,17'd31173,17'd31174,17'd31175,17'd31176,17'd31177,17'd31178,17'd31179,17'd31180,17'd31181,17'd31182,17'd31183,17'd31184,17'd31185,17'd31186,17'd31187,17'd30572,17'd31188,17'd30574,17'd31189,17'd30577,17'd25696,17'd28978,17'd28723,17'd25178,17'd24742,17'd24090,17'd30275,17'd23733,17'd31190,17'd31191,17'd30426,17'd23222,17'd31030,17'd31192,17'd31193,17'd31194,17'd31195,17'd23733,17'd24087,17'd24086,17'd23733,17'd29531,17'd23731,17'd29103,17'd27638,17'd25708,17'd28978,17'd30586,17'd31035,17'd29245,17'd27642,17'd27885,17'd27885,17'd28370,17'd29247,17'd28856,17'd31196,17'd29978,17'd31036,17'd30736,17'd30280,17'd31037,17'd30739,17'd31038,17'd31197,17'd31198,17'd31199,17'd31200,17'd26909,17'd29988,17'd30288,17'd31201,17'd27034,17'd28503,17'd31202,17'd28739,17'd28613,17'd31203,17'd31204,17'd31205,17'd23917,17'd29116,17'd31206,17'd31207,17'd28731,17'd24753,17'd28739,17'd25961,17'd27533,17'd31208,17'd28620,17'd28505,17'd31209,17'd28389,17'd26791,17'd30443,17'd31053,17'd31210,17'd31211,17'd31212,17'd31213,17'd31214,17'd31215,17'd31216,17'd31217,17'd23055,17'd25857,17'd31218,17'd31219,17'd31220,17'd31221,17'd31222,17'd31223,17'd31224,17'd31225,17'd31226,17'd31227,17'd31228,17'd31229,17'd31230,17'd31231,17'd31232,17'd31233,17'd31234,17'd31235,17'd31236,17'd31079,17'd31237,17'd31238,17'd31239,17'd31240,17'd31241,17'd31242,17'd31086,17'd31087,17'd22393,17'd23106,17'd23108,17'd24794,17'd6545,17'd5479,17'd5758,17'd5759,17'd26451,17'd5482,17'd5158,17'd5332,17'd6553,17'd9090,17'd10777,17'd10641,17'd27932,17'd10897,17'd10897,17'd10897,17'd29593,17'd28183,17'd31243,17'd28057,17'd12160,17'd6220,17'd31244,17'd31245,17'd5335,17'd5762,17'd6220,17'd27696,17'd28306,17'd28305,17'd11181,17'd11709,17'd14049,17'd11853,17'd11316,17'd11037,17'd10515,17'd27815,17'd10516,17'd10517,17'd8155,17'd7502,17'd6712,17'd7504,17'd12627,17'd30033,17'd20855,17'd13053,17'd31246,17'd24318,17'd27312,17'd31247,17'd31248,17'd31098,17'd27579,17'd31249,17'd241,17'd31250,17'd1823,17'd24323,17'd8317,17'd3392,17'd28315,17'd29039,17'd31251,17'd31101,17'd31101,17'd31101,17'd31101,17'd31101,17'd27708,17'd27708,17'd28792,17'd27711,17'd27711,17'd31102,17'd30650,17'd29893,17'd30190,17'd30042,17'd26967,17'd26465,17'd31252,17'd31253,17'd14061,17'd948,17'd3086,17'd1677,17'd12915,17'd31254,17'd3586,17'd610,17'd15741,17'd615,17'd16388,17'd31255
},
'{
17'd31256,17'd7046,17'd6422,17'd5053,17'd4735,17'd4426,17'd4891,17'd4892,17'd3427,17'd3252,17'd2594,17'd2595,17'd2595,17'd2594,17'd1688,17'd1688,17'd1414,17'd2257,17'd2257,17'd2257,17'd468,17'd468,17'd653,17'd653,17'd7060,17'd7061,17'd7388,17'd7388,17'd7388,17'd7388,17'd6600,17'd6904,17'd6279,17'd12337,17'd5661,17'd31257,17'd31258,17'd5665,17'd26014,17'd30198,17'd31259,17'd31260,17'd3758,17'd24969,17'd30050,17'd15368,17'd31261,17'd31262,17'd28435,17'd20282,17'd31263,17'd31264,17'd15253,17'd31265,17'd31266,17'd31267,17'd31268,17'd15902,17'd16168,17'd14626,17'd14893,17'd14892,17'd17811,17'd16987,17'd17445,17'd17319,17'd18656,17'd19383,17'd18655,17'd20886,17'd30058,17'd13211,17'd19890,17'd19890,17'd14621,17'd14764,17'd12361,17'd12532,17'd17941,17'd16410,17'd31269,17'd14896,17'd31270,17'd31271,17'd31272,17'd12816,17'd10120,17'd9989,17'd10569,17'd9444,17'd9584,17'd9585,17'd9585,17'd9585,17'd10292,17'd18897,17'd15537,17'd7429,17'd9021,17'd31273,17'd31115,17'd8082,17'd29184,17'd31274,17'd31275,17'd31276,17'd31277,17'd31278,17'd31279,17'd31280,17'd28564,17'd31281,17'd31282,17'd31283,17'd31284,17'd11962,17'd14262,17'd10990,17'd11132,17'd25530,17'd24211,17'd12118,17'd30969,17'd12425,17'd24711,17'd9887,17'd8099,17'd8246,17'd8722,17'd25525,17'd14928,17'd19282,17'd11808,17'd18443,17'd21671,17'd27123,17'd28345,17'd28686,17'd31285,17'd29067,17'd31286,17'd30072,17'd30973,17'd31287,17'd31288,17'd31289,17'd31290,17'd26873,17'd25671,17'd17722,17'd18917,17'd12996,17'd11961,17'd11806,17'd11667,17'd14673,17'd11400,17'd10169,17'd9480,17'd11809,17'd11277,17'd11134,17'd10476,17'd14810,17'd10990,17'd14263,17'd19282,17'd14134,17'd11399,17'd13138,17'd13137,17'd12862,17'd10477,17'd15431,17'd15944,17'd9482,17'd12725,17'd9886,17'd31291,17'd31292,17'd31293,17'd30077,17'd29337,17'd29483,17'd31294,17'd29483,17'd31295,17'd31295,17'd29930,17'd31296,17'd28823,17'd23855,17'd19158,17'd10854,17'd14263,17'd20451,17'd31297,17'd11957,17'd12576,17'd13760,17'd29340,17'd30232,17'd30233,17'd30234,17'd30235,17'd31298,17'd31141,17'd30986,17'd31299,17'd31300,17'd30384,17'd31145,17'd10984,17'd31301,17'd31302,17'd29348,17'd29800,17'd31001,17'd30391,17'd31303,17'd31304,17'd31305,17'd31306,17'd31307,17'd30699,17'd31308,17'd31309,17'd31158,17'd30703,17'd30858,17'd31309,17'd31310,17'd31311,17'd31312,17'd31313,17'd31314,17'd31315,17'd31316,17'd31317,17'd31318,17'd31319,17'd31320,17'd31321,17'd31322,17'd31323,17'd31324,17'd31325,17'd31326,17'd31327,17'd31328,17'd31329,17'd31330,17'd31331,17'd31332,17'd31333,17'd31334,17'd31335,17'd31336,17'd31337,17'd31338,17'd31339,17'd31026,17'd30575,17'd31340,17'd31028,17'd25696,17'd28724,17'd28723,17'd25178,17'd24742,17'd29100,17'd23564,17'd23918,17'd31341,17'd31342,17'd31343,17'd31344,17'd31345,17'd31346,17'd31347,17'd31348,17'd31349,17'd31350,17'd31032,17'd23733,17'd23733,17'd29531,17'd30275,17'd29103,17'd27638,17'd27766,17'd31351,17'd27146,17'd31035,17'd31352,17'd31353,17'd31354,17'd27885,17'd28133,17'd29247,17'd29105,17'd31196,17'd29978,17'd31036,17'd30736,17'd30736,17'd31037,17'd30739,17'd30738,17'd31197,17'd31355,17'd31356,17'd29990,17'd26909,17'd29839,17'd30288,17'd31201,17'd27893,17'd28732,17'd31202,17'd25328,17'd31357,17'd31358,17'd29689,17'd31359,17'd24085,17'd31360,17'd31361,17'd27771,17'd31362,17'd30892,17'd28739,17'd25961,17'd27533,17'd30296,17'd28024,17'd27785,17'd31363,17'd28028,17'd26792,17'd27270,17'd30758,17'd30604,17'd31364,17'd31365,17'd31366,17'd31367,17'd31368,17'd30760,17'd31369,17'd31370,17'd22525,17'd22183,17'd31371,17'd31372,17'd31373,17'd31374,17'd31375,17'd31376,17'd31377,17'd31378,17'd31379,17'd31380,17'd31381,17'd31382,17'd31383,17'd31384,17'd31385,17'd31386,17'd31387,17'd31388,17'd31389,17'd31390,17'd31391,17'd31392,17'd31393,17'd31394,17'd31395,17'd31396,17'd31397,17'd31398,17'd23625,17'd31399,17'd10881,17'd6381,17'd5326,17'd5610,17'd5759,17'd26451,17'd5482,17'd5158,17'd5331,17'd6218,17'd8154,17'd10513,17'd10777,17'd27932,17'd27932,17'd10897,17'd10897,17'd27933,17'd27933,17'd27933,17'd27934,17'd28183,17'd10514,17'd31400,17'd31401,17'd5160,17'd5614,17'd7499,17'd27696,17'd28306,17'd28305,17'd11181,17'd14049,17'd14049,17'd11853,17'd11037,17'd31402,17'd27815,17'd27815,17'd10516,17'd10517,17'd6854,17'd6710,17'd8156,17'd7182,17'd31403,17'd25882,17'd21008,17'd22427,17'd31246,17'd25636,17'd31404,17'd31405,17'd31406,17'd31407,17'd30498,17'd18386,17'd240,17'd31408,17'd1396,17'd2740,17'd4401,17'd3074,17'd28315,17'd29441,17'd31101,17'd31101,17'd31101,17'd31101,17'd31101,17'd31101,17'd31409,17'd31409,17'd27822,17'd31410,17'd31410,17'd31411,17'd30650,17'd30042,17'd30190,17'd24324,17'd24955,17'd2396,17'd14979,17'd31253,17'd14061,17'd13809,17'd1677,17'd2762,17'd2921,17'd2577,17'd9790,17'd594,17'd614,17'd615,17'd31412,17'd31413
},
'{
17'd9262,17'd7046,17'd6422,17'd5053,17'd4735,17'd4426,17'd3902,17'd4892,17'd2934,17'd3252,17'd2594,17'd2595,17'd2595,17'd2594,17'd1831,17'd3250,17'd2596,17'd2257,17'd2257,17'd2257,17'd1692,17'd468,17'd653,17'd653,17'd7060,17'd7061,17'd7388,17'd7388,17'd7388,17'd7388,17'd6600,17'd6904,17'd6279,17'd12337,17'd5660,17'd31414,17'd31258,17'd31415,17'd26014,17'd30048,17'd31259,17'd31260,17'd3758,17'd24832,17'd23826,17'd15368,17'd31416,17'd29900,17'd30053,17'd4754,17'd31417,17'd15252,17'd15504,17'd31418,17'd31419,17'd31420,17'd18776,17'd14346,17'd14626,17'd14626,17'd15384,17'd14892,17'd17811,17'd16987,17'd17445,17'd17319,17'd18656,17'd19383,17'd18774,17'd20424,17'd24347,17'd13211,17'd13599,17'd13210,17'd14621,17'd12361,17'd12531,17'd17204,17'd16766,17'd15765,17'd14896,17'd31421,17'd31422,17'd31423,17'd31424,17'd21489,17'd9845,17'd18179,17'd9992,17'd9850,17'd9584,17'd9585,17'd9585,17'd9585,17'd10292,17'd31425,17'd15537,17'd7429,17'd8858,17'd31426,17'd31427,17'd31428,17'd31429,17'd31430,17'd31431,17'd31432,17'd31433,17'd31434,17'd31435,17'd31436,17'd30366,17'd10586,17'd31437,17'd11273,17'd31284,17'd11963,17'd10989,17'd10739,17'd11132,17'd26759,17'd24040,17'd8410,17'd31438,17'd8570,17'd24545,17'd24213,17'd17126,17'd12723,17'd8875,17'd15569,17'd11135,17'd11132,17'd11397,17'd16325,17'd25671,17'd28227,17'd29067,17'd31439,17'd31440,17'd30072,17'd30072,17'd30676,17'd31441,17'd31442,17'd31288,17'd30677,17'd28462,17'd31443,17'd24362,17'd21361,17'd18917,17'd11806,17'd13363,17'd12861,17'd16068,17'd10476,17'd11671,17'd11136,17'd9742,17'd9741,17'd9883,17'd10326,17'd10739,17'd10990,17'd10854,17'd11669,17'd11400,17'd15176,17'd11524,17'd12720,17'd16064,17'd14931,17'd17720,17'd16065,17'd8886,17'd12587,17'd9887,17'd31444,17'd31445,17'd31446,17'd26872,17'd28466,17'd30679,17'd31447,17'd30976,17'd30079,17'd31448,17'd30073,17'd29926,17'd30376,17'd27736,17'd17722,17'd11130,17'd13886,17'd10474,17'd29203,17'd11962,17'd12258,17'd13518,17'd30378,17'd30232,17'd30232,17'd30840,17'd31449,17'd31450,17'd31451,17'd31452,17'd30536,17'd31144,17'd31453,17'd31454,17'd31455,17'd31456,17'd29809,17'd31457,17'd31458,17'd30249,17'd31459,17'd31460,17'd31311,17'd30854,17'd31461,17'd31462,17'd30549,17'd31309,17'd30998,17'd31158,17'd30858,17'd31463,17'd30549,17'd31464,17'd31465,17'd31466,17'd31467,17'd31468,17'd31315,17'd31469,17'd31470,17'd31471,17'd31472,17'd31473,17'd31474,17'd31475,17'd31476,17'd31477,17'd31478,17'd31479,17'd31480,17'd31327,17'd31481,17'd31482,17'd31483,17'd31484,17'd31485,17'd31486,17'd31487,17'd31488,17'd31489,17'd31490,17'd31491,17'd30271,17'd30573,17'd31492,17'd31493,17'd31494,17'd27369,17'd28978,17'd28723,17'd25320,17'd28851,17'd24415,17'd23732,17'd23920,17'd31341,17'd31495,17'd31496,17'd31497,17'd23041,17'd23041,17'd31498,17'd31499,17'd31500,17'd31501,17'd24592,17'd30127,17'd31502,17'd29975,17'd29689,17'd25320,17'd27765,17'd28720,17'd28252,17'd27372,17'd31035,17'd31352,17'd31353,17'd31503,17'd27885,17'd28133,17'd29247,17'd29105,17'd31504,17'd29979,17'd30736,17'd31505,17'd31506,17'd31037,17'd30885,17'd30738,17'd30588,17'd31507,17'd31356,17'd29990,17'd27034,17'd27379,17'd30890,17'd31508,17'd30899,17'd28732,17'd31509,17'd31510,17'd28261,17'd31511,17'd29972,17'd26527,17'd26397,17'd31512,17'd31513,17'd31514,17'd31515,17'd29546,17'd28739,17'd25961,17'd25458,17'd27661,17'd28024,17'd27785,17'd31516,17'd31517,17'd31052,17'd31518,17'd29987,17'd30758,17'd28260,17'd31519,17'd31520,17'd23912,17'd31521,17'd31522,17'd31523,17'd31524,17'd23232,17'd25974,17'd31525,17'd31526,17'd31527,17'd31528,17'd31529,17'd31530,17'd31531,17'd31532,17'd31533,17'd31534,17'd31535,17'd31536,17'd31537,17'd31538,17'd31539,17'd31540,17'd31541,17'd31542,17'd31543,17'd31543,17'd31544,17'd31545,17'd31546,17'd31547,17'd31548,17'd31396,17'd31397,17'd31549,17'd31550,17'd23796,17'd23109,17'd6544,17'd5326,17'd5758,17'd5759,17'd5760,17'd5482,17'd5158,17'd5158,17'd6389,17'd8303,17'd9657,17'd10777,17'd27932,17'd27932,17'd27932,17'd10897,17'd27933,17'd29592,17'd27933,17'd28057,17'd31551,17'd28183,17'd28185,17'd31552,17'd31553,17'd6554,17'd7499,17'd27696,17'd28650,17'd27932,17'd11576,17'd11853,17'd11853,17'd30332,17'd31402,17'd11038,17'd27815,17'd27815,17'd10516,17'd10517,17'd6854,17'd7013,17'd7838,17'd7330,17'd12472,17'd31554,17'd21008,17'd12314,17'd31246,17'd31555,17'd31556,17'd31557,17'd31558,17'd31098,17'd31559,17'd22264,17'd31560,17'd31408,17'd1666,17'd1668,17'd4401,17'd31561,17'd31562,17'd29441,17'd31101,17'd31101,17'd31101,17'd31101,17'd31101,17'd31101,17'd31409,17'd31409,17'd29040,17'd31410,17'd27822,17'd31563,17'd30650,17'd30042,17'd30650,17'd30190,17'd26967,17'd26465,17'd2561,17'd1385,17'd14179,17'd13809,17'd2762,17'd2762,17'd2921,17'd2922,17'd19607,17'd610,17'd791,17'd20000,17'd31564,17'd31255
},
'{
17'd9262,17'd7046,17'd5375,17'd5053,17'd5201,17'd4426,17'd3902,17'd4892,17'd2934,17'd3252,17'd4247,17'd2595,17'd2595,17'd2594,17'd1831,17'd2422,17'd2596,17'd2597,17'd2257,17'd2257,17'd1692,17'd468,17'd653,17'd653,17'd7060,17'd7061,17'd7388,17'd7388,17'd7388,17'd7388,17'd6600,17'd6904,17'd6279,17'd12337,17'd5659,17'd31565,17'd31566,17'd31415,17'd31567,17'd30048,17'd31259,17'd31259,17'd3919,17'd24832,17'd13190,17'd13955,17'd31416,17'd2279,17'd29453,17'd31568,17'd31569,17'd26243,17'd31570,17'd31571,17'd31572,17'd31573,17'd16290,17'd14474,17'd31574,17'd15519,17'd15384,17'd14892,17'd16987,17'd15902,17'd17320,17'd17319,17'd18656,17'd18655,17'd19006,17'd30058,17'd29904,17'd13211,17'd13210,17'd13210,17'd14621,17'd14622,17'd16658,17'd19753,17'd16766,17'd17097,17'd31575,17'd31576,17'd31577,17'd31271,17'd31424,17'd12067,17'd31578,17'd14358,17'd18667,17'd9850,17'd9584,17'd9585,17'd9585,17'd9585,17'd10570,17'd31425,17'd15537,17'd7429,17'd8858,17'd31426,17'd8227,17'd31428,17'd31429,17'd31579,17'd31580,17'd31581,17'd31582,17'd31583,17'd31584,17'd31585,17'd30366,17'd29320,17'd28682,17'd24702,17'd16797,17'd19157,17'd10853,17'd10475,17'd19282,17'd16070,17'd15430,17'd9482,17'd8411,17'd31586,17'd11531,17'd14812,17'd17126,17'd11137,17'd9038,17'd9619,17'd10479,17'd21206,17'd11522,17'd15055,17'd26036,17'd28344,17'd31439,17'd30834,17'd31439,17'd31587,17'd30972,17'd31588,17'd31589,17'd31590,17'd31591,17'd29785,17'd28943,17'd26493,17'd21505,17'd21361,17'd17722,17'd11958,17'd12857,17'd11963,17'd10604,17'd10164,17'd9885,17'd10025,17'd9742,17'd12116,17'd12863,17'd11132,17'd10854,17'd11131,17'd11669,17'd11669,17'd15176,17'd14134,17'd17236,17'd12862,17'd11520,17'd20910,17'd10479,17'd13887,17'd10177,17'd14812,17'd14812,17'd31592,17'd31593,17'd31594,17'd29336,17'd29485,17'd31595,17'd31596,17'd29201,17'd30073,17'd31597,17'd30371,17'd29642,17'd31598,17'd22819,17'd18444,17'd19282,17'd17720,17'd27743,17'd20910,17'd28695,17'd12576,17'd29208,17'd31599,17'd30683,17'd31600,17'd31601,17'd31602,17'd31603,17'd31604,17'd31142,17'd31299,17'd31605,17'd31606,17'd31607,17'd31608,17'd31609,17'd29662,17'd31610,17'd31611,17'd31612,17'd31613,17'd31614,17'd31615,17'd31616,17'd31617,17'd31159,17'd31618,17'd31619,17'd30999,17'd31620,17'd31621,17'd31310,17'd31622,17'd31623,17'd31624,17'd31625,17'd31626,17'd31627,17'd31628,17'd31629,17'd31630,17'd31631,17'd31632,17'd31633,17'd31634,17'd31635,17'd31636,17'd31637,17'd31638,17'd31639,17'd31640,17'd31327,17'd31641,17'd31642,17'd31643,17'd31644,17'd31645,17'd31646,17'd31647,17'd31648,17'd31488,17'd31649,17'd31650,17'd31651,17'd31652,17'd31653,17'd31654,17'd31494,17'd27369,17'd28978,17'd28720,17'd25178,17'd24416,17'd24415,17'd30275,17'd31029,17'd31655,17'd31656,17'd31657,17'd31658,17'd31659,17'd31660,17'd31661,17'd31662,17'd23391,17'd31663,17'd31664,17'd31502,17'd29376,17'd29975,17'd23385,17'd29976,17'd27765,17'd28594,17'd25707,17'd27146,17'd30586,17'd30735,17'd31353,17'd31503,17'd31354,17'd28255,17'd28133,17'd28981,17'd28856,17'd29831,17'd30736,17'd31505,17'd31506,17'd31037,17'd30885,17'd30738,17'd30588,17'd31507,17'd31665,17'd30747,17'd27034,17'd27379,17'd30289,17'd31666,17'd31667,17'd25849,17'd31509,17'd31668,17'd31669,17'd31670,17'd31671,17'd31672,17'd31673,17'd30446,17'd26065,17'd31674,17'd31675,17'd31676,17'd24909,17'd27043,17'd25342,17'd27661,17'd27391,17'd28620,17'd31677,17'd27785,17'd31678,17'd29557,17'd31679,17'd31680,17'd29263,17'd31681,17'd31682,17'd25175,17'd25026,17'd27512,17'd31683,17'd31684,17'd31685,17'd31686,17'd31687,17'd31688,17'd31689,17'd31690,17'd31691,17'd31692,17'd31693,17'd31694,17'd31695,17'd31696,17'd31697,17'd31698,17'd31699,17'd31700,17'd31701,17'd31702,17'd31703,17'd31704,17'd31705,17'd31706,17'd31707,17'd31708,17'd31709,17'd31710,17'd31711,17'd31712,17'd31397,17'd31549,17'd31713,17'd31714,17'd9637,17'd24649,17'd5480,17'd5758,17'd24799,17'd5482,17'd5760,17'd5332,17'd5612,17'd26218,17'd6218,17'd9090,17'd10513,17'd10897,17'd11181,17'd27932,17'd10897,17'd27933,17'd27933,17'd10515,17'd27933,17'd31715,17'd31551,17'd6221,17'd31716,17'd31400,17'd31717,17'd7499,17'd27696,17'd10897,17'd27932,17'd10641,17'd11853,17'd12160,17'd30332,17'd31402,17'd11038,17'd29592,17'd29592,17'd29592,17'd31718,17'd8002,17'd7179,17'd6394,17'd10898,17'd8158,17'd31719,17'd13052,17'd12314,17'd31720,17'd31721,17'd31722,17'd31723,17'd31724,17'd31725,17'd31559,17'd29749,17'd31726,17'd31727,17'd1112,17'd192,17'd3712,17'd31728,17'd28066,17'd31409,17'd31729,17'd31729,17'd31729,17'd31101,17'd31101,17'd31101,17'd31409,17'd31409,17'd29039,17'd27822,17'd27822,17'd31563,17'd27320,17'd29041,17'd30650,17'd2563,17'd24955,17'd2395,17'd14978,17'd1385,17'd14179,17'd13573,17'd2762,17'd780,17'd8165,17'd26595,17'd10073,17'd404,17'd433,17'd19864,17'd586,17'd31730
},
'{
17'd9262,17'd7046,17'd6422,17'd5053,17'd5200,17'd4087,17'd3902,17'd4892,17'd3101,17'd3252,17'd4247,17'd4247,17'd4247,17'd2594,17'd1831,17'd2422,17'd2596,17'd2596,17'd2257,17'd2257,17'd1692,17'd468,17'd653,17'd653,17'd7060,17'd7061,17'd7388,17'd7388,17'd7388,17'd7388,17'd6600,17'd6904,17'd6279,17'd12786,17'd26847,17'd26471,17'd26236,17'd31731,17'd31567,17'd25903,17'd30654,17'd31260,17'd31732,17'd31733,17'd31734,17'd13955,17'd31735,17'd30202,17'd31736,17'd31737,17'd31569,17'd31738,17'd31739,17'd31740,17'd31741,17'd17575,17'd14346,17'd15384,17'd31742,17'd31743,17'd15641,17'd14892,17'd16987,17'd15902,17'd16519,17'd17319,17'd18656,17'd18774,17'd18884,17'd30058,17'd24347,17'd13211,17'd14621,17'd15383,17'd14764,17'd14622,17'd12681,17'd18655,17'd20426,17'd16883,17'd31744,17'd31745,17'd31577,17'd31746,17'd31747,17'd31748,17'd19020,17'd18178,17'd14903,17'd9850,17'd9584,17'd9585,17'd9585,17'd9311,17'd10570,17'd31425,17'd15537,17'd7266,17'd8858,17'd31749,17'd31750,17'd31751,17'd31752,17'd31753,17'd31754,17'd31755,17'd31756,17'd9329,17'd31757,17'd31758,17'd29467,17'd29469,17'd10322,17'd28696,17'd16797,17'd15810,17'd20910,17'd10475,17'd19532,17'd11277,17'd9188,17'd15568,17'd31759,17'd31760,17'd11811,17'd14812,17'd9483,17'd10607,17'd10174,17'd12116,17'd11670,17'd11399,17'd14264,17'd30229,17'd26872,17'd30071,17'd31761,17'd31762,17'd31763,17'd31764,17'd31765,17'd31128,17'd31766,17'd31589,17'd31767,17'd31768,17'd28816,17'd24538,17'd21505,17'd21361,17'd17603,17'd12420,17'd12260,17'd14262,17'd10991,17'd9740,17'd9480,17'd9480,17'd18556,17'd11671,17'd10478,17'd13886,17'd10854,17'd14263,17'd24996,17'd19282,17'd14134,17'd12584,17'd12720,17'd16068,17'd10736,17'd10991,17'd22131,17'd9194,17'd10178,17'd21208,17'd31769,17'd17606,17'd31770,17'd28106,17'd31771,17'd30977,17'd31772,17'd30078,17'd30530,17'd30677,17'd31773,17'd29785,17'd28824,17'd19283,17'd12582,17'd11275,17'd10477,17'd15300,17'd27743,17'd11666,17'd12577,17'd14523,17'd31774,17'd31775,17'd31776,17'd30840,17'd31777,17'd31778,17'd31779,17'd31142,17'd31780,17'd31781,17'd31782,17'd31783,17'd31784,17'd29501,17'd29806,17'd31785,17'd31612,17'd31786,17'd31787,17'd31788,17'd31789,17'd31790,17'd30998,17'd31791,17'd31792,17'd31793,17'd30999,17'd31620,17'd31160,17'd31794,17'd30854,17'd31795,17'd31796,17'd31797,17'd31626,17'd31798,17'd31628,17'd31629,17'd31799,17'd31800,17'd31801,17'd31802,17'd31803,17'd31804,17'd31805,17'd31806,17'd31807,17'd31808,17'd31809,17'd31810,17'd31811,17'd31812,17'd31813,17'd31814,17'd31815,17'd31816,17'd31817,17'd31818,17'd31819,17'd31820,17'd31821,17'd31822,17'd31338,17'd31823,17'd31824,17'd31825,17'd31826,17'd30423,17'd31827,17'd25566,17'd25438,17'd25032,17'd23916,17'd31033,17'd31029,17'd31828,17'd22857,17'd31829,17'd31830,17'd31659,17'd31831,17'd31832,17'd31833,17'd31834,17'd31835,17'd31836,17'd24421,17'd23387,17'd29374,17'd29687,17'd25180,17'd28369,17'd27638,17'd25833,17'd27146,17'd26901,17'd30735,17'd31352,17'd31503,17'd27885,17'd28256,17'd29247,17'd28855,17'd28856,17'd29536,17'd30736,17'd31837,17'd31506,17'd31838,17'd31839,17'd31839,17'd30588,17'd31840,17'd31665,17'd31841,17'd27034,17'd27269,17'd31201,17'd31666,17'd30899,17'd25849,17'd31509,17'd31668,17'd31842,17'd31843,17'd24903,17'd29828,17'd31844,17'd24742,17'd25835,17'd31845,17'd31846,17'd31847,17'd25585,17'd27043,17'd25853,17'd27533,17'd31848,17'd28620,17'd31849,17'd31850,17'd31851,17'd31852,17'd31853,17'd31854,17'd30594,17'd31855,17'd31856,17'd23725,17'd25174,17'd31857,17'd29115,17'd31858,17'd31859,17'd23939,17'd31860,17'd31861,17'd31862,17'd31863,17'd31527,17'd31864,17'd31865,17'd31866,17'd31867,17'd31868,17'd31869,17'd31870,17'd31871,17'd31872,17'd31873,17'd31874,17'd31875,17'd31876,17'd31877,17'd31878,17'd31879,17'd31880,17'd31239,17'd31881,17'd31882,17'd31883,17'd31884,17'd31885,17'd31886,17'd23794,17'd31887,17'd5322,17'd5325,17'd5610,17'd5760,17'd5331,17'd6388,17'd6387,17'd5158,17'd5331,17'd6218,17'd8154,17'd10513,17'd10897,17'd11181,17'd27932,17'd10897,17'd27815,17'd10642,17'd10515,17'd31888,17'd31889,17'd31551,17'd25084,17'd4842,17'd31890,17'd31891,17'd7499,17'd27696,17'd27931,17'd10897,17'd27932,17'd11853,17'd12160,17'd10642,17'd11038,17'd11038,17'd29592,17'd29593,17'd29592,17'd31718,17'd8002,17'd7013,17'd7670,17'd6712,17'd7183,17'd31892,17'd29600,17'd12171,17'd31720,17'd31893,17'd31894,17'd31895,17'd31558,17'd31896,17'd31559,17'd31897,17'd210,17'd31898,17'd1112,17'd5957,17'd6888,17'd31728,17'd31899,17'd31409,17'd31729,17'd31729,17'd31729,17'd31101,17'd31101,17'd31101,17'd31409,17'd31900,17'd29039,17'd29040,17'd29040,17'd31901,17'd27320,17'd29171,17'd27583,17'd27208,17'd26967,17'd31902,17'd2561,17'd31903,17'd14179,17'd13573,17'd2762,17'd780,17'd2576,17'd4084,17'd1678,17'd1096,17'd249,17'd435,17'd219,17'd31904
},
'{
17'd7543,17'd7542,17'd7043,17'd5199,17'd5200,17'd31905,17'd4243,17'd6420,17'd3101,17'd3252,17'd1831,17'd4247,17'd2594,17'd1831,17'd1831,17'd1688,17'd1414,17'd1414,17'd1414,17'd2257,17'd468,17'd289,17'd652,17'd28,17'd7060,17'd7555,17'd7557,17'd7388,17'd7388,17'd7388,17'd6904,17'd27592,17'd5809,17'd5659,17'd26733,17'd26471,17'd31906,17'd31907,17'd31908,17'd31909,17'd4097,17'd30812,17'd3601,17'd3109,17'd31910,17'd13955,17'd31911,17'd31912,17'd31107,17'd31108,17'd17432,17'd31913,17'd31914,17'd31915,17'd31916,17'd18175,17'd14892,17'd31917,17'd31918,17'd16029,17'd14892,17'd14768,17'd15902,17'd17445,17'd18060,17'd19255,17'd18655,17'd22630,17'd17940,17'd17096,17'd17096,17'd13211,17'd13211,17'd14621,17'd18411,17'd15764,17'd19006,17'd21649,17'd31919,17'd31920,17'd31921,17'd31922,17'd31923,17'd31924,17'd31925,17'd31926,17'd31927,17'd15022,17'd31928,17'd31928,17'd18421,17'd9584,17'd18786,17'd10292,17'd18786,17'd31929,17'd15537,17'd29457,17'd31930,17'd8859,17'd31931,17'd31932,17'd8707,17'd31933,17'd31934,17'd31935,17'd31936,17'd31937,17'd29915,17'd31938,17'd28220,17'd31939,17'd27001,17'd16435,17'd11807,17'd13516,17'd10738,17'd10603,17'd10330,17'd16549,17'd12722,17'd14135,17'd8576,17'd23173,17'd19923,17'd13139,17'd9744,17'd9348,17'd9344,17'd17719,17'd11400,17'd25280,17'd28112,17'd26149,17'd27984,17'd31940,17'd31765,17'd31761,17'd31761,17'd31941,17'd30973,17'd31942,17'd31943,17'd31127,17'd29925,17'd27984,17'd26493,17'd23170,17'd21362,17'd18198,17'd12420,17'd11958,17'd13362,17'd10990,17'd11134,17'd9479,17'd9620,17'd9742,17'd17719,17'd11670,17'd10477,17'd11132,17'd11669,17'd19532,17'd10326,17'd10326,17'd21206,17'd11274,17'd11396,17'd14673,17'd17715,17'd14928,17'd24361,17'd30217,17'd17483,17'd10178,17'd31944,17'd31945,17'd31946,17'd31947,17'd30979,17'd31948,17'd31949,17'd31950,17'd30678,17'd30677,17'd30972,17'd29779,17'd30082,17'd15053,17'd20451,17'd10738,17'd31951,17'd31952,17'd14262,17'd14131,17'd12253,17'd21057,17'd31774,17'd31953,17'd30234,17'd31954,17'd31955,17'd31956,17'd31957,17'd31958,17'd31959,17'd31960,17'd31961,17'd31609,17'd31457,17'd29806,17'd31610,17'd31613,17'd31613,17'd31962,17'd31963,17'd31964,17'd30398,17'd30701,17'd31791,17'd31965,17'd31966,17'd31619,17'd31160,17'd31967,17'd31968,17'd30853,17'd31969,17'd31970,17'd31971,17'd31972,17'd31973,17'd31974,17'd31975,17'd31976,17'd31977,17'd31978,17'd31979,17'd31980,17'd31981,17'd31982,17'd31983,17'd31984,17'd31985,17'd31986,17'd31987,17'd31988,17'd31989,17'd31990,17'd31991,17'd31992,17'd31993,17'd31994,17'd31995,17'd31996,17'd31997,17'd31998,17'd31999,17'd32000,17'd32001,17'd31651,17'd32002,17'd32003,17'd32004,17'd32005,17'd32006,17'd25565,17'd25317,17'd25320,17'd32007,17'd23731,17'd29527,17'd32008,17'd22506,17'd23040,17'd32009,17'd31345,17'd32010,17'd32011,17'd32012,17'd32013,17'd32014,17'd32015,17'd29829,17'd29686,17'd29686,17'd29685,17'd28851,17'd28850,17'd27765,17'd28602,17'd27258,17'd31035,17'd32016,17'd31353,17'd27885,17'd28134,17'd32017,17'd32017,17'd27885,17'd27885,17'd32018,17'd32019,17'd31505,17'd32020,17'd32021,17'd32022,17'd32022,17'd32023,17'd32024,17'd32025,17'd30288,17'd26911,17'd27378,17'd26911,17'd27270,17'd30144,17'd28732,17'd25334,17'd32026,17'd32027,17'd32028,17'd32029,17'd32030,17'd23739,17'd24090,17'd25177,17'd27766,17'd32031,17'd32032,17'd32033,17'd26675,17'd26547,17'd32034,17'd27168,17'd31208,17'd30601,17'd31677,17'd32035,17'd28387,17'd26192,17'd32036,17'd32037,17'd32038,17'd32039,17'd31520,17'd25709,17'd28480,17'd32040,17'd32041,17'd32042,17'd32043,17'd32044,17'd32045,17'd32046,17'd32047,17'd32048,17'd32049,17'd32050,17'd32051,17'd32052,17'd32053,17'd32054,17'd32055,17'd32056,17'd32057,17'd32058,17'd32059,17'd32060,17'd32061,17'd32062,17'd32063,17'd32064,17'd31544,17'd32065,17'd32066,17'd32067,17'd32068,17'd32069,17'd7160,17'd32070,17'd32071,17'd32072,17'd7656,17'd4682,17'd5610,17'd5331,17'd26218,17'd8303,17'd6553,17'd5158,17'd5481,17'd5481,17'd6553,17'd9394,17'd8780,17'd27815,17'd10642,17'd10515,17'd28184,17'd28184,17'd29592,17'd30933,17'd31551,17'd27934,17'd30487,17'd5335,17'd31401,17'd30333,17'd32073,17'd32074,17'd9933,17'd10515,17'd10515,17'd10642,17'd10642,17'd28183,17'd28183,17'd28183,17'd10515,17'd27815,17'd10380,17'd10517,17'd7012,17'd6559,17'd11040,17'd6856,17'd7183,17'd31403,17'd12311,17'd32075,17'd4215,17'd32076,17'd32077,17'd32078,17'd32079,17'd32080,17'd32081,17'd2770,17'd17661,17'd17547,17'd1112,17'd4084,17'd6888,17'd3570,17'd32082,17'd32083,17'd31101,17'd27949,17'd27949,17'd27949,17'd31101,17'd31101,17'd31101,17'd31101,17'd29441,17'd29039,17'd27822,17'd31410,17'd27320,17'd27320,17'd27208,17'd27208,17'd27095,17'd27095,17'd2561,17'd31903,17'd24498,17'd5941,17'd780,17'd951,17'd2576,17'd26595,17'd409,17'd32084,17'd280,17'd19864,17'd31412,17'd32085
},
'{
17'd7543,17'd7542,17'd7044,17'd32086,17'd5200,17'd31905,17'd4243,17'd6420,17'd3101,17'd3252,17'd1688,17'd1688,17'd1831,17'd1831,17'd1831,17'd1831,17'd1414,17'd1414,17'd2257,17'd2257,17'd468,17'd289,17'd652,17'd28,17'd7060,17'd7555,17'd7557,17'd7388,17'd7388,17'd7388,17'd6904,17'd27592,17'd5809,17'd5383,17'd32087,17'd31906,17'd26013,17'd32088,17'd32089,17'd25792,17'd30348,17'd30812,17'd3440,17'd32090,17'd2443,17'd32091,17'd32092,17'd32093,17'd4909,17'd32094,17'd26983,17'd32095,17'd32096,17'd32097,17'd31573,17'd17811,17'd15520,17'd32098,17'd32099,17'd32100,17'd32101,17'd14768,17'd15902,17'd17445,17'd18060,17'd19255,17'd32102,17'd13969,17'd13211,17'd13599,17'd13211,17'd13094,17'd14470,17'd14470,17'd15383,17'd15764,17'd19382,17'd21037,17'd32103,17'd32104,17'd32105,17'd32106,17'd32107,17'd32108,17'd32109,17'd32110,17'd15655,17'd32111,17'd32112,17'd32113,17'd9584,17'd9584,17'd10292,17'd18786,17'd11239,17'd10818,17'd7428,17'd29457,17'd9022,17'd32114,17'd29183,17'd31932,17'd32115,17'd32116,17'd32117,17'd32118,17'd32119,17'd32120,17'd30826,17'd10718,17'd10835,17'd28225,17'd11273,17'd11520,17'd11807,17'd13645,17'd24708,17'd10740,17'd11134,17'd15569,17'd10607,17'd8418,17'd32121,17'd23343,17'd8249,17'd13139,17'd11404,17'd9041,17'd10742,17'd16796,17'd19282,17'd13367,17'd24539,17'd26493,17'd28344,17'd32122,17'd31765,17'd31761,17'd31762,17'd31127,17'd31441,17'd31942,17'd31942,17'd30973,17'd29924,17'd26757,17'd24538,17'd21505,17'd17722,17'd13883,17'd11958,17'd12858,17'd14262,17'd11132,17'd12116,17'd9480,17'd16328,17'd17965,17'd9883,17'd10326,17'd14518,17'd11133,17'd19532,17'd19532,17'd10164,17'd10326,17'd10854,17'd11274,17'd11964,17'd16068,17'd11528,17'd32123,17'd9195,17'd32124,17'd8419,17'd32125,17'd32126,17'd32127,17'd32128,17'd29926,17'd32129,17'd32130,17'd32131,17'd32132,17'd30678,17'd30073,17'd32133,17'd32134,17'd27861,17'd13762,17'd24708,17'd32135,17'd32136,17'd32137,17'd12111,17'd12109,17'd13515,17'd14525,17'd32138,17'd31138,17'd31140,17'd32139,17'd32140,17'd32141,17'd32142,17'd31605,17'd30091,17'd28939,17'd29809,17'd29216,17'd30850,17'd30103,17'd31962,17'd31962,17'd32143,17'd32144,17'd32145,17'd30701,17'd32146,17'd31791,17'd31158,17'd31619,17'd31619,17'd32147,17'd32148,17'd32149,17'd31312,17'd32150,17'd32151,17'd32152,17'd32153,17'd32154,17'd32155,17'd32156,17'd32157,17'd32158,17'd32159,17'd32160,17'd32161,17'd32162,17'd32163,17'd32164,17'd32165,17'd32166,17'd32167,17'd32168,17'd32169,17'd32170,17'd32171,17'd32172,17'd32173,17'd32174,17'd32175,17'd32176,17'd31994,17'd32177,17'd32178,17'd32179,17'd32180,17'd32181,17'd32001,17'd32182,17'd32183,17'd31824,17'd32184,17'd32185,17'd28978,17'd26174,17'd28130,17'd25438,17'd25031,17'd24415,17'd32186,17'd30128,17'd22506,17'd22163,17'd32009,17'd31497,17'd32010,17'd32187,17'd32188,17'd31344,17'd32189,17'd32190,17'd23569,17'd30128,17'd32191,17'd30278,17'd24742,17'd29103,17'd27882,17'd27513,17'd28725,17'd28486,17'd31035,17'd31352,17'd30279,17'd32192,17'd32193,17'd32017,17'd31354,17'd27885,17'd29248,17'd30885,17'd31505,17'd32020,17'd32021,17'd32194,17'd32022,17'd32195,17'd32196,17'd32197,17'd30889,17'd27378,17'd32198,17'd27893,17'd27270,17'd30891,17'd32199,17'd25042,17'd32026,17'd32027,17'd32200,17'd32201,17'd32202,17'd30882,17'd29100,17'd25177,17'd24584,17'd32203,17'd30138,17'd32204,17'd32205,17'd32206,17'd26920,17'd27168,17'd31208,17'd30451,17'd31677,17'd31516,17'd32207,17'd27162,17'd25849,17'd32208,17'd29711,17'd32209,17'd32210,17'd25709,17'd25437,17'd30139,17'd32211,17'd32212,17'd32213,17'd32214,17'd25958,17'd32215,17'd32216,17'd32217,17'd32218,17'd32219,17'd32220,17'd32221,17'd32222,17'd32223,17'd32224,17'd32225,17'd32226,17'd32227,17'd32228,17'd32229,17'd32230,17'd32231,17'd32232,17'd9760,17'd32233,17'd32234,17'd32235,17'd32236,17'd32237,17'd32238,17'd32239,17'd32240,17'd32241,17'd12601,17'd32242,17'd5756,17'd5609,17'd5159,17'd32243,17'd8933,17'd8303,17'd5331,17'd5481,17'd5481,17'd6387,17'd9090,17'd8780,17'd27815,17'd10642,17'd27815,17'd28184,17'd28184,17'd29592,17'd30933,17'd31551,17'd28057,17'd30487,17'd27935,17'd30796,17'd30333,17'd6554,17'd32074,17'd29593,17'd29592,17'd10515,17'd11037,17'd28183,17'd28183,17'd28305,17'd28306,17'd27815,17'd9933,17'd10380,17'd10517,17'd6854,17'd7836,17'd7501,17'd6561,17'd7016,17'd12472,17'd31892,17'd21006,17'd32244,17'd32245,17'd32246,17'd32247,17'd32248,17'd32249,17'd25894,17'd2111,17'd1538,17'd32250,17'd425,17'd4084,17'd6886,17'd3570,17'd32082,17'd28544,17'd27949,17'd27949,17'd28066,17'd27949,17'd31729,17'd31101,17'd31101,17'd31729,17'd29441,17'd29039,17'd27822,17'd31410,17'd27320,17'd27320,17'd27208,17'd27208,17'd32251,17'd31902,17'd28546,17'd27709,17'd2741,17'd27094,17'd1383,17'd951,17'd24323,17'd4084,17'd1240,17'd610,17'd250,17'd19864,17'd31412,17'd32252
},
'{
17'd7543,17'd7366,17'd5643,17'd5199,17'd5200,17'd31905,17'd4243,17'd15746,17'd3252,17'd2422,17'd1688,17'd1688,17'd1831,17'd10535,17'd1831,17'd1831,17'd1414,17'd1414,17'd2257,17'd2257,17'd468,17'd289,17'd652,17'd980,17'd20570,17'd7385,17'd7388,17'd7388,17'd7388,17'd7388,17'd6904,17'd27592,17'd12786,17'd32253,17'd26471,17'd31906,17'd26013,17'd4585,17'd32089,17'd25792,17'd30348,17'd3441,17'd32254,17'd32255,17'd32256,17'd32091,17'd32092,17'd32257,17'd4909,17'd25119,17'd15252,17'd31570,17'd32258,17'd32259,17'd17575,17'd16768,17'd14893,17'd32098,17'd32260,17'd15767,17'd15008,17'd16768,17'd18776,17'd17320,17'd19255,17'd25512,17'd32261,17'd14622,17'd17809,17'd13599,17'd13211,17'd14621,17'd14622,17'd14470,17'd14470,17'd22630,17'd18774,17'd21809,17'd32262,17'd32263,17'd32264,17'd31922,17'd32265,17'd32266,17'd32267,17'd32268,17'd15655,17'd32269,17'd32270,17'd32271,17'd9445,17'd9584,17'd10292,17'd11239,17'd32272,17'd10818,17'd15274,17'd7267,17'd8081,17'd32273,17'd31428,17'd32274,17'd8553,17'd32275,17'd32276,17'd32277,17'd32278,17'd32279,17'd32280,17'd10587,17'd32281,17'd10152,17'd11394,17'd11666,17'd11807,17'd13645,17'd16555,17'd10326,17'd11671,17'd15807,17'd14675,17'd24042,17'd9196,17'd12119,17'd14384,17'd8100,17'd12264,17'd16067,17'd24037,17'd16796,17'd21206,17'd23171,17'd24992,17'd29196,17'd30673,17'd32282,17'd30676,17'd31761,17'd32283,17'd31442,17'd31441,17'd31942,17'd31441,17'd30972,17'd27984,17'd24856,17'd22819,17'd20314,17'd17722,17'd13883,17'd11962,17'd19157,17'd10739,17'd10165,17'd9885,17'd9340,17'd9620,17'd18556,17'd11134,17'd10479,17'd11528,17'd11670,17'd19532,17'd10474,17'd10326,17'd11133,17'd11524,17'd14673,17'd11964,17'd14931,17'd12116,17'd17716,17'd10177,17'd21823,17'd32284,17'd16437,17'd32285,17'd32286,17'd32287,17'd29930,17'd30681,17'd32288,17'd32289,17'd32289,17'd30678,17'd30074,17'd32290,17'd31443,17'd18443,17'd11275,17'd16555,17'd32291,17'd32292,17'd32293,17'd12412,17'd13760,17'd30379,17'd31953,17'd30838,17'd32294,17'd32295,17'd31141,17'd32296,17'd32297,17'd32298,17'd32299,17'd29670,17'd32300,17'd29667,17'd29663,17'd30103,17'd32301,17'd32302,17'd32303,17'd30252,17'd31463,17'd30858,17'd31791,17'd32304,17'd31619,17'd32305,17'd32306,17'd31967,17'd32307,17'd31311,17'd31304,17'd32308,17'd32309,17'd32310,17'd32311,17'd32312,17'd32313,17'd32314,17'd32315,17'd32316,17'd32317,17'd32318,17'd32319,17'd32320,17'd32321,17'd32322,17'd32323,17'd32324,17'd32325,17'd32326,17'd32327,17'd32328,17'd32329,17'd32330,17'd32331,17'd32332,17'd32333,17'd32334,17'd32335,17'd32336,17'd32337,17'd32338,17'd32339,17'd32340,17'd32341,17'd32342,17'd31186,17'd32183,17'd31824,17'd32184,17'd32343,17'd26903,17'd26174,17'd28600,17'd28850,17'd25179,17'd24742,17'd30431,17'd23388,17'd32344,17'd32345,17'd32346,17'd21846,17'd32010,17'd32347,17'd32348,17'd23041,17'd32349,17'd32350,17'd22328,17'd32351,17'd23215,17'd32352,17'd24090,17'd32353,17'd25438,17'd28599,17'd28725,17'd28486,17'd28486,17'd31352,17'd30279,17'd32354,17'd32017,17'd32355,17'd32356,17'd31354,17'd32355,17'd30130,17'd32357,17'd31837,17'd32021,17'd32358,17'd31839,17'd29982,17'd32196,17'd32359,17'd30889,17'd30747,17'd27378,17'd26911,17'd30290,17'd29698,17'd25586,17'd25042,17'd32360,17'd24599,17'd32361,17'd32362,17'd32202,17'd32363,17'd24902,17'd25178,17'd30606,17'd32364,17'd32365,17'd32366,17'd26301,17'd29559,17'd27660,17'd27782,17'd30296,17'd28386,17'd28620,17'd31516,17'd32367,17'd32368,17'd26074,17'd32369,17'd32370,17'd32371,17'd32372,17'd25709,17'd25437,17'd25710,17'd32373,17'd32374,17'd32375,17'd31842,17'd32376,17'd32377,17'd32378,17'd32379,17'd32380,17'd32381,17'd32382,17'd32383,17'd32384,17'd32385,17'd32386,17'd32387,17'd32388,17'd32389,17'd32390,17'd32391,17'd28528,17'd32392,17'd9365,17'd32393,17'd32394,17'd32395,17'd32396,17'd32397,17'd9499,17'd7988,17'd5910,17'd7160,17'd31397,17'd32398,17'd32399,17'd4681,17'd4687,17'd25627,17'd26708,17'd26709,17'd6218,17'd6388,17'd5482,17'd5482,17'd5332,17'd8154,17'd8780,17'd10515,17'd10515,17'd28184,17'd30487,17'd28184,17'd29592,17'd30933,17'd30933,17'd28183,17'd10514,17'd5615,17'd31245,17'd31553,17'd31717,17'd9091,17'd9933,17'd29593,17'd27815,17'd11037,17'd28183,17'd28183,17'd28305,17'd28306,17'd10897,17'd9933,17'd10380,17'd10517,17'd6854,17'd7836,17'd7501,17'd30032,17'd7182,17'd30489,17'd31892,17'd11714,17'd32400,17'd3549,17'd32401,17'd32402,17'd32403,17'd32404,17'd32405,17'd32406,17'd1111,17'd424,17'd1111,17'd4084,17'd6886,17'd3570,17'd32082,17'd29751,17'd27707,17'd28066,17'd28066,17'd28066,17'd31729,17'd31729,17'd31729,17'd31729,17'd29441,17'd29039,17'd27822,17'd31410,17'd27320,17'd27320,17'd27320,17'd27208,17'd32251,17'd31902,17'd28546,17'd25238,17'd5498,17'd5941,17'd780,17'd951,17'd24323,17'd191,17'd641,17'd404,17'd770,17'd29442,17'd32407,17'd32408
},
'{
17'd7543,17'd7366,17'd5790,17'd5199,17'd5200,17'd31905,17'd4892,17'd4245,17'd2935,17'd2422,17'd1688,17'd1688,17'd1831,17'd10535,17'd10535,17'd1831,17'd1414,17'd1414,17'd2257,17'd2257,17'd468,17'd289,17'd653,17'd980,17'd20570,17'd7385,17'd7388,17'd7388,17'd7388,17'd7556,17'd6904,17'd6279,17'd12786,17'd12787,17'd5059,17'd26013,17'd4585,17'd32409,17'd25792,17'd31259,17'd32410,17'd3603,17'd3438,17'd2620,17'd30351,17'd32091,17'd32411,17'd30816,17'd32412,17'd19745,17'd26243,17'd32413,17'd32414,17'd32415,17'd18175,17'd17811,17'd31917,17'd32416,17'd32100,17'd15767,17'd15385,17'd16768,17'd18534,17'd17320,17'd19255,17'd27461,17'd12681,17'd14621,17'd13599,17'd13599,17'd14621,17'd14621,17'd14622,17'd14470,17'd14622,17'd19382,17'd21964,17'd32417,17'd32418,17'd32419,17'd32264,17'd32420,17'd31923,17'd32421,17'd32422,17'd32423,17'd32424,17'd32425,17'd32270,17'd18421,17'd9310,17'd9445,17'd10292,17'd18786,17'd11239,17'd19521,17'd15274,17'd7267,17'd8081,17'd32426,17'd32427,17'd8228,17'd32428,17'd32429,17'd32430,17'd32431,17'd9329,17'd32432,17'd32433,17'd10719,17'd32434,17'd10320,17'd11664,17'd11667,17'd15185,17'd13645,17'd16555,17'd10164,17'd14928,17'd15944,17'd8246,17'd8417,17'd25148,17'd12588,17'd13005,17'd17126,17'd8728,17'd17123,17'd15048,17'd10329,17'd11398,17'd29488,17'd24538,17'd32435,17'd30971,17'd32436,17'd30676,17'd32437,17'd32438,17'd31442,17'd31127,17'd31127,17'd31941,17'd29330,17'd26872,17'd24030,17'd22818,17'd18198,17'd15053,17'd11806,17'd11520,17'd10852,17'd11133,17'd17719,17'd11136,17'd9340,17'd9480,17'd11277,17'd16070,17'd19642,17'd11276,17'd11134,17'd10165,17'd10474,17'd19282,17'd11132,17'd13886,17'd17236,17'd14673,17'd19282,17'd15048,17'd15297,17'd22474,17'd10178,17'd32439,17'd17479,17'd30975,17'd32440,17'd31295,17'd30371,17'd32441,17'd32442,17'd32443,17'd32444,17'd30974,17'd31290,17'd28692,17'd24992,17'd30532,17'd14132,17'd10474,17'd31952,17'd15186,17'd15809,17'd13881,17'd13759,17'd32445,17'd29933,17'd32446,17'd32447,17'd32448,17'd32449,17'd32450,17'd32451,17'd32452,17'd31283,17'd32300,17'd32453,17'd30250,17'd30249,17'd30249,17'd30249,17'd32454,17'd32455,17'd31620,17'd32456,17'd30858,17'd31966,17'd31159,17'd32147,17'd31160,17'd30248,17'd30545,17'd30694,17'd32457,17'd32458,17'd32459,17'd32460,17'd32461,17'd32462,17'd32463,17'd32464,17'd32465,17'd32466,17'd32467,17'd32468,17'd32469,17'd32470,17'd32471,17'd32472,17'd32473,17'd32474,17'd32475,17'd32476,17'd32477,17'd32478,17'd32479,17'd32480,17'd32481,17'd32482,17'd32483,17'd32484,17'd32485,17'd32486,17'd32487,17'd32488,17'd32489,17'd32490,17'd32491,17'd32492,17'd31649,17'd31650,17'd32493,17'd32494,17'd32495,17'd32496,17'd28724,17'd25707,17'd28721,17'd29101,17'd30432,17'd28851,17'd29534,17'd23387,17'd22677,17'd32497,17'd32346,17'd31658,17'd32498,17'd32499,17'd32500,17'd32501,17'd32502,17'd32503,17'd22331,17'd22328,17'd22329,17'd32504,17'd28722,17'd32353,17'd25438,17'd31055,17'd27259,17'd28486,17'd28486,17'd31353,17'd29977,17'd32192,17'd32193,17'd32505,17'd32506,17'd27885,17'd32507,17'd32508,17'd31036,17'd31837,17'd32358,17'd32358,17'd31839,17'd29982,17'd32509,17'd32510,17'd32511,17'd27036,17'd32512,17'd26911,17'd30290,17'd29837,17'd25586,17'd24910,17'd32360,17'd24599,17'd32361,17'd32201,17'd32513,17'd32514,17'd23384,17'd25030,17'd28594,17'd32364,17'd32515,17'd32516,17'd29126,17'd26676,17'd27660,17'd25853,17'd25721,17'd28026,17'd28620,17'd32517,17'd32518,17'd32519,17'd26195,17'd32520,17'd32521,17'd32522,17'd32523,17'd25177,17'd31367,17'd31367,17'd32040,17'd32524,17'd32525,17'd32526,17'd31669,17'd32527,17'd32528,17'd32529,17'd32530,17'd32531,17'd32532,17'd32533,17'd32534,17'd32535,17'd32536,17'd32537,17'd32538,17'd32539,17'd32540,17'd32541,17'd32542,17'd32543,17'd32544,17'd32545,17'd32546,17'd32547,17'd32548,17'd32549,17'd9366,17'd6065,17'd32550,17'd32239,17'd31884,17'd32551,17'd10358,17'd5755,17'd32552,17'd25627,17'd26708,17'd26709,17'd6389,17'd6553,17'd5332,17'd5331,17'd6389,17'd8303,17'd8780,17'd10515,17'd10515,17'd27815,17'd28184,17'd28184,17'd29592,17'd31243,17'd31243,17'd27933,17'd10514,17'd6391,17'd31553,17'd32553,17'd31891,17'd7499,17'd9933,17'd29593,17'd27815,17'd28057,17'd28183,17'd28183,17'd28306,17'd28650,17'd27931,17'd9933,17'd10380,17'd10517,17'd10517,17'd8002,17'd6559,17'd7502,17'd7181,17'd31090,17'd12167,17'd25229,17'd32554,17'd3549,17'd32555,17'd32556,17'd32557,17'd32558,17'd32559,17'd2112,17'd603,17'd423,17'd192,17'd5957,17'd6885,17'd4559,17'd29169,17'd28544,17'd28066,17'd28066,17'd28066,17'd28066,17'd31729,17'd31101,17'd31101,17'd31729,17'd29441,17'd29039,17'd29040,17'd27822,17'd27320,17'd27320,17'd27320,17'd27320,17'd32251,17'd31902,17'd28545,17'd27580,17'd29037,17'd27094,17'd1383,17'd951,17'd24323,17'd2764,17'd1240,17'd610,17'd251,17'd20266,17'd32560,17'd176
},
'{
17'd32561,17'd7043,17'd5790,17'd5199,17'd5200,17'd31905,17'd4892,17'd14743,17'd3252,17'd2422,17'd1688,17'd1831,17'd1831,17'd10535,17'd10535,17'd1831,17'd1415,17'd1414,17'd2257,17'd2257,17'd468,17'd289,17'd652,17'd980,17'd20570,17'd7385,17'd7388,17'd7388,17'd6904,17'd9970,17'd6904,17'd27445,17'd5808,17'd32562,17'd31906,17'd26013,17'd4585,17'd32409,17'd32409,17'd31259,17'd30812,17'd3268,17'd32563,17'd2620,17'd30351,17'd32564,17'd21480,17'd4908,17'd20018,17'd18047,17'd32565,17'd32566,17'd32567,17'd32568,17'd16768,17'd14767,17'd32569,17'd32098,17'd16029,17'd15767,17'd15385,17'd16411,17'd18060,17'd19008,17'd25512,17'd30511,17'd16658,17'd13211,17'd13599,17'd32570,17'd19890,17'd15383,17'd14470,17'd14622,17'd22630,17'd19382,17'd32571,17'd31744,17'd32572,17'd32573,17'd32264,17'd32420,17'd32574,17'd32575,17'd32576,17'd32268,17'd32577,17'd32578,17'd32579,17'd18421,17'd9445,17'd11095,17'd9311,17'd9585,17'd9311,17'd19521,17'd16666,17'd7267,17'd32580,17'd32426,17'd32427,17'd32581,17'd32582,17'd32583,17'd32584,17'd32585,17'd32586,17'd32587,17'd32588,17'd32589,17'd10723,17'd10844,17'd32590,17'd11667,17'd19158,17'd13645,17'd16555,17'd17720,17'd16070,17'd10174,17'd18808,17'd8417,17'd8733,17'd9888,17'd13004,17'd17481,17'd8569,17'd16553,17'd25673,17'd10326,17'd11396,17'd24539,17'd26493,17'd32591,17'd32133,17'd32282,17'd31765,17'd32437,17'd32438,17'd32592,17'd31287,17'd30973,17'd31440,17'd28345,17'd24856,17'd22819,17'd17474,17'd12106,17'd13135,17'd11666,17'd24860,17'd10606,17'd9739,17'd9885,17'd13255,17'd13255,17'd9741,17'd14928,17'd26759,17'd26759,17'd9884,17'd11671,17'd25811,17'd10472,17'd11132,17'd10476,17'd12721,17'd10605,17'd10739,17'd10741,17'd25814,17'd32125,17'd22298,17'd32593,17'd32594,17'd32595,17'd28692,17'd32596,17'd32597,17'd32598,17'd32599,17'd32599,17'd32600,17'd32601,17'd30974,17'd32602,17'd28468,17'd21361,17'd11275,17'd10473,17'd27738,17'd18560,17'd12111,17'd13763,17'd32603,17'd32604,17'd32605,17'd32606,17'd32607,17'd32608,17'd32609,17'd32610,17'd32611,17'd32612,17'd32613,17'd32614,17'd29808,17'd32615,17'd30396,17'd32616,17'd32454,17'd32617,17'd29800,17'd32618,17'd32147,17'd32147,17'd32619,17'd32619,17'd32147,17'd32620,17'd32621,17'd32457,17'd32622,17'd32623,17'd32624,17'd32624,17'd32625,17'd32626,17'd32627,17'd32628,17'd32629,17'd32630,17'd32631,17'd32632,17'd32633,17'd32634,17'd32635,17'd32636,17'd32637,17'd32638,17'd32639,17'd32640,17'd32641,17'd32642,17'd32643,17'd32644,17'd32645,17'd32646,17'd32647,17'd32648,17'd32332,17'd32649,17'd32650,17'd32651,17'd32652,17'd32653,17'd32654,17'd32655,17'd32489,17'd31487,17'd32656,17'd31822,17'd32657,17'd32003,17'd32495,17'd32185,17'd29535,17'd31351,17'd32658,17'd25317,17'd29244,17'd24745,17'd32659,17'd23566,17'd22678,17'd32660,17'd32661,17'd23220,17'd32662,17'd32663,17'd32664,17'd21695,17'd32665,17'd32666,17'd22681,17'd22500,17'd22500,17'd32667,17'd29243,17'd32668,17'd25438,17'd32669,17'd27515,17'd27027,17'd28486,17'd31353,17'd30279,17'd32354,17'd32355,17'd32505,17'd28258,17'd27885,17'd32507,17'd29979,17'd32357,17'd32670,17'd31506,17'd32671,17'd31839,17'd29982,17'd32672,17'd32673,17'd32674,17'd27036,17'd32512,17'd32675,17'd30297,17'd28148,17'd28147,17'd27033,17'd32676,17'd32677,17'd32361,17'd32678,17'd32679,17'd32680,17'd28976,17'd24745,17'd27765,17'd32364,17'd32681,17'd32682,17'd29986,17'd32683,17'd25843,17'd25844,17'd32684,17'd27045,17'd27785,17'd32517,17'd32518,17'd29707,17'd26913,17'd31202,17'd32685,17'd32686,17'd32687,17'd27512,17'd25177,17'd25177,17'd32688,17'd32689,17'd32690,17'd32691,17'd32692,17'd28500,17'd32693,17'd32694,17'd32695,17'd32696,17'd32697,17'd32698,17'd32699,17'd32700,17'd32701,17'd32702,17'd32703,17'd32704,17'd32705,17'd32706,17'd32707,17'd32708,17'd32709,17'd32710,17'd32711,17'd9902,17'd32712,17'd32713,17'd12278,17'd32714,17'd32715,17'd7821,17'd32716,17'd32716,17'd32717,17'd5605,17'd32552,17'd5329,17'd6218,17'd26709,17'd6218,17'd6707,17'd6388,17'd5332,17'd26218,17'd26709,17'd7668,17'd10514,17'd10515,17'd27815,17'd28184,17'd8780,17'd29592,17'd29592,17'd29593,17'd10515,17'd30332,17'd25084,17'd5335,17'd32553,17'd32718,17'd9091,17'd9933,17'd27696,17'd29592,17'd28057,17'd28183,17'd31551,17'd28306,17'd32719,17'd10897,17'd9933,17'd10380,17'd10517,17'd10517,17'd8002,17'd6559,17'd6710,17'd7671,17'd7183,17'd12166,17'd27698,17'd32720,17'd3853,17'd32721,17'd32722,17'd32723,17'd27316,17'd32724,17'd8483,17'd1099,17'd422,17'd598,17'd11062,17'd6415,17'd4559,17'd29169,17'd32082,17'd27949,17'd28066,17'd28066,17'd28066,17'd31729,17'd31101,17'd31101,17'd31101,17'd27708,17'd29170,17'd29040,17'd27822,17'd27822,17'd27822,17'd27320,17'd27320,17'd31902,17'd32725,17'd28545,17'd27318,17'd5498,17'd27094,17'd1383,17'd951,17'd24323,17'd191,17'd641,17'd404,17'd280,17'd29753,17'd32726,17'd31104
},
'{
17'd32561,17'd32727,17'd5199,17'd5200,17'd32728,17'd31905,17'd4428,17'd4245,17'd2935,17'd2422,17'd1688,17'd1831,17'd10535,17'd10535,17'd10535,17'd1831,17'd1415,17'd1414,17'd2257,17'd2257,17'd468,17'd289,17'd652,17'd980,17'd20570,17'd7385,17'd7388,17'd7388,17'd6904,17'd9970,17'd6439,17'd27445,17'd32729,17'd5381,17'd4897,17'd32088,17'd32409,17'd32730,17'd32730,17'd31260,17'd30812,17'd3440,17'd32731,17'd32732,17'd32733,17'd14453,17'd27597,17'd31107,17'd32734,17'd19116,17'd32735,17'd32736,17'd32737,17'd32738,17'd16768,17'd15008,17'd32098,17'd24194,17'd15767,17'd15384,17'd32739,17'd15902,17'd18060,17'd19255,17'd27461,17'd19128,17'd16765,17'd17096,17'd13599,17'd32570,17'd19890,17'd19005,17'd29904,17'd16765,17'd19382,17'd32740,17'd32417,17'd32741,17'd32742,17'd32743,17'd32744,17'd32745,17'd32266,17'd32422,17'd32423,17'd32746,17'd32747,17'd32748,17'd18421,17'd9584,17'd9311,17'd11095,17'd11095,17'd9585,17'd9311,17'd12370,17'd8702,17'd8224,17'd32580,17'd32749,17'd7928,17'd32750,17'd32751,17'd32752,17'd32753,17'd32754,17'd32755,17'd32756,17'd32757,17'd32758,17'd9878,17'd27001,17'd11519,17'd11667,17'd16326,17'd24029,17'd16555,17'd17720,17'd15431,17'd9041,17'd12724,17'd19780,17'd11674,17'd17849,17'd23685,17'd8413,17'd8569,17'd24361,17'd16319,17'd11132,17'd14264,17'd26628,17'd32759,17'd32760,17'd32282,17'd32761,17'd30973,17'd32283,17'd32592,17'd31442,17'd31287,17'd31765,17'd29779,17'd27857,17'd24030,17'd19408,17'd17348,17'd12106,17'd12996,17'd11519,17'd10477,17'd25675,17'd10742,17'd10743,17'd13255,17'd10992,17'd9740,17'd17839,17'd16070,17'd14928,17'd17841,17'd11671,17'd10741,17'd10472,17'd11132,17'd11524,17'd12721,17'd12721,17'd11133,17'd22131,17'd9348,17'd32762,17'd9745,17'd32763,17'd32764,17'd32765,17'd29926,17'd32766,17'd32767,17'd32768,17'd32769,17'd32768,17'd32770,17'd32597,17'd31295,17'd28825,17'd23168,17'd16326,17'd10853,17'd27738,17'd25144,17'd12861,17'd13136,17'd18684,17'd32604,17'd31139,17'd32606,17'd32771,17'd32772,17'd32773,17'd32774,17'd32775,17'd32776,17'd32777,17'd32778,17'd32779,17'd32780,17'd30250,17'd32781,17'd32782,17'd32455,17'd30860,17'd32455,17'd31160,17'd31160,17'd32618,17'd32783,17'd32783,17'd31160,17'd30392,17'd32784,17'd32785,17'd32786,17'd32787,17'd32788,17'd32789,17'd32790,17'd32791,17'd32792,17'd32793,17'd32794,17'd32795,17'd32796,17'd32797,17'd32798,17'd32799,17'd32800,17'd32801,17'd32802,17'd32803,17'd32804,17'd32805,17'd32806,17'd32807,17'd32808,17'd32809,17'd32810,17'd32811,17'd32812,17'd32813,17'd32814,17'd32815,17'd32816,17'd32817,17'd32818,17'd32819,17'd32820,17'd32655,17'd32821,17'd32822,17'd32823,17'd32824,17'd32825,17'd32003,17'd32495,17'd32826,17'd32006,17'd27260,17'd28253,17'd28484,17'd29103,17'd24895,17'd32659,17'd23565,17'd32827,17'd30427,17'd31031,17'd32502,17'd21694,17'd32187,17'd32828,17'd23044,17'd31345,17'd32829,17'd22160,17'd22325,17'd22504,17'd32830,17'd30732,17'd25031,17'd25438,17'd31366,17'd25949,17'd28725,17'd30586,17'd31352,17'd30279,17'd32192,17'd32355,17'd32505,17'd32831,17'd32832,17'd32193,17'd32833,17'd30736,17'd31505,17'd32358,17'd32671,17'd31839,17'd32834,17'd32835,17'd32836,17'd32837,17'd29988,17'd30890,17'd32838,17'd30286,17'd28272,17'd28271,17'd27898,17'd25049,17'd32839,17'd32840,17'd32841,17'd23389,17'd32842,17'd23385,17'd24742,17'd28369,17'd32364,17'd32843,17'd32844,17'd29696,17'd26302,17'd25961,17'd25844,17'd32684,17'd25721,17'd27785,17'd32517,17'd32845,17'd32367,17'd32368,17'd26419,17'd32846,17'd30447,17'd32847,17'd28254,17'd25320,17'd25177,17'd32688,17'd25436,17'd25435,17'd32848,17'd32849,17'd32850,17'd32212,17'd32851,17'd32852,17'd32853,17'd32854,17'd32855,17'd32856,17'd32857,17'd32858,17'd32859,17'd32860,17'd32861,17'd32862,17'd32863,17'd32864,17'd32865,17'd32866,17'd32867,17'd32868,17'd32869,17'd32712,17'd32870,17'd32871,17'd32872,17'd4987,17'd32873,17'd32874,17'd9500,17'd32717,17'd4522,17'd4839,17'd5329,17'd6218,17'd6553,17'd6553,17'd6707,17'd6553,17'd6218,17'd26218,17'd26708,17'd7668,17'd28184,17'd27815,17'd10515,17'd28184,17'd9933,17'd29592,17'd29592,17'd29593,17'd27815,17'd30332,17'd30487,17'd27935,17'd32553,17'd32718,17'd6390,17'd7668,17'd27696,17'd29592,17'd28183,17'd31551,17'd32875,17'd32876,17'd32719,17'd10897,17'd27931,17'd9933,17'd10380,17'd10517,17'd8001,17'd6558,17'd6710,17'd7671,17'd7841,17'd11580,17'd26713,17'd32877,17'd3853,17'd32878,17'd32879,17'd32880,17'd32881,17'd32882,17'd1679,17'd1099,17'd421,17'd602,17'd6868,17'd6415,17'd6889,17'd5030,17'd28066,17'd27949,17'd28066,17'd28066,17'd28066,17'd31729,17'd31101,17'd31101,17'd31101,17'd27708,17'd29170,17'd29040,17'd29040,17'd29040,17'd27822,17'd27319,17'd27319,17'd31902,17'd32725,17'd28545,17'd27580,17'd29169,17'd2394,17'd1383,17'd2589,17'd2409,17'd1667,17'd1679,17'd403,17'd613,17'd435,17'd32883,17'd32884
},
'{
17'd32885,17'd5643,17'd5199,17'd5200,17'd5646,17'd3902,17'd4428,17'd4246,17'd3252,17'd2422,17'd1688,17'd1831,17'd10535,17'd10535,17'd3252,17'd1831,17'd1415,17'd2257,17'd2425,17'd2257,17'd468,17'd652,17'd980,17'd980,17'd20570,17'd7385,17'd7388,17'd7388,17'd6904,17'd9970,17'd6439,17'd26731,17'd4741,17'd5220,17'd4744,17'd32088,17'd32409,17'd32730,17'd32730,17'd31260,17'd3758,17'd24969,17'd32886,17'd32732,17'd32887,17'd14453,17'd32888,17'd4909,17'd25509,17'd32889,17'd32890,17'd32891,17'd32892,17'd32893,17'd17321,17'd32894,17'd32895,17'd15520,17'd15767,17'd15519,17'd14768,17'd15524,17'd18060,17'd17206,17'd18774,17'd19006,17'd12362,17'd17809,17'd32896,17'd32897,17'd13210,17'd17809,17'd29904,17'd16765,17'd19893,17'd32571,17'd16661,17'd32898,17'd32899,17'd32900,17'd32901,17'd31923,17'd32902,17'd32903,17'd32268,17'd32577,17'd32904,17'd32112,17'd9584,17'd9445,17'd9311,17'd9311,17'd9311,17'd11095,17'd11095,17'd19521,17'd12071,17'd8224,17'd32580,17'd32749,17'd32905,17'd32906,17'd32907,17'd32908,17'd32909,17'd32910,17'd32911,17'd32912,17'd32913,17'd32914,17'd9879,17'd32915,17'd11519,17'd11807,17'd24029,17'd11275,17'd16555,17'd11528,17'd32916,17'd8880,17'd10178,17'd10028,17'd16691,17'd17849,17'd13004,17'd10607,17'd9348,17'd15569,17'd9740,17'd13886,17'd24858,17'd27622,17'd32917,17'd32918,17'd32919,17'd31765,17'd30973,17'd32283,17'd32592,17'd32920,17'd31287,17'd30972,17'd28345,17'd25528,17'd23168,17'd11959,17'd16321,17'd11958,17'd13362,17'd10990,17'd11528,17'd19279,17'd9344,17'd9344,17'd9341,17'd9473,17'd10023,17'd17839,17'd11277,17'd9619,17'd9741,17'd11277,17'd26034,17'd10164,17'd11132,17'd11524,17'd13886,17'd10991,17'd25675,17'd25525,17'd32921,17'd32922,17'd32923,17'd32924,17'd32925,17'd30829,17'd32926,17'd32927,17'd32928,17'd32929,17'd32930,17'd32931,17'd32932,17'd32933,17'd29642,17'd26758,17'd18198,17'd12262,17'd32137,17'd32934,17'd15810,17'd12111,17'd13881,17'd30983,17'd32935,17'd32936,17'd32937,17'd32938,17'd32939,17'd32940,17'd32941,17'd32942,17'd32777,17'd28953,17'd32943,17'd32944,17'd32945,17'd32781,17'd30399,17'd32946,17'd32947,17'd32948,17'd32949,17'd31462,17'd32148,17'd31794,17'd32950,17'd31794,17'd31311,17'd32951,17'd32952,17'd32953,17'd32954,17'd32955,17'd32956,17'd32957,17'd32958,17'd32959,17'd32960,17'd32961,17'd32962,17'd32963,17'd32964,17'd32965,17'd32966,17'd32967,17'd32968,17'd32969,17'd32970,17'd32971,17'd32972,17'd32973,17'd32974,17'd32975,17'd32976,17'd32977,17'd32978,17'd32979,17'd32980,17'd32981,17'd32982,17'd32983,17'd32984,17'd32985,17'd32986,17'd32987,17'd32654,17'd32988,17'd32989,17'd32990,17'd32991,17'd32992,17'd32993,17'd32003,17'd32495,17'd32994,17'd32343,17'd32006,17'd32995,17'd32996,17'd29825,17'd25180,17'd24416,17'd23733,17'd22328,17'd22506,17'd31031,17'd32502,17'd32997,17'd22511,17'd32998,17'd32347,17'd31831,17'd31497,17'd22683,17'd32999,17'd22504,17'd32830,17'd29526,17'd28977,17'd29103,17'd33000,17'd28481,17'd27640,17'd30586,17'd29245,17'd33001,17'd32192,17'd32017,17'd32505,17'd32831,17'd32354,17'd32193,17'd29690,17'd30737,17'd32670,17'd31506,17'd32671,17'd31506,17'd29981,17'd33002,17'd32024,17'd33003,17'd27154,17'd30288,17'd33004,17'd30286,17'd28272,17'd28383,17'd33005,17'd27527,17'd32839,17'd26290,17'd33006,17'd23218,17'd33007,17'd23386,17'd24090,17'd33008,17'd33009,17'd33010,17'd33011,17'd33012,17'd33013,17'd25447,17'd25718,17'd26542,17'd25458,17'd28505,17'd33014,17'd33015,17'd32518,17'd28505,17'd28745,17'd33016,17'd33017,17'd33018,17'd24898,17'd23558,17'd27509,17'd25177,17'd31366,17'd23554,17'd25708,17'd32515,17'd27645,17'd33019,17'd33020,17'd33021,17'd33022,17'd24423,17'd33023,17'd23932,17'd33024,17'd31531,17'd33025,17'd33026,17'd33027,17'd33028,17'd33029,17'd33030,17'd33031,17'd33032,17'd33033,17'd33034,17'd6060,17'd33035,17'd33036,17'd5318,17'd33037,17'd33038,17'd8141,17'd33039,17'd32240,17'd33040,17'd33041,17'd6067,17'd4845,17'd5336,17'd5615,17'd6707,17'd6553,17'd6553,17'd6553,17'd6389,17'd26708,17'd7499,17'd8780,17'd27815,17'd10515,17'd27815,17'd9933,17'd29593,17'd29592,17'd29592,17'd10515,17'd10514,17'd30487,17'd5615,17'd31553,17'd33042,17'd6390,17'd7499,17'd9933,17'd29592,17'd27933,17'd31551,17'd31551,17'd28305,17'd32876,17'd28306,17'd29592,17'd10380,17'd10380,17'd10380,17'd8001,17'd11039,17'd6709,17'd30032,17'd11433,17'd33043,17'd25881,17'd33044,17'd33045,17'd33046,17'd33047,17'd33048,17'd33049,17'd32882,17'd642,17'd2116,17'd415,17'd1383,17'd2393,17'd5630,17'd3073,17'd5030,17'd33050,17'd28066,17'd33051,17'd28066,17'd28066,17'd27949,17'd27949,17'd31729,17'd31729,17'd28315,17'd27708,17'd29039,17'd29040,17'd29040,17'd29040,17'd27822,17'd27319,17'd31902,17'd2561,17'd27709,17'd27318,17'd26965,17'd2394,17'd413,17'd602,17'd1668,17'd1823,17'd607,17'd404,17'd613,17'd177,17'd32252,17'd397
},
'{
17'd32885,17'd5643,17'd5199,17'd5200,17'd5646,17'd4243,17'd6420,17'd4246,17'd3252,17'd2422,17'd1831,17'd1831,17'd10535,17'd10535,17'd3252,17'd2422,17'd2936,17'd2257,17'd2425,17'd2257,17'd468,17'd29,17'd28,17'd980,17'd20570,17'd7385,17'd7388,17'd7388,17'd6904,17'd6904,17'd6439,17'd26731,17'd4741,17'd5058,17'd4743,17'd33052,17'd33053,17'd32730,17'd33054,17'd33055,17'd3603,17'd24969,17'd32886,17'd33056,17'd22790,17'd33057,17'd33058,17'd25507,17'd18161,17'd33059,17'd33060,17'd33061,17'd33062,17'd17811,17'd14767,17'd32569,17'd32416,17'd24013,17'd15767,17'd15385,17'd16987,17'd16519,17'd19255,17'd27461,17'd20422,17'd22630,17'd14621,17'd13093,17'd21184,17'd32897,17'd13210,17'd23325,17'd24347,17'd28925,17'd27107,17'd33063,17'd33064,17'd33065,17'd32573,17'd33066,17'd33067,17'd32108,17'd33068,17'd33069,17'd33070,17'd33071,17'd32747,17'd15150,17'd9584,17'd9310,17'd9311,17'd18307,17'd9585,17'd18542,17'd18542,17'd9019,17'd8548,17'd7924,17'd32580,17'd33072,17'd33073,17'd33074,17'd33075,17'd33076,17'd33077,17'd33078,17'd33079,17'd33080,17'd32913,17'd33081,17'd10020,17'd33082,17'd11395,17'd11807,17'd19533,17'd11275,17'd19282,17'd26759,17'd32123,17'd10338,17'd12867,17'd10028,17'd16691,17'd17849,17'd10178,17'd8569,17'd9194,17'd33083,17'd9739,17'd17236,17'd33084,17'd33085,17'd33086,17'd33087,17'd31763,17'd31128,17'd32283,17'd32438,17'd33088,17'd32920,17'd30973,17'd31285,17'd27858,17'd12254,17'd21671,17'd11959,17'd16321,17'd13883,17'd11964,17'd10476,17'd14928,17'd22814,17'd10174,17'd9346,17'd10743,17'd16796,17'd10023,17'd9883,17'd12116,17'd17011,17'd9741,17'd11277,17'd17839,17'd11528,17'd11132,17'd11524,17'd10476,17'd12863,17'd29090,17'd9040,17'd23685,17'd23685,17'd33089,17'd33090,17'd33091,17'd33092,17'd33093,17'd32770,17'd32929,17'd32930,17'd33094,17'd33095,17'd33096,17'd30677,17'd28462,17'd23855,17'd12719,17'd16548,17'd33097,17'd21670,17'd14002,17'd14521,17'd33098,17'd33099,17'd30234,17'd33100,17'd33101,17'd33102,17'd33103,17'd32610,17'd33104,17'd33105,17'd33106,17'd32943,17'd32144,17'd30251,17'd29952,17'd32781,17'd33107,17'd33108,17'd30399,17'd33109,17'd32950,17'd31461,17'd33110,17'd33111,17'd33112,17'd33113,17'd33114,17'd33115,17'd33116,17'd33117,17'd33118,17'd33119,17'd33120,17'd33121,17'd33122,17'd33123,17'd33124,17'd33125,17'd33126,17'd33127,17'd33128,17'd33129,17'd33130,17'd33131,17'd33132,17'd33133,17'd33134,17'd33135,17'd33136,17'd33137,17'd33138,17'd33139,17'd33140,17'd33141,17'd33142,17'd33143,17'd33144,17'd33145,17'd33146,17'd33147,17'd32984,17'd33148,17'd32487,17'd33149,17'd33150,17'd32820,17'd32988,17'd32989,17'd33151,17'd33152,17'd33153,17'd32003,17'd32495,17'd32005,17'd32496,17'd33154,17'd33155,17'd33156,17'd33157,17'd25320,17'd24416,17'd23920,17'd33158,17'd22332,17'd33159,17'd32502,17'd32997,17'd32010,17'd33160,17'd33161,17'd33162,17'd31344,17'd22507,17'd32999,17'd22325,17'd32830,17'd29531,17'd30733,17'd31034,17'd28597,17'd30606,17'd27515,17'd33163,17'd29245,17'd33001,17'd33164,17'd32017,17'd33165,17'd28373,17'd32354,17'd32193,17'd33166,17'd30280,17'd31505,17'd32021,17'd32358,17'd31506,17'd33167,17'd30588,17'd32024,17'd33003,17'd32511,17'd30593,17'd33168,17'd30438,17'd33169,17'd33170,17'd28870,17'd27655,17'd33171,17'd33172,17'd24746,17'd30277,17'd33173,17'd23923,17'd28722,17'd31367,17'd33174,17'd33175,17'd33176,17'd33177,17'd30135,17'd33178,17'd25718,17'd26542,17'd25458,17'd28505,17'd29261,17'd32517,17'd32517,17'd29261,17'd25458,17'd33179,17'd28613,17'd33180,17'd24745,17'd24894,17'd27509,17'd28717,17'd31856,17'd26660,17'd23908,17'd30455,17'd33181,17'd31513,17'd33182,17'd28977,17'd30127,17'd33183,17'd33184,17'd33185,17'd33186,17'd33187,17'd33188,17'd33189,17'd33190,17'd33191,17'd33192,17'd33193,17'd33194,17'd33195,17'd33196,17'd33197,17'd33198,17'd33199,17'd33200,17'd33201,17'd33202,17'd33203,17'd33204,17'd33205,17'd33206,17'd33207,17'd33208,17'd5144,17'd4845,17'd5334,17'd26949,17'd9090,17'd8303,17'd8303,17'd8154,17'd26708,17'd26708,17'd7499,17'd8780,17'd9933,17'd10642,17'd10515,17'd27696,17'd29593,17'd29592,17'd29592,17'd27933,17'd10515,17'd28184,17'd6219,17'd31553,17'd33042,17'd6554,17'd7499,17'd9933,17'd27933,17'd27933,17'd31551,17'd32875,17'd33209,17'd32876,17'd28306,17'd28650,17'd9933,17'd10380,17'd10380,17'd10380,17'd11039,17'd8002,17'd7502,17'd8634,17'd33210,17'd12474,17'd10646,17'd7189,17'd33211,17'd33212,17'd33213,17'd33049,17'd32882,17'd607,17'd1099,17'd194,17'd778,17'd413,17'd12496,17'd3073,17'd5777,17'd33050,17'd33051,17'd33051,17'd31899,17'd28066,17'd28066,17'd27949,17'd31729,17'd31729,17'd28315,17'd27708,17'd29039,17'd29039,17'd29040,17'd29040,17'd29040,17'd27822,17'd27710,17'd31902,17'd28545,17'd27580,17'd29169,17'd2394,17'd413,17'd2589,17'd2409,17'd1823,17'd1679,17'd1960,17'd613,17'd19240,17'd33214,17'd397
},
'{
17'd33215,17'd5790,17'd33216,17'd4890,17'd5646,17'd4892,17'd4733,17'd4887,17'd3252,17'd2422,17'd1831,17'd10535,17'd14070,17'd14070,17'd3252,17'd1831,17'd2257,17'd2257,17'd2257,17'd2257,17'd468,17'd652,17'd980,17'd980,17'd7385,17'd7555,17'd7388,17'd7388,17'd6904,17'd6904,17'd27592,17'd12931,17'd32729,17'd5220,17'd4744,17'd32088,17'd32409,17'd32730,17'd33054,17'd33055,17'd3601,17'd31733,17'd32255,17'd33056,17'd33217,17'd2277,17'd4752,17'd25507,17'd19372,17'd15253,17'd33218,17'd33219,17'd33220,17'd17811,17'd14893,17'd33221,17'd24194,17'd15520,17'd15008,17'd32894,17'd16033,17'd18060,17'd17206,17'd18774,17'd12532,17'd12815,17'd17096,17'd13599,17'd13463,17'd32897,17'd13210,17'd33222,17'd33223,17'd19387,17'd21186,17'd31575,17'd32263,17'd33224,17'd33225,17'd33226,17'd33227,17'd32902,17'd32903,17'd33069,17'd33228,17'd33229,17'd33230,17'd15023,17'd9445,17'd9445,17'd9311,17'd9311,17'd11095,17'd11095,17'd9165,17'd9165,17'd8387,17'd8857,17'd7594,17'd33072,17'd33073,17'd33231,17'd33232,17'd33233,17'd33234,17'd33235,17'd33236,17'd32912,17'd32589,17'd31437,17'd33105,17'd10604,17'd14810,17'd14673,17'd11130,17'd17236,17'd12863,17'd33237,17'd33238,17'd12586,17'd12588,17'd17352,17'd18203,17'd17849,17'd9887,17'd8886,17'd15944,17'd9619,17'd10606,17'd14673,17'd26035,17'd29327,17'd30675,17'd33087,17'd30973,17'd31287,17'd32283,17'd32283,17'd32920,17'd32920,17'd30834,17'd28461,17'd28689,17'd12253,17'd14130,17'd13761,17'd11958,17'd16204,17'd10989,17'd10991,17'd11277,17'd10335,17'd8874,17'd10173,17'd9741,17'd9883,17'd10023,17'd9883,17'd12116,17'd10742,17'd9741,17'd9473,17'd19642,17'd20756,17'd11132,17'd10604,17'd21206,17'd19642,17'd17347,17'd18808,17'd33239,17'd32762,17'd33240,17'd33241,17'd33242,17'd31767,17'd33096,17'd32930,17'd32931,17'd32770,17'd32930,17'd33243,17'd31288,17'd30972,17'd28229,17'd12254,17'd12260,17'd33244,17'd33245,17'd33246,17'd18192,17'd32603,17'd33247,17'd30234,17'd33248,17'd33249,17'd32608,17'd33250,17'd33251,17'd33252,17'd33253,17'd33254,17'd32943,17'd33255,17'd32615,17'd33256,17'd33257,17'd30703,17'd33108,17'd30702,17'd31308,17'd33258,17'd31153,17'd33259,17'd33260,17'd33261,17'd33262,17'd33263,17'd33264,17'd32310,17'd33265,17'd33266,17'd33267,17'd33268,17'd33269,17'd33270,17'd33271,17'd33272,17'd33273,17'd33274,17'd33275,17'd33276,17'd33277,17'd33278,17'd33279,17'd33280,17'd33281,17'd33282,17'd33283,17'd33284,17'd33285,17'd33286,17'd33287,17'd33288,17'd33289,17'd33290,17'd33291,17'd33292,17'd33293,17'd33294,17'd33295,17'd33296,17'd33297,17'd33298,17'd33299,17'd33300,17'd33301,17'd33150,17'd33302,17'd33303,17'd33304,17'd33305,17'd33306,17'd33307,17'd33308,17'd32005,17'd32826,17'd33309,17'd33310,17'd33155,17'd32996,17'd28850,17'd25032,17'd29241,17'd22501,17'd33311,17'd31348,17'd33312,17'd33313,17'd22510,17'd33314,17'd33160,17'd32997,17'd32009,17'd22157,17'd32999,17'd33315,17'd33316,17'd29531,17'd33317,17'd33318,17'd28717,17'd27638,17'd26174,17'd27258,17'd31352,17'd33319,17'd32192,17'd28373,17'd33165,17'd33320,17'd32017,17'd33321,17'd29691,17'd30433,17'd32357,17'd33322,17'd32358,17'd33323,17'd33167,17'd30281,17'd32196,17'd33324,17'd29700,17'd30441,17'd30592,17'd33325,17'd33326,17'd33327,17'd28022,17'd33328,17'd33329,17'd33330,17'd33331,17'd30277,17'd33332,17'd31844,17'd23564,17'd29702,17'd33333,17'd27640,17'd33334,17'd33335,17'd33336,17'd25586,17'd25576,17'd25967,17'd32368,17'd33337,17'd27904,17'd27785,17'd27665,17'd32517,17'd28505,17'd25718,17'd33338,17'd29549,17'd33339,17'd33340,17'd23558,17'd33341,17'd31213,17'd33342,17'd26174,17'd32843,17'd33343,17'd33344,17'd33345,17'd24081,17'd24084,17'd33346,17'd33347,17'd33348,17'd33349,17'd33350,17'd33351,17'd33352,17'd33353,17'd33354,17'd33355,17'd33356,17'd33357,17'd33358,17'd33359,17'd33360,17'd33361,17'd33362,17'd5906,17'd33201,17'd33363,17'd4182,17'd33364,17'd4522,17'd33365,17'd33208,17'd33366,17'd33367,17'd32552,17'd29739,17'd26949,17'd6391,17'd7668,17'd7668,17'd6220,17'd6390,17'd6554,17'd6390,17'd7668,17'd27815,17'd10515,17'd27815,17'd27815,17'd29593,17'd29593,17'd29592,17'd27933,17'd10515,17'd10514,17'd6391,17'd31717,17'd33368,17'd33369,17'd7499,17'd8780,17'd9933,17'd28183,17'd31551,17'd31551,17'd28305,17'd32876,17'd28305,17'd28306,17'd29592,17'd29592,17'd10516,17'd9934,17'd10238,17'd6558,17'd6561,17'd7503,17'd12310,17'd12168,17'd33370,17'd5769,17'd33371,17'd33372,17'd33373,17'd27092,17'd33374,17'd608,17'd1099,17'd778,17'd1672,17'd33375,17'd2393,17'd14178,17'd5183,17'd11061,17'd33051,17'd33051,17'd33051,17'd33051,17'd28066,17'd27949,17'd31729,17'd31101,17'd27708,17'd29170,17'd29039,17'd29039,17'd29039,17'd29040,17'd29040,17'd29040,17'd27710,17'd28545,17'd27709,17'd27318,17'd26965,17'd2394,17'd413,17'd414,17'd11062,17'd3743,17'd607,17'd442,17'd1397,17'd436,17'd33376,17'd33377
},
'{
17'd10397,17'd6421,17'd30047,17'd32728,17'd4425,17'd4892,17'd4733,17'd4887,17'd2422,17'd2422,17'd1831,17'd10535,17'd14070,17'd14070,17'd3252,17'd2422,17'd2597,17'd2257,17'd2257,17'd2257,17'd468,17'd29,17'd652,17'd980,17'd7385,17'd7555,17'd7388,17'd7388,17'd6904,17'd10408,17'd6279,17'd12931,17'd4741,17'd5058,17'd4743,17'd32409,17'd4260,17'd4260,17'd33378,17'd33055,17'd3267,17'd24334,17'd2952,17'd2444,17'd32091,17'd27103,17'd21030,17'd14995,17'd18878,17'd15754,17'd32891,17'd33379,17'd33380,17'd14893,17'd15519,17'd33381,17'd24194,17'd14893,17'd15008,17'd24012,17'd17445,17'd21185,17'd18655,17'd19382,17'd13969,17'd13211,17'd13093,17'd13093,17'd13209,17'd19890,17'd13210,17'd33222,17'd33382,17'd33383,17'd33384,17'd33385,17'd32742,17'd33224,17'd33386,17'd33387,17'd33388,17'd33389,17'd33069,17'd32268,17'd33390,17'd33391,17'd33392,17'd15023,17'd9445,17'd9445,17'd9311,17'd9311,17'd11095,17'd11095,17'd9165,17'd8387,17'd7922,17'd33393,17'd8859,17'd33072,17'd33394,17'd33395,17'd33396,17'd33397,17'd33398,17'd33399,17'd33400,17'd32912,17'd32589,17'd10592,17'd33401,17'd17236,17'd13138,17'd10990,17'd14132,17'd10476,17'd11135,17'd32916,17'd25531,17'd12724,17'd8419,17'd16691,17'd17609,17'd17849,17'd11531,17'd25677,17'd24361,17'd11277,17'd10476,17'd17478,17'd26494,17'd33402,17'd30833,17'd33403,17'd31287,17'd31287,17'd32283,17'd31287,17'd32920,17'd31127,17'd31439,17'd28345,17'd18084,17'd12109,17'd13761,17'd11960,17'd13135,17'd12262,17'd10854,17'd11134,17'd9479,17'd9743,17'd14811,17'd15807,17'd9741,17'd9883,17'd17719,17'd16796,17'd10742,17'd10742,17'd10856,17'd9740,17'd11135,17'd19155,17'd14518,17'd10476,17'd19282,17'd21669,17'd33404,17'd9745,17'd33405,17'd33406,17'd33407,17'd33408,17'd32133,17'd33409,17'd33243,17'd32930,17'd32931,17'd33096,17'd33096,17'd31288,17'd30973,17'd29067,17'd27121,17'd15570,17'd33410,17'd30841,17'd33411,17'd33412,17'd30086,17'd33413,17'd33414,17'd33415,17'd33416,17'd33417,17'd33418,17'd33419,17'd33420,17'd33421,17'd33422,17'd29508,17'd29952,17'd30250,17'd32781,17'd33257,17'd30858,17'd31157,17'd33423,17'd33424,17'd33425,17'd33426,17'd33427,17'd33428,17'd33429,17'd33430,17'd32151,17'd33431,17'd33432,17'd33433,17'd33434,17'd33435,17'd33436,17'd33437,17'd33438,17'd33439,17'd33440,17'd33441,17'd33442,17'd33443,17'd33444,17'd33445,17'd33446,17'd33447,17'd33448,17'd33449,17'd33450,17'd33451,17'd33452,17'd33453,17'd33454,17'd33455,17'd33456,17'd33457,17'd33458,17'd33459,17'd33460,17'd33461,17'd33462,17'd33463,17'd33464,17'd33465,17'd33466,17'd33467,17'd33468,17'd33469,17'd33470,17'd33471,17'd33472,17'd33473,17'd33151,17'd33152,17'd33474,17'd33307,17'd33475,17'd33476,17'd32994,17'd32826,17'd33477,17'd33478,17'd28483,17'd29970,17'd25032,17'd29375,17'd32351,17'd22678,17'd33479,17'd33480,17'd31192,17'd32011,17'd33481,17'd33314,17'd31660,17'd32829,17'd30580,17'd22324,17'd33315,17'd33316,17'd32352,17'd33482,17'd33483,17'd33484,17'd28599,17'd26174,17'd27258,17'd30735,17'd30279,17'd32192,17'd28134,17'd33485,17'd33165,17'd32017,17'd33321,17'd33486,17'd29978,17'd30736,17'd33487,17'd32358,17'd33488,17'd33489,17'd30434,17'd33490,17'd33491,17'd29989,17'd33492,17'd33493,17'd29985,17'd29696,17'd29110,17'd33494,17'd29128,17'd33329,17'd33495,17'd33496,17'd30277,17'd33497,17'd33498,17'd23564,17'd29548,17'd30456,17'd33499,17'd33500,17'd33501,17'd33502,17'd33503,17'd26074,17'd27162,17'd32368,17'd33337,17'd27904,17'd28505,17'd27785,17'd32517,17'd27785,17'd25721,17'd25040,17'd33504,17'd33505,17'd24898,17'd23558,17'd33341,17'd33506,17'd33507,17'd26174,17'd33508,17'd33509,17'd33510,17'd28850,17'd26899,17'd24901,17'd33511,17'd33512,17'd33513,17'd33514,17'd33515,17'd33516,17'd33517,17'd33518,17'd33519,17'd33520,17'd33521,17'd33522,17'd33523,17'd33524,17'd33525,17'd33526,17'd33527,17'd7320,17'd33528,17'd33529,17'd33530,17'd33531,17'd4676,17'd33532,17'd33533,17'd33534,17'd4187,17'd4840,17'd29739,17'd26949,17'd6391,17'd7668,17'd7668,17'd7499,17'd32073,17'd6554,17'd6390,17'd6220,17'd8780,17'd10515,17'd10515,17'd27815,17'd29593,17'd29593,17'd29592,17'd29592,17'd10515,17'd10515,17'd8780,17'd6554,17'd31553,17'd30333,17'd6219,17'd7668,17'd9933,17'd27933,17'd31551,17'd31551,17'd28305,17'd32876,17'd28305,17'd28306,17'd29592,17'd29593,17'd10380,17'd9934,17'd10238,17'd6558,17'd6561,17'd29433,17'd7184,17'd11859,17'd33370,17'd4544,17'd33535,17'd33536,17'd33537,17'd33538,17'd33539,17'd609,17'd192,17'd194,17'd777,17'd941,17'd12644,17'd2098,17'd5183,17'd2906,17'd11882,17'd33051,17'd33051,17'd33051,17'd28066,17'd27949,17'd31729,17'd31101,17'd27708,17'd29170,17'd29039,17'd29039,17'd29039,17'd29040,17'd29040,17'd29040,17'd27710,17'd28545,17'd27580,17'd26228,17'd29169,17'd2394,17'd413,17'd414,17'd11062,17'd3743,17'd607,17'd442,17'd1397,17'd218,17'd33540,17'd33377
},
'{
17'd5053,17'd5199,17'd30047,17'd32728,17'd4425,17'd4892,17'd4733,17'd4887,17'd2422,17'd2422,17'd1831,17'd10535,17'd14070,17'd14070,17'd3252,17'd1831,17'd2257,17'd2257,17'd2257,17'd2257,17'd468,17'd652,17'd980,17'd27,17'd7385,17'd7555,17'd7388,17'd7388,17'd6904,17'd10408,17'd6279,17'd5809,17'd5215,17'd26235,17'd33541,17'd25791,17'd4436,17'd4260,17'd30811,17'd33542,17'd33543,17'd24181,17'd33544,17'd2444,17'd32091,17'd3116,17'd5233,17'd25119,17'd33545,17'd33060,17'd33061,17'd33546,17'd33547,17'd33548,17'd33549,17'd33381,17'd14893,17'd15008,17'd24521,17'd16411,17'd17319,17'd16986,17'd19753,17'd12681,17'd14764,17'd12955,17'd13093,17'd13093,17'd13599,17'd13210,17'd13599,17'd33550,17'd19755,17'd6768,17'd33551,17'd33552,17'd33553,17'd33554,17'd33555,17'd32901,17'd33556,17'd33557,17'd33069,17'd32423,17'd32577,17'd33558,17'd33559,17'd9444,17'd10570,17'd10570,17'd9311,17'd9311,17'd11095,17'd11095,17'd12370,17'd12370,17'd8702,17'd8224,17'd7594,17'd33072,17'd33394,17'd33560,17'd33561,17'd33562,17'd33563,17'd33564,17'd33565,17'd32912,17'd10720,17'd33566,17'd27002,17'd17236,17'd17236,17'd21206,17'd19281,17'd11133,17'd11276,17'd32123,17'd23861,17'd13139,17'd9888,17'd8581,17'd7949,17'd9888,17'd8572,17'd15684,17'd15569,17'd11134,17'd17236,17'd14259,17'd24857,17'd30526,17'd32919,17'd33567,17'd32592,17'd32592,17'd33568,17'd31288,17'd31441,17'd31765,17'd29067,17'd28104,17'd25671,17'd14130,17'd13761,17'd11806,17'd13362,17'd11965,17'd19532,17'd21503,17'd9340,17'd9743,17'd15807,17'd14674,17'd12116,17'd11277,17'd9741,17'd11136,17'd9480,17'd10742,17'd9740,17'd17839,17'd11276,17'd19155,17'd10478,17'd11133,17'd10479,17'd32123,17'd12587,17'd33569,17'd33570,17'd33571,17'd33572,17'd33573,17'd31765,17'd33574,17'd33243,17'd32930,17'd33096,17'd33575,17'd33409,17'd33576,17'd30972,17'd28818,17'd25279,17'd14670,17'd33577,17'd33578,17'd32448,17'd33579,17'd31139,17'd33580,17'd33581,17'd33582,17'd33583,17'd33418,17'd33419,17'd33420,17'd33584,17'd33585,17'd33586,17'd33587,17'd32454,17'd32949,17'd30397,17'd31463,17'd30701,17'd33588,17'd33589,17'd33590,17'd33591,17'd33592,17'd33593,17'd33594,17'd33595,17'd33596,17'd33597,17'd33598,17'd33599,17'd33600,17'd33601,17'd33602,17'd33603,17'd33604,17'd33605,17'd33606,17'd33607,17'd33608,17'd33609,17'd33610,17'd33611,17'd33612,17'd33613,17'd33614,17'd33615,17'd33616,17'd33617,17'd33618,17'd33619,17'd33620,17'd33621,17'd33622,17'd33623,17'd33624,17'd33625,17'd33626,17'd33627,17'd33628,17'd33629,17'd33630,17'd33631,17'd33632,17'd33466,17'd33633,17'd33634,17'd33635,17'd33636,17'd33637,17'd33471,17'd33638,17'd33303,17'd33639,17'd33305,17'd33640,17'd33641,17'd31654,17'd32004,17'd32826,17'd33154,17'd27260,17'd33642,17'd33643,17'd32353,17'd33644,17'd23736,17'd32827,17'd33645,17'd23394,17'd31658,17'd21695,17'd33646,17'd33647,17'd33648,17'd33649,17'd32497,17'd33650,17'd22326,17'd33316,17'd33651,17'd33652,17'd33653,17'd28719,17'd31366,17'd27766,17'd28853,17'd31035,17'd29977,17'd33319,17'd32832,17'd33485,17'd33165,17'd33654,17'd33655,17'd33656,17'd29979,17'd30130,17'd33487,17'd33487,17'd33489,17'd33489,17'd31037,17'd32672,17'd32673,17'd29989,17'd33492,17'd30592,17'd30454,17'd33657,17'd28605,17'd28376,17'd33658,17'd33329,17'd33495,17'd33659,17'd32513,17'd33660,17'd33661,17'd23565,17'd31512,17'd25951,17'd27883,17'd33500,17'd33662,17'd33663,17'd33169,17'd25966,17'd26081,17'd32368,17'd26671,17'd28276,17'd27904,17'd27785,17'd32517,17'd29393,17'd27784,17'd33664,17'd33665,17'd25711,17'd33666,17'd25179,17'd31367,17'd33667,17'd33668,17'd32364,17'd33669,17'd33670,17'd33671,17'd27765,17'd23557,17'd33672,17'd33673,17'd33674,17'd33675,17'd33676,17'd33677,17'd33678,17'd33679,17'd33680,17'd33681,17'd33682,17'd33683,17'd33684,17'd33685,17'd21432,17'd33686,17'd10497,17'd33687,17'd33527,17'd33688,17'd33689,17'd33690,17'd33038,17'd5755,17'd5144,17'd4515,17'd33533,17'd33691,17'd4525,17'd33692,17'd26828,17'd8780,17'd27696,17'd27696,17'd27696,17'd7499,17'd9091,17'd6390,17'd6219,17'd8780,17'd10515,17'd10642,17'd27933,17'd9933,17'd9933,17'd9933,17'd27815,17'd27933,17'd10515,17'd28184,17'd6220,17'd30333,17'd31553,17'd6390,17'd7668,17'd9933,17'd27933,17'd31551,17'd31551,17'd32875,17'd32875,17'd28305,17'd28306,17'd29592,17'd31718,17'd10380,17'd9934,17'd7177,17'd6558,17'd6561,17'd7016,17'd33693,17'd11858,17'd20700,17'd5346,17'd24318,17'd33694,17'd33695,17'd33538,17'd763,17'd30342,17'd410,17'd780,17'd777,17'd1671,17'd15233,17'd14586,17'd4559,17'd2906,17'd11882,17'd33051,17'd33051,17'd33051,17'd28066,17'd27949,17'd31729,17'd31101,17'd31101,17'd31101,17'd29170,17'd29170,17'd29039,17'd29039,17'd29040,17'd29040,17'd28546,17'd28545,17'd27580,17'd1949,17'd26965,17'd2394,17'd413,17'd2589,17'd11062,17'd3743,17'd607,17'd442,17'd33696,17'd218,17'd33540,17'd33377
},
'{
17'd6421,17'd5200,17'd29756,17'd32728,17'd4425,17'd4892,17'd4733,17'd4887,17'd2422,17'd2422,17'd1831,17'd10535,17'd14070,17'd14070,17'd3252,17'd2422,17'd2597,17'd2257,17'd2257,17'd2257,17'd468,17'd29,17'd28,17'd27,17'd7385,17'd7555,17'd7388,17'd7556,17'd10408,17'd10408,17'd6279,17'd12931,17'd4740,17'd5217,17'd4584,17'd4436,17'd4260,17'd33378,17'd31732,17'd3603,17'd24334,17'd2952,17'd33056,17'd2273,17'd14453,17'd33697,17'd5234,17'd33698,17'd33059,17'd33218,17'd33219,17'd33699,17'd32101,17'd33548,17'd33549,17'd33221,17'd14892,17'd32739,17'd18059,17'd17690,17'd21185,17'd18774,17'd19382,17'd13969,17'd12955,17'd13599,17'd12813,17'd12813,17'd13599,17'd17096,17'd23325,17'd33700,17'd20150,17'd33384,17'd33701,17'd32899,17'd33702,17'd33703,17'd33704,17'd33705,17'd33557,17'd32903,17'd32268,17'd33706,17'd32577,17'd33707,17'd15023,17'd9444,17'd10570,17'd10570,17'd9311,17'd11095,17'd11095,17'd9165,17'd12370,17'd8548,17'd8078,17'd8079,17'd8859,17'd33072,17'd33394,17'd33708,17'd33709,17'd33710,17'd8712,17'd33711,17'd33565,17'd33712,17'd33713,17'd10314,17'd10606,17'd33714,17'd33714,17'd19282,17'd10328,17'd11134,17'd19531,17'd24366,17'd22473,17'd33715,17'd8581,17'd33716,17'd8253,17'd8419,17'd24368,17'd17480,17'd11809,17'd11670,17'd11396,17'd24539,17'd29065,17'd33717,17'd33718,17'd33719,17'd32592,17'd32592,17'd33720,17'd33721,17'd33576,17'd31440,17'd28571,17'd27121,17'd22819,17'd14130,17'd11960,17'd12996,17'd10989,17'd10739,17'd9883,17'd11136,17'd23679,17'd10335,17'd10173,17'd9480,17'd16549,17'd11277,17'd10742,17'd9340,17'd9344,17'd24037,17'd25673,17'd17839,17'd10331,17'd14668,17'd14134,17'd11528,17'd33722,17'd15684,17'd33723,17'd33569,17'd33724,17'd33725,17'd33726,17'd29785,17'd33727,17'd33095,17'd33728,17'd33729,17'd33730,17'd33731,17'd33732,17'd33733,17'd29330,17'd28103,17'd12417,17'd33734,17'd33418,17'd32448,17'd33249,17'd30085,17'd30084,17'd32936,17'd33735,17'd33736,17'd33737,17'd33419,17'd33097,17'd33738,17'd10600,17'd33422,17'd33739,17'd30252,17'd32782,17'd31621,17'd32456,17'd33740,17'd30700,17'd33741,17'd33742,17'd33743,17'd33592,17'd33428,17'd33594,17'd33744,17'd33745,17'd33746,17'd33747,17'd33748,17'd33749,17'd33750,17'd33751,17'd33752,17'd33753,17'd33754,17'd33755,17'd33756,17'd33757,17'd33758,17'd33759,17'd33612,17'd33760,17'd33761,17'd33762,17'd33763,17'd33764,17'd33765,17'd33766,17'd33767,17'd33768,17'd33769,17'd33770,17'd33771,17'd33772,17'd33773,17'd33774,17'd33775,17'd33776,17'd33777,17'd33778,17'd33779,17'd33780,17'd33632,17'd33781,17'd33782,17'd33634,17'd33468,17'd33783,17'd33784,17'd33470,17'd33472,17'd33473,17'd33785,17'd33786,17'd33787,17'd33788,17'd33789,17'd33790,17'd33791,17'd32496,17'd32006,17'd33792,17'd28253,17'd31034,17'd33793,17'd33794,17'd23215,17'd33795,17'd30728,17'd32502,17'd33796,17'd33797,17'd33647,17'd33798,17'd31497,17'd30727,17'd33650,17'd22326,17'd33799,17'd33800,17'd33801,17'd33802,17'd25029,17'd33803,17'd25566,17'd28978,17'd28486,17'd29977,17'd33319,17'd27885,17'd32831,17'd33165,17'd33654,17'd33655,17'd33656,17'd29690,17'd29978,17'd33487,17'd33487,17'd31506,17'd33489,17'd31037,17'd32835,17'd33804,17'd33805,17'd29700,17'd31199,17'd33806,17'd33807,17'd33808,17'd28145,17'd33809,17'd24752,17'd33810,17'd33811,17'd32030,17'd32191,17'd33812,17'd33813,17'd28851,17'd33814,17'd33815,17'd26781,17'd33816,17'd33501,17'd33817,17'd31854,17'd27161,17'd26671,17'd26671,17'd32368,17'd27904,17'd29261,17'd32517,17'd28620,17'd25731,17'd25737,17'd33818,17'd29257,17'd33180,17'd29842,17'd25318,17'd25437,17'd33506,17'd26661,17'd26287,17'd27028,17'd33819,17'd30456,17'd24244,17'd24740,17'd23920,17'd33820,17'd33821,17'd33822,17'd33823,17'd33824,17'd33825,17'd33826,17'd33827,17'd33828,17'd33829,17'd33830,17'd33831,17'd21279,17'd30932,17'd33832,17'd6063,17'd33833,17'd33834,17'd33835,17'd33836,17'd4183,17'd33837,17'd6067,17'd33838,17'd33839,17'd33840,17'd33841,17'd27570,17'd27081,17'd28184,17'd29593,17'd29593,17'd29593,17'd27696,17'd7499,17'd6390,17'd6390,17'd7668,17'd10515,17'd28183,17'd27933,17'd27815,17'd9933,17'd9933,17'd9933,17'd29592,17'd27933,17'd27815,17'd6391,17'd28185,17'd5004,17'd27935,17'd7668,17'd27815,17'd31243,17'd30933,17'd31551,17'd32875,17'd32875,17'd28305,17'd28306,17'd29592,17'd31718,17'd10380,17'd9934,17'd7177,17'd7011,17'd8156,17'd8003,17'd7184,17'd19990,17'd20700,17'd33842,17'd23638,17'd33843,17'd33844,17'd33845,17'd33846,17'd9102,17'd1962,17'd7027,17'd26965,17'd33847,17'd15233,17'd15233,17'd5631,17'd12495,17'd11882,17'd33051,17'd33051,17'd33051,17'd28066,17'd28066,17'd31729,17'd31729,17'd31101,17'd31101,17'd29170,17'd29170,17'd29039,17'd29039,17'd29040,17'd29040,17'd28546,17'd28545,17'd27580,17'd26228,17'd29169,17'd2394,17'd1383,17'd2589,17'd11062,17'd3743,17'd607,17'd442,17'd33696,17'd585,17'd33848,17'd33377
},
'{
17'd5200,17'd5200,17'd4426,17'd4425,17'd27713,17'd25384,17'd2935,17'd2784,17'd2422,17'd2422,17'd1831,17'd10535,17'd14070,17'd14070,17'd2935,17'd2422,17'd2597,17'd2257,17'd2257,17'd2257,17'd468,17'd652,17'd27,17'd27,17'd7385,17'd7555,17'd7388,17'd6600,17'd6441,17'd10672,17'd27445,17'd26605,17'd5380,17'd33849,17'd25791,17'd4436,17'd33378,17'd33850,17'd33851,17'd3440,17'd24181,17'd33852,17'd30199,17'd32887,17'd2132,17'd26242,17'd4909,17'd33853,17'd33854,17'd33855,17'd33379,17'd33856,17'd32101,17'd33857,17'd33857,17'd31918,17'd14892,17'd32894,17'd24685,17'd17207,17'd16986,17'd17941,17'd12681,17'd14764,17'd13209,17'd13209,17'd12813,17'd13093,17'd17096,17'd17096,17'd33858,17'd33859,17'd7408,17'd33551,17'd33860,17'd33861,17'd33702,17'd33386,17'd33862,17'd33863,17'd33557,17'd33069,17'd33864,17'd33390,17'd33865,17'd31928,17'd9583,17'd9445,17'd10570,17'd10570,17'd11095,17'd11095,17'd9165,17'd9165,17'd12370,17'd8548,17'd7924,17'd8388,17'd33866,17'd31428,17'd33394,17'd33867,17'd33868,17'd33869,17'd33870,17'd33711,17'd33565,17'd30966,17'd33871,17'd33872,17'd10991,17'd24364,17'd20610,17'd19280,17'd16796,17'd17839,17'd19279,17'd33873,17'd8573,17'd8102,17'd8420,17'd33874,17'd8253,17'd8580,17'd8569,17'd10173,17'd12116,17'd21206,17'd23513,17'd24209,17'd26757,17'd30971,17'd31765,17'd31287,17'd32592,17'd32592,17'd33875,17'd33721,17'd33733,17'd29067,17'd27857,17'd24991,17'd21671,17'd14130,17'd11960,17'd13762,17'd10854,17'd11133,17'd9741,17'd23679,17'd9339,17'd9345,17'd9620,17'd9479,17'd16549,17'd16549,17'd9345,17'd9339,17'd13887,17'd24037,17'd33876,17'd9739,17'd11670,17'd14134,17'd11400,17'd17599,17'd33877,17'd8247,17'd16563,17'd33878,17'd33879,17'd33880,17'd31947,17'd31597,17'd33881,17'd33882,17'd33728,17'd33728,17'd33730,17'd33883,17'd33409,17'd33884,17'd28462,17'd23511,17'd12856,17'd30685,17'd33578,17'd32295,17'd33248,17'd30234,17'd30084,17'd33885,17'd33582,17'd33736,17'd30088,17'd33886,17'd33887,17'd33421,17'd33888,17'd29495,17'd33889,17'd30399,17'd30399,17'd33257,17'd31463,17'd33890,17'd33891,17'd33892,17'd33893,17'd33894,17'd33895,17'd33896,17'd33897,17'd32786,17'd33898,17'd33899,17'd33119,17'd33900,17'd33901,17'd33902,17'd33903,17'd33904,17'd33905,17'd33906,17'd33907,17'd33908,17'd33909,17'd33910,17'd33911,17'd33912,17'd33913,17'd33914,17'd33915,17'd33916,17'd33917,17'd33918,17'd33919,17'd33920,17'd33921,17'd33917,17'd33922,17'd33923,17'd33924,17'd33925,17'd33926,17'd33927,17'd33928,17'd33929,17'd33930,17'd33931,17'd33932,17'd33933,17'd33467,17'd33934,17'd33935,17'd33468,17'd33936,17'd33783,17'd33470,17'd33472,17'd33473,17'd33303,17'd33937,17'd33938,17'd33939,17'd33940,17'd33476,17'd33941,17'd32826,17'd33942,17'd31827,17'd25565,17'd25317,17'd32668,17'd33652,17'd29829,17'd33943,17'd33944,17'd33945,17'd33796,17'd33946,17'd33947,17'd23044,17'd31497,17'd30727,17'd33948,17'd33315,17'd33949,17'd32680,17'd33950,17'd33802,17'd28596,17'd33951,17'd25435,17'd28724,17'd26901,17'd33952,17'd33319,17'd27885,17'd32831,17'd33165,17'd32017,17'd33321,17'd29248,17'd28857,17'd29831,17'd30885,17'd33487,17'd31506,17'd33323,17'd29981,17'd33953,17'd33954,17'd33805,17'd29700,17'd31199,17'd33806,17'd33955,17'd33956,17'd33957,17'd33958,17'd33959,17'd33960,17'd33961,17'd32030,17'd30128,17'd33962,17'd33813,17'd24416,17'd30903,17'd26530,17'd33963,17'd28486,17'd33964,17'd33965,17'd30758,17'd26074,17'd26671,17'd26671,17'd32368,17'd27904,17'd28505,17'd27785,17'd31208,17'd27784,17'd25579,17'd25049,17'd33966,17'd33967,17'd33968,17'd33969,17'd25438,17'd28480,17'd25435,17'd25708,17'd27028,17'd27028,17'd33970,17'd23723,17'd23726,17'd24090,17'd33971,17'd33972,17'd33973,17'd33974,17'd33975,17'd33976,17'd33977,17'd33978,17'd33979,17'd33980,17'd33981,17'd33982,17'd21581,17'd33983,17'd33984,17'd33985,17'd33986,17'd33987,17'd33988,17'd33989,17'd33990,17'd4361,17'd4836,17'd4836,17'd33991,17'd33691,17'd33992,17'd5157,17'd29159,17'd28184,17'd29592,17'd29592,17'd29593,17'd9933,17'd7668,17'd6219,17'd6390,17'd7499,17'd10514,17'd11037,17'd28183,17'd27815,17'd9933,17'd9933,17'd9933,17'd29592,17'd10515,17'd28184,17'd28058,17'd27935,17'd5004,17'd28185,17'd6391,17'd29592,17'd30933,17'd33993,17'd30934,17'd32875,17'd32875,17'd28305,17'd27933,17'd10516,17'd10380,17'd10380,17'd9934,17'd7011,17'd8630,17'd6395,17'd7016,17'd33693,17'd11435,17'd11436,17'd33842,17'd33994,17'd33995,17'd33996,17'd33997,17'd33998,17'd33999,17'd16858,17'd6888,17'd27094,17'd33847,17'd34000,17'd12644,17'd14586,17'd34001,17'd11882,17'd33051,17'd34002,17'd34002,17'd28066,17'd28066,17'd31729,17'd31729,17'd31101,17'd31101,17'd29170,17'd29170,17'd29039,17'd29039,17'd29039,17'd29039,17'd28546,17'd28545,17'd27580,17'd1949,17'd26965,17'd2394,17'd15233,17'd2589,17'd11062,17'd3743,17'd1539,17'd442,17'd33696,17'd585,17'd33848,17'd34003
},
'{
17'd5200,17'd5200,17'd4426,17'd4426,17'd3902,17'd4428,17'd2593,17'd2784,17'd2422,17'd2422,17'd10535,17'd27714,17'd14188,17'd14070,17'd2935,17'd2422,17'd2597,17'd2257,17'd2257,17'd2257,17'd468,17'd29,17'd28,17'd27,17'd7385,17'd7388,17'd6600,17'd6904,17'd10672,17'd27592,17'd27445,17'd34004,17'd5380,17'd4584,17'd4436,17'd4260,17'd33850,17'd34005,17'd34006,17'd32254,17'd34007,17'd34008,17'd2444,17'd34009,17'd34010,17'd16013,17'd25796,17'd34011,17'd25393,17'd34012,17'd34013,17'd34014,17'd16029,17'd33857,17'd33857,17'd16029,17'd14892,17'd32739,17'd16411,17'd16289,17'd16986,17'd19382,17'd16765,17'd13211,17'd13209,17'd13968,17'd13092,17'd13093,17'd13211,17'd34015,17'd33550,17'd19388,17'd34016,17'd34017,17'd34018,17'd34019,17'd33861,17'd34020,17'd34021,17'd34022,17'd34023,17'd32576,17'd33228,17'd33390,17'd34024,17'd15150,17'd9445,17'd9445,17'd10570,17'd10570,17'd11095,17'd11095,17'd9165,17'd9165,17'd8387,17'd8702,17'd8224,17'd34025,17'd34026,17'd31428,17'd32581,17'd34027,17'd34028,17'd34029,17'd34030,17'd34031,17'd33565,17'd34032,17'd34033,17'd34034,17'd10991,17'd34035,17'd12721,17'd10330,17'd16796,17'd22131,17'd16065,17'd33238,17'd14135,17'd8103,17'd33716,17'd34036,17'd16566,17'd19780,17'd25677,17'd10334,17'd9883,17'd11398,17'd24706,17'd24857,17'd28106,17'd30832,17'd31941,17'd31442,17'd33088,17'd31766,17'd34037,17'd31288,17'd31765,17'd28571,17'd26629,17'd12255,17'd21671,17'd13761,17'd11961,17'd14262,17'd11132,17'd9883,17'd9480,17'd9191,17'd9339,17'd9620,17'd10743,17'd17011,17'd16549,17'd14674,17'd8874,17'd9189,17'd12117,17'd25525,17'd23857,17'd9739,17'd11400,17'd12584,17'd11525,17'd34038,17'd34039,17'd25813,17'd34040,17'd34041,17'd34042,17'd34043,17'd29930,17'd32930,17'd33243,17'd34044,17'd34045,17'd34046,17'd34047,17'd33881,17'd31289,17'd31285,17'd27857,17'd14003,17'd34048,17'd33419,17'd33578,17'd31140,17'd31449,17'd30234,17'd32606,17'd33736,17'd33582,17'd31140,17'd34049,17'd30090,17'd34050,17'd10020,17'd34051,17'd34052,17'd33108,17'd34053,17'd34053,17'd33107,17'd30550,17'd34054,17'd34055,17'd33893,17'd33893,17'd34056,17'd33428,17'd34057,17'd34058,17'd34059,17'd34060,17'd34061,17'd34062,17'd34063,17'd34064,17'd33903,17'd34065,17'd34066,17'd34067,17'd34068,17'd34069,17'd34070,17'd34071,17'd34072,17'd34073,17'd34074,17'd33768,17'd34075,17'd34076,17'd34077,17'd34078,17'd34079,17'd33917,17'd34080,17'd34080,17'd34081,17'd34082,17'd34083,17'd34084,17'd34085,17'd34086,17'd34087,17'd34088,17'd34089,17'd34090,17'd34091,17'd34092,17'd34093,17'd34094,17'd33781,17'd34094,17'd34095,17'd33936,17'd34096,17'd34097,17'd34098,17'd34099,17'd34099,17'd34100,17'd34101,17'd34102,17'd34103,17'd34104,17'd34105,17'd32005,17'd32826,17'd32006,17'd25707,17'd28600,17'd29244,17'd34106,17'd31502,17'd30582,17'd34107,17'd34108,17'd31659,17'd34109,17'd33947,17'd34110,17'd31345,17'd23222,17'd23742,17'd34111,17'd33949,17'd33799,17'd34112,17'd34113,17'd24896,17'd28974,17'd28600,17'd25707,17'd26901,17'd33952,17'd33001,17'd27885,17'd28258,17'd33165,17'd32017,17'd33321,17'd29248,17'd28857,17'd34114,17'd34115,17'd34116,17'd32021,17'd34117,17'd29981,17'd33953,17'd33954,17'd33003,17'd32837,17'd31199,17'd33336,17'd31207,17'd34118,17'd33957,17'd34119,17'd34120,17'd34121,17'd34122,17'd34123,17'd34124,17'd34125,17'd34126,17'd32659,17'd34127,17'd28482,17'd33963,17'd26901,17'd34128,17'd34129,17'd34130,17'd28732,17'd26297,17'd32368,17'd32519,17'd31517,17'd28505,17'd31208,17'd30296,17'd28026,17'd25199,17'd28625,17'd34131,17'd34132,17'd34133,17'd25180,17'd26399,17'd23726,17'd28130,17'd25708,17'd27028,17'd34134,17'd34135,17'd23909,17'd34136,17'd24589,17'd34137,17'd34138,17'd34139,17'd23927,17'd34140,17'd34141,17'd34142,17'd34143,17'd34144,17'd34145,17'd34146,17'd34147,17'd20825,17'd34148,17'd34149,17'd34150,17'd34151,17'd3828,17'd34152,17'd34153,17'd34154,17'd4365,17'd34155,17'd34156,17'd4524,17'd34157,17'd4998,17'd4846,17'd5763,17'd27815,17'd27933,17'd30933,17'd29592,17'd9933,17'd8780,17'd6220,17'd6219,17'd7499,17'd27815,17'd28183,17'd28183,17'd10515,17'd27815,17'd9933,17'd9933,17'd29592,17'd27933,17'd27815,17'd28058,17'd5614,17'd25627,17'd28185,17'd6220,17'd29593,17'd30933,17'd34158,17'd30934,17'd32875,17'd32875,17'd28305,17'd28306,17'd27815,17'd10380,17'd9934,17'd9934,17'd7011,17'd8630,17'd6069,17'd10899,17'd8635,17'd11042,17'd34159,17'd34160,17'd34161,17'd33995,17'd34162,17'd34163,17'd34164,17'd22263,17'd2250,17'd2905,17'd2394,17'd29440,17'd34000,17'd29750,17'd14586,17'd33050,17'd33051,17'd33051,17'd34002,17'd34002,17'd28066,17'd28066,17'd31729,17'd31729,17'd31101,17'd31101,17'd29170,17'd29170,17'd29039,17'd29039,17'd29039,17'd29039,17'd28546,17'd28545,17'd27580,17'd26228,17'd29169,17'd2394,17'd12644,17'd33375,17'd34165,17'd3743,17'd1539,17'd442,17'd33696,17'd585,17'd33848,17'd34003
},
'{
17'd4890,17'd4890,17'd5646,17'd4891,17'd4243,17'd6420,17'd2935,17'd2784,17'd2422,17'd2422,17'd3252,17'd14070,17'd14188,17'd14188,17'd2935,17'd2422,17'd2596,17'd2257,17'd2257,17'd2257,17'd468,17'd652,17'd27,17'd27,17'd7385,17'd7388,17'd6600,17'd6600,17'd6440,17'd27592,17'd26731,17'd4895,17'd5216,17'd34166,17'd4436,17'd4096,17'd33850,17'd34167,17'd34168,17'd3438,17'd34007,17'd31910,17'd34169,17'd34170,17'd34010,17'd34171,17'd25655,17'd34172,17'd34173,17'd34174,17'd34175,17'd34176,17'd34177,17'd34178,17'd34179,17'd16029,17'd14893,17'd24012,17'd17448,17'd16164,17'd17205,17'd20423,17'd12362,17'd13210,17'd13462,17'd13968,17'd13092,17'd13093,17'd13094,17'd34180,17'd34181,17'd19388,17'd34182,17'd34183,17'd34184,17'd34185,17'd34186,17'd34187,17'd34188,17'd34189,17'd34190,17'd34191,17'd33228,17'd33390,17'd34192,17'd12822,17'd9445,17'd9310,17'd18786,17'd11239,17'd11239,17'd11095,17'd9165,17'd9165,17'd8387,17'd8702,17'd7267,17'd8389,17'd34026,17'd31428,17'd34193,17'd34027,17'd34194,17'd34195,17'd34196,17'd34197,17'd34198,17'd29632,17'd34199,17'd34200,17'd11132,17'd34201,17'd15176,17'd9883,17'd9741,17'd15048,17'd15569,17'd17123,17'd12867,17'd8104,17'd8253,17'd34036,17'd9622,17'd23864,17'd16071,17'd9479,17'd11134,17'd16068,17'd21363,17'd26493,17'd32128,17'd34202,17'd31765,17'd32920,17'd33088,17'd31766,17'd34037,17'd34203,17'd31440,17'd28818,17'd24704,17'd12108,17'd21671,17'd13883,17'd12260,17'd11965,17'd10165,17'd10742,17'd12117,17'd9192,17'd9339,17'd9341,17'd27003,17'd17011,17'd15187,17'd9189,17'd19033,17'd8720,17'd26626,17'd18080,17'd34204,17'd17839,17'd19282,17'd13521,17'd34205,17'd17718,17'd8571,17'd7949,17'd16688,17'd34206,17'd34207,17'd34208,17'd30372,17'd34209,17'd33094,17'd34046,17'd34210,17'd34210,17'd34211,17'd34212,17'd30221,17'd30373,17'd34213,17'd15570,17'd29793,17'd34214,17'd33250,17'd34215,17'd30085,17'd33248,17'd33582,17'd31954,17'd33736,17'd34216,17'd33245,17'd34217,17'd10160,17'd34051,17'd34218,17'd31302,17'd34219,17'd34219,17'd34219,17'd34220,17'd34221,17'd34222,17'd33894,17'd34056,17'd34223,17'd34224,17'd34225,17'd34226,17'd34227,17'd34228,17'd34229,17'd34230,17'd34231,17'd34232,17'd34233,17'd34234,17'd34235,17'd34236,17'd34237,17'd34238,17'd34239,17'd34240,17'd34241,17'd34242,17'd34243,17'd34244,17'd34245,17'd34246,17'd34247,17'd34248,17'd34249,17'd34250,17'd34251,17'd34252,17'd34253,17'd34254,17'd34081,17'd34255,17'd34256,17'd34257,17'd34258,17'd34259,17'd34260,17'd34261,17'd34262,17'd34263,17'd34264,17'd34265,17'd34266,17'd34267,17'd34268,17'd34268,17'd34269,17'd33783,17'd34270,17'd34271,17'd33638,17'd34099,17'd34100,17'd34101,17'd34272,17'd34273,17'd34274,17'd34275,17'd33790,17'd32994,17'd33477,17'd31351,17'd28720,17'd27511,17'd34276,17'd23733,17'd34277,17'd34278,17'd34279,17'd31659,17'd34280,17'd33947,17'd32348,17'd31346,17'd22005,17'd34281,17'd34111,17'd22859,17'd31495,17'd24421,17'd34282,17'd34283,17'd34284,17'd28484,17'd26174,17'd26902,17'd29246,17'd33952,17'd31503,17'd28258,17'd33485,17'd32017,17'd33321,17'd29248,17'd32018,17'd34285,17'd34115,17'd31839,17'd33323,17'd34117,17'd34286,17'd34287,17'd34288,17'd34289,17'd34290,17'd31199,17'd33336,17'd34291,17'd33956,17'd34292,17'd34293,17'd34294,17'd34295,17'd34296,17'd34297,17'd34298,17'd26527,17'd34299,17'd23916,17'd25318,17'd34300,17'd34301,17'd26781,17'd34302,17'd34303,17'd29541,17'd32199,17'd28745,17'd28028,17'd31517,17'd31517,17'd28505,17'd34304,17'd34304,17'd34305,17'd34305,17'd34306,17'd34307,17'd34308,17'd34309,17'd25032,17'd34310,17'd25026,17'd23724,17'd27766,17'd34311,17'd33964,17'd34312,17'd24737,17'd23550,17'd34313,17'd31033,17'd34314,17'd34315,17'd34316,17'd24096,17'd34317,17'd34318,17'd34319,17'd34320,17'd34321,17'd34322,17'd34323,17'd34324,17'd34325,17'd34326,17'd33984,17'd34327,17'd4825,17'd4352,17'd34328,17'd34329,17'd34330,17'd34331,17'd34332,17'd34333,17'd33838,17'd4998,17'd4684,17'd34334,17'd28184,17'd28183,17'd30933,17'd31243,17'd9933,17'd28184,17'd6391,17'd6219,17'd7499,17'd27815,17'd28183,17'd28183,17'd10515,17'd27815,17'd9933,17'd9933,17'd29592,17'd29592,17'd27815,17'd8780,17'd5614,17'd5160,17'd28185,17'd6219,17'd31888,17'd30933,17'd34158,17'd34335,17'd31551,17'd32875,17'd28305,17'd27933,17'd10516,17'd10380,17'd9934,17'd9934,17'd7011,17'd34336,17'd6069,17'd34337,17'd8308,17'd11042,17'd34338,17'd34339,17'd34340,17'd34341,17'd34342,17'd34343,17'd34344,17'd24164,17'd1959,17'd2559,17'd14178,17'd34000,17'd33847,17'd34000,17'd14586,17'd5777,17'd11882,17'd33051,17'd34002,17'd34002,17'd34002,17'd33051,17'd28066,17'd27949,17'd31729,17'd31101,17'd29170,17'd29170,17'd29039,17'd29039,17'd29039,17'd29039,17'd28546,17'd28545,17'd27580,17'd1949,17'd26965,17'd2394,17'd12644,17'd414,17'd11337,17'd3743,17'd1539,17'd442,17'd33696,17'd31730,17'd34345,17'd34003
},
'{
17'd4890,17'd4890,17'd5646,17'd4426,17'd4892,17'd4245,17'd2935,17'd2422,17'd2422,17'd3252,17'd3252,17'd3101,17'd3251,17'd3251,17'd2935,17'd2422,17'd2596,17'd2257,17'd2257,17'd22965,17'd468,17'd652,17'd28,17'd286,17'd7061,17'd7388,17'd7388,17'd6904,17'd6439,17'd6279,17'd12931,17'd4741,17'd5217,17'd3914,17'd4256,17'd4095,17'd34167,17'd34346,17'd34347,17'd32731,17'd34348,17'd31910,17'd34349,17'd34170,17'd34350,17'd34351,17'd29045,17'd34352,17'd34353,17'd34354,17'd34355,17'd34356,17'd34177,17'd34357,17'd34179,17'd16029,17'd15008,17'd17321,17'd17320,17'd21650,17'd18774,17'd12681,17'd14621,17'd13599,17'd13462,17'd13968,17'd13092,17'd13093,17'd13094,17'd34358,17'd34359,17'd34360,17'd34361,17'd32418,17'd34362,17'd34363,17'd33225,17'd34364,17'd34365,17'd34366,17'd32576,17'd34367,17'd33706,17'd32746,17'd33559,17'd9309,17'd9584,17'd18542,17'd10818,17'd19521,17'd11239,17'd11095,17'd11095,17'd9165,17'd8387,17'd8702,17'd8388,17'd34368,17'd34026,17'd8860,17'd34369,17'd34370,17'd34371,17'd34372,17'd34373,17'd34374,17'd34375,17'd34376,17'd10458,17'd34377,17'd11133,17'd34378,17'd12585,17'd10024,17'd10742,17'd9619,17'd14674,17'd29920,17'd13005,17'd7950,17'd9889,17'd9889,17'd18203,17'd24862,17'd14811,17'd18556,17'd11400,17'd14133,17'd23170,17'd29196,17'd34379,17'd32282,17'd31287,17'd32920,17'd31766,17'd31589,17'd34380,17'd34381,17'd29330,17'd27857,17'd23681,17'd22819,17'd14130,17'd15053,17'd12262,17'd25144,17'd17719,17'd9620,17'd8874,17'd9189,17'd9346,17'd10743,17'd10743,17'd9479,17'd15944,17'd9621,17'd11530,17'd9040,17'd17964,17'd34382,17'd34204,17'd17839,17'd19282,17'd28352,17'd15176,17'd17232,17'd8248,17'd8581,17'd33878,17'd34383,17'd34384,17'd30673,17'd34385,17'd34386,17'd34387,17'd33729,17'd34388,17'd34389,17'd34211,17'd33093,17'd30220,17'd34390,17'd16556,17'd15433,17'd34391,17'd33578,17'd33737,17'd30235,17'd31449,17'd34392,17'd33583,17'd34393,17'd30088,17'd33886,17'd34394,17'd32612,17'd34395,17'd34396,17'd31302,17'd29496,17'd34397,17'd34398,17'd31301,17'd34399,17'd33424,17'd33892,17'd34400,17'd34401,17'd34402,17'd34403,17'd34404,17'd34405,17'd34406,17'd34407,17'd34408,17'd34409,17'd34410,17'd34411,17'd34412,17'd34413,17'd34414,17'd34415,17'd34416,17'd34417,17'd34418,17'd34419,17'd34420,17'd34421,17'd34422,17'd34422,17'd34423,17'd34424,17'd34425,17'd34426,17'd34426,17'd34426,17'd34426,17'd34427,17'd34428,17'd34428,17'd34429,17'd34430,17'd34431,17'd34432,17'd34433,17'd34434,17'd34435,17'd34436,17'd34437,17'd34438,17'd34439,17'd34440,17'd34441,17'd34442,17'd34268,17'd34443,17'd34444,17'd34096,17'd33784,17'd33470,17'd34098,17'd34445,17'd34446,17'd34447,17'd34448,17'd34449,17'd34450,17'd34451,17'd33790,17'd33791,17'd32185,17'd31827,17'd25565,17'd29970,17'd32668,17'd24087,17'd34452,17'd34453,17'd34454,17'd34455,17'd22512,17'd33647,17'd34456,17'd34457,17'd22010,17'd22006,17'd34111,17'd34458,17'd31495,17'd23736,17'd34459,17'd34283,17'd27763,17'd28850,17'd27766,17'd26902,17'd28980,17'd33952,17'd30279,17'd32832,17'd32355,17'd33654,17'd33321,17'd29248,17'd32018,17'd34285,17'd34115,17'd31839,17'd34460,17'd34461,17'd32508,17'd34287,17'd32024,17'd33324,17'd34290,17'd31199,17'd34462,17'd31207,17'd33956,17'd33957,17'd34293,17'd34463,17'd34464,17'd34465,17'd34297,17'd34466,17'd31359,17'd34299,17'd34467,17'd25710,17'd33174,17'd27883,17'd26782,17'd26781,17'd34468,17'd34469,17'd34470,17'd26195,17'd28028,17'd34471,17'd31517,17'd28505,17'd27904,17'd34304,17'd34472,17'd34305,17'd34473,17'd34474,17'd34475,17'd34476,17'd34477,17'd34478,17'd25026,17'd24585,17'd24242,17'd25707,17'd34479,17'd34480,17'd24891,17'd34481,17'd25026,17'd24590,17'd34482,17'd34483,17'd34139,17'd34484,17'd34485,17'd34486,17'd34487,17'd34488,17'd34489,17'd34490,17'd34491,17'd20508,17'd34492,17'd34493,17'd34494,17'd34495,17'd34496,17'd34497,17'd34498,17'd34499,17'd34500,17'd4362,17'd34332,17'd34501,17'd4999,17'd33992,17'd4684,17'd5168,17'd28184,17'd28057,17'd31551,17'd31243,17'd9933,17'd28184,17'd28058,17'd6219,17'd7499,17'd9933,17'd31551,17'd31551,17'd10515,17'd27815,17'd9933,17'd9933,17'd29593,17'd29592,17'd27933,17'd8780,17'd5614,17'd28185,17'd27935,17'd6390,17'd29740,17'd31243,17'd33993,17'd31551,17'd31551,17'd34502,17'd28305,17'd27933,17'd29592,17'd10516,17'd9934,17'd7500,17'd6223,17'd34336,17'd9093,17'd34337,17'd8635,17'd34503,17'd34504,17'd34160,17'd34505,17'd34506,17'd34507,17'd34508,17'd34509,17'd34510,17'd1257,17'd1680,17'd2393,17'd15233,17'd2560,17'd28428,17'd15233,17'd28657,17'd11882,17'd33051,17'd34002,17'd34002,17'd34002,17'd33051,17'd28066,17'd27949,17'd31729,17'd31101,17'd29170,17'd29170,17'd29039,17'd29039,17'd29039,17'd29039,17'd28545,17'd28545,17'd27580,17'd26228,17'd29169,17'd2394,17'd33375,17'd12496,17'd11337,17'd3743,17'd1539,17'd442,17'd33696,17'd585,17'd34511,17'd34003
},
'{
17'd4890,17'd4889,17'd4890,17'd29756,17'd4892,17'd6420,17'd5508,17'd7214,17'd10535,17'd3252,17'd3101,17'd3251,17'd34512,17'd3101,17'd2422,17'd1688,17'd2597,17'd2425,17'd1416,17'd26344,17'd2938,17'd28,17'd652,17'd286,17'd7061,17'd7556,17'd7557,17'd6600,17'd6904,17'd11211,17'd12507,17'd4742,17'd4092,17'd4433,17'd3915,17'd4095,17'd34167,17'd34513,17'd32731,17'd2952,17'd34514,17'd33056,17'd34169,17'd32091,17'd3116,17'd34515,17'd19744,17'd34516,17'd34517,17'd34518,17'd34519,17'd34520,17'd34521,17'd34522,17'd33548,17'd15384,17'd32894,17'd16033,17'd17319,17'd17205,17'd20423,17'd13969,17'd13211,17'd13092,17'd13462,17'd13968,17'd13209,17'd13093,17'd27458,17'd9155,17'd21486,17'd34182,17'd34523,17'd34524,17'd34525,17'd32742,17'd33555,17'd34526,17'd34527,17'd34528,17'd34529,17'd34367,17'd33390,17'd15149,17'd10291,17'd11238,17'd11095,17'd10818,17'd12071,17'd12685,17'd15273,17'd11095,17'd11095,17'd13611,17'd14359,17'd7265,17'd34530,17'd34531,17'd8227,17'd7596,17'd34532,17'd34533,17'd34534,17'd34535,17'd34536,17'd34537,17'd32279,17'd34538,17'd34539,17'd26870,17'd10606,17'd11528,17'd18556,17'd9479,17'd17011,17'd24037,17'd25408,17'd9195,17'd18203,17'd17972,17'd34540,17'd23686,17'd12426,17'd16562,17'd34541,17'd19779,17'd17236,17'd14264,17'd24705,17'd34542,17'd31940,17'd34543,17'd31589,17'd34544,17'd34545,17'd33875,17'd31289,17'd30974,17'd31768,17'd26629,17'd23515,17'd21671,17'd13761,17'd15185,17'd11274,17'd10326,17'd10992,17'd10335,17'd8874,17'd9038,17'd13887,17'd15187,17'd9345,17'd24361,17'd9045,17'd34546,17'd10027,17'd15684,17'd15180,17'd9478,17'd14928,17'd20756,17'd19532,17'd10166,17'd33083,17'd29920,17'd12588,17'd34547,17'd34548,17'd34549,17'd34550,17'd34551,17'd33730,17'd34552,17'd34553,17'd34554,17'd34555,17'd34556,17'd33882,17'd34557,17'd28944,17'd24704,17'd34558,17'd34559,17'd34560,17'd33417,17'd34215,17'd33415,17'd33416,17'd33249,17'd33737,17'd30380,17'd34561,17'd32941,17'd34562,17'd10160,17'd31783,17'd34218,17'd31147,17'd30849,17'd29496,17'd30400,17'd32145,17'd34563,17'd34564,17'd34565,17'd34566,17'd34567,17'd34568,17'd34569,17'd34570,17'd34571,17'd34572,17'd34573,17'd34574,17'd34575,17'd34576,17'd34577,17'd34578,17'd34579,17'd34580,17'd34581,17'd34582,17'd34583,17'd34584,17'd34585,17'd33920,17'd34586,17'd34587,17'd34588,17'd34589,17'd34590,17'd34591,17'd34247,17'd34592,17'd34592,17'd34593,17'd34428,17'd34594,17'd34079,17'd34251,17'd34595,17'd34596,17'd34597,17'd34598,17'd34599,17'd34600,17'd34601,17'd34602,17'd34603,17'd34604,17'd34605,17'd34606,17'd34607,17'd34608,17'd33935,17'd34609,17'd34444,17'd34610,17'd34611,17'd34098,17'd34612,17'd34100,17'd34447,17'd34272,17'd34613,17'd34449,17'd34614,17'd34105,17'd33941,17'd32826,17'd33154,17'd32995,17'd28600,17'd29244,17'd30733,17'd31502,17'd23389,17'd34111,17'd22156,17'd21695,17'd34615,17'd34616,17'd34617,17'd34618,17'd31345,17'd34619,17'd34620,17'd33949,17'd29829,17'd34621,17'd28595,17'd34622,17'd29244,17'd32658,17'd28724,17'd28486,17'd29246,17'd29977,17'd33654,17'd32355,17'd32193,17'd33654,17'd32355,17'd28728,17'd29537,17'd29833,17'd30885,17'd31838,17'd34286,17'd32508,17'd30435,17'd34623,17'd33804,17'd34290,17'd30887,17'd28860,17'd34624,17'd34625,17'd34626,17'd32042,17'd34627,17'd34628,17'd34629,17'd34630,17'd24421,17'd28976,17'd34631,17'd24418,17'd24893,17'd25176,17'd24583,17'd25311,17'd26781,17'd34632,17'd34633,17'd30297,17'd26192,17'd26920,17'd26671,17'd32207,17'd28505,17'd28505,17'd27661,17'd25342,17'd28276,17'd34473,17'd34634,17'd24103,17'd34635,17'd26404,17'd34636,17'd28850,17'd23911,17'd24243,17'd26285,17'd27146,17'd34637,17'd25833,17'd25566,17'd28484,17'd24417,17'd23387,17'd34638,17'd34639,17'd34640,17'd34641,17'd30467,17'd34642,17'd34643,17'd34644,17'd34645,17'd34646,17'd34647,17'd22726,17'd21900,17'd34648,17'd34649,17'd34650,17'd34651,17'd34652,17'd34653,17'd34654,17'd34655,17'd4525,17'd34656,17'd5156,17'd34657,17'd4995,17'd5334,17'd25084,17'd11317,17'd31551,17'd30933,17'd27933,17'd28184,17'd30487,17'd28058,17'd34658,17'd27933,17'd31551,17'd31551,17'd10515,17'd28184,17'd8780,17'd8780,17'd29593,17'd29593,17'd29592,17'd9933,17'd6219,17'd28185,17'd28185,17'd31717,17'd9091,17'd27815,17'd27933,17'd27933,17'd28183,17'd28183,17'd31551,17'd27933,17'd29592,17'd27815,17'd9934,17'd7011,17'd8630,17'd9093,17'd8783,17'd6858,17'd34659,17'd10782,17'd8161,17'd34660,17'd34661,17'd34662,17'd34663,17'd1938,17'd34664,17'd34665,17'd622,17'd190,17'd192,17'd413,17'd15233,17'd15233,17'd34000,17'd28916,17'd33050,17'd5030,17'd11336,17'd11336,17'd11061,17'd11882,17'd33051,17'd33051,17'd31729,17'd31101,17'd29170,17'd29170,17'd31409,17'd31409,17'd31900,17'd29039,17'd27710,17'd28545,17'd29610,17'd29037,17'd27094,17'd15233,17'd2393,17'd12026,17'd11337,17'd1396,17'd608,17'd34666,17'd440,17'd31730,17'd34667,17'd34668
},
'{
17'd4890,17'd4890,17'd4890,17'd29756,17'd4892,17'd14743,17'd7545,17'd4886,17'd10535,17'd3252,17'd3101,17'd3428,17'd3428,17'd3101,17'd2422,17'd1688,17'd2597,17'd2425,17'd1416,17'd26344,17'd34669,17'd27,17'd28,17'd287,17'd7061,17'd7728,17'd7388,17'd7556,17'd6439,17'd11211,17'd12507,17'd4742,17'd3597,17'd4433,17'd4259,17'd1978,17'd34167,17'd34670,17'd3109,17'd2952,17'd34514,17'd34671,17'd2444,17'd32091,17'd26608,17'd31736,17'd19371,17'd34672,17'd34174,17'd32892,17'd34673,17'd34356,17'd34674,17'd34521,17'd16029,17'd15384,17'd32739,17'd16034,17'd16289,17'd18774,17'd20423,17'd14764,17'd13599,17'd12678,17'd13462,17'd13462,17'd13209,17'd13093,17'd34675,17'd19756,17'd34676,17'd16523,17'd34677,17'd32572,17'd34525,17'd34678,17'd34679,17'd34680,17'd34681,17'd34682,17'd34683,17'd34367,17'd15913,17'd34684,17'd10291,17'd12070,17'd19521,17'd11920,17'd8702,17'd14640,17'd14231,17'd11095,17'd11095,17'd14231,17'd14640,17'd12686,17'd34685,17'd34686,17'd31750,17'd34687,17'd7597,17'd34688,17'd34689,17'd34690,17'd34691,17'd34537,17'd32432,17'd34692,17'd34693,17'd12116,17'd15688,17'd17839,17'd9479,17'd9480,17'd9478,17'd24037,17'd22814,17'd8729,17'd17609,17'd14932,17'd34694,17'd7952,17'd10339,17'd10337,17'd34695,17'd29782,17'd25280,17'd14259,17'd24031,17'd34696,17'd30675,17'd33567,17'd34544,17'd34697,17'd34545,17'd34037,17'd34698,17'd30074,17'd28462,17'd27121,17'd23515,17'd21671,17'd14261,17'd11522,17'd11399,17'd9883,17'd9620,17'd9743,17'd8874,17'd9038,17'd15944,17'd24361,17'd15944,17'd23859,17'd16562,17'd34699,17'd17729,17'd15684,17'd15180,17'd17011,17'd11277,17'd10479,17'd10326,17'd25675,17'd24211,17'd8571,17'd34700,17'd34701,17'd34702,17'd34703,17'd29328,17'd34704,17'd33095,17'd33728,17'd34553,17'd34209,17'd34705,17'd34556,17'd31288,17'd30974,17'd28229,17'd23855,17'd13517,17'd34706,17'd34707,17'd34708,17'd33248,17'd33579,17'd33416,17'd31140,17'd33412,17'd34709,17'd30090,17'd34710,17'd34711,17'd29940,17'd34712,17'd34218,17'd29496,17'd29496,17'd30253,17'd33257,17'd33890,17'd34713,17'd33892,17'd34566,17'd34714,17'd34568,17'd34715,17'd34716,17'd34717,17'd33599,17'd34718,17'd34719,17'd34720,17'd34721,17'd34722,17'd34723,17'd34724,17'd34725,17'd34726,17'd34727,17'd34728,17'd34729,17'd34730,17'd33920,17'd34731,17'd34731,17'd34731,17'd34731,17'd34732,17'd33768,17'd34733,17'd34734,17'd34593,17'd34592,17'd34735,17'd34593,17'd34429,17'd34079,17'd34736,17'd34737,17'd34738,17'd34739,17'd34257,17'd34740,17'd34741,17'd34742,17'd34743,17'd34744,17'd34745,17'd34746,17'd34093,17'd34442,17'd34607,17'd34747,17'd34748,17'd34749,17'd34750,17'd34751,17'd34271,17'd34098,17'd34101,17'd34752,17'd34753,17'd34754,17'd34755,17'd34756,17'd34104,17'd33790,17'd32994,17'd32496,17'd27260,17'd25566,17'd27882,17'd32007,17'd23920,17'd23215,17'd33315,17'd22157,17'd32501,17'd34757,17'd33481,17'd34758,17'd34617,17'd32997,17'd34759,17'd34620,17'd31495,17'd23388,17'd30733,17'd23561,17'd28008,17'd25179,17'd25435,17'd25707,17'd27027,17'd29245,17'd33001,17'd32192,17'd32507,17'd32193,17'd33654,17'd32355,17'd28728,17'd29536,17'd29981,17'd31037,17'd31838,17'd34286,17'd32508,17'd30435,17'd34760,17'd34761,17'd34290,17'd30887,17'd33326,17'd34762,17'd28990,17'd32692,17'd32042,17'd34763,17'd34764,17'd34765,17'd25034,17'd24421,17'd29689,17'd34766,17'd24418,17'd24893,17'd23724,17'd24583,17'd25312,17'd34767,17'd34768,17'd34769,17'd34770,17'd34771,17'd27664,17'd26913,17'd32207,17'd28505,17'd29261,17'd27391,17'd28617,17'd28276,17'd34473,17'd34772,17'd25964,17'd34773,17'd34463,17'd34774,17'd29256,17'd28597,17'd23723,17'd26285,17'd25560,17'd25559,17'd28724,17'd32364,17'd28600,17'd24898,17'd26396,17'd22859,17'd34775,17'd34776,17'd34777,17'd34778,17'd34779,17'd34780,17'd34781,17'd34782,17'd34783,17'd34784,17'd23084,17'd22397,17'd31883,17'd34785,17'd34786,17'd34651,17'd34787,17'd34788,17'd34789,17'd34790,17'd4525,17'd5157,17'd4846,17'd34791,17'd4683,17'd33692,17'd6392,17'd13800,17'd34792,17'd30933,17'd27933,17'd28184,17'd30487,17'd28058,17'd32074,17'd31243,17'd34793,17'd31551,17'd10515,17'd28184,17'd28058,17'd7668,17'd9933,17'd29593,17'd29592,17'd9933,17'd9091,17'd31717,17'd28185,17'd30638,17'd6390,17'd8780,17'd10515,17'd27933,17'd28183,17'd28183,17'd31551,17'd30933,17'd29592,17'd29592,17'd9934,17'd7011,17'd8630,17'd9093,17'd34794,17'd8938,17'd34795,17'd34796,17'd8310,17'd34660,17'd34797,17'd34798,17'd34799,17'd34800,17'd34801,17'd34665,17'd244,17'd410,17'd411,17'd602,17'd1383,17'd2394,17'd34000,17'd28916,17'd34001,17'd5777,17'd11336,17'd11336,17'd11061,17'd11882,17'd33051,17'd33051,17'd31729,17'd31101,17'd29170,17'd29170,17'd31409,17'd31409,17'd31900,17'd31900,17'd29039,17'd30649,17'd27708,17'd27707,17'd28916,17'd15233,17'd2393,17'd12026,17'd5371,17'd1262,17'd609,17'd34666,17'd440,17'd585,17'd34511,17'd34668
},
'{
17'd5200,17'd4890,17'd4890,17'd29756,17'd4892,17'd4246,17'd7545,17'd4886,17'd10535,17'd3252,17'd3101,17'd3428,17'd3428,17'd3101,17'd2422,17'd1688,17'd2597,17'd2425,17'd1416,17'd26344,17'd34669,17'd27,17'd28,17'd2424,17'd7061,17'd7728,17'd7388,17'd7226,17'd6440,17'd27445,17'd13067,17'd4581,17'd3597,17'd4583,17'd2786,17'd1978,17'd34167,17'd34802,17'd3109,17'd2952,17'd34008,17'd34671,17'd2444,17'd34803,17'd33697,17'd4593,17'd15371,17'd31913,17'd34804,17'd34805,17'd34806,17'd34807,17'd34674,17'd34177,17'd15767,17'd15641,17'd14767,17'd17445,17'd16986,17'd19382,17'd22630,17'd14621,17'd13599,17'd12678,17'd13968,17'd14344,17'd16284,17'd13093,17'd34181,17'd19261,17'd34808,17'd31575,17'd34183,17'd34809,17'd33553,17'd34810,17'd34811,17'd34812,17'd34813,17'd34814,17'd34367,17'd33228,17'd16293,17'd34815,17'd10125,17'd12070,17'd19521,17'd12071,17'd8702,17'd14640,17'd14231,17'd9165,17'd9165,17'd13611,17'd14359,17'd12686,17'd34816,17'd34686,17'd34817,17'd34687,17'd7597,17'd34818,17'd34819,17'd34820,17'd34821,17'd34822,17'd34823,17'd34824,17'd27983,17'd16796,17'd10164,17'd9740,17'd10026,17'd10026,17'd9478,17'd9478,17'd16795,17'd11966,17'd8253,17'd7789,17'd34694,17'd34825,17'd9887,17'd16440,17'd26875,17'd34826,17'd23337,17'd24363,17'd26371,17'd30673,17'd34827,17'd33719,17'd34828,17'd34697,17'd34545,17'd31288,17'd34698,17'd29930,17'd28818,17'd28107,17'd23515,17'd21671,17'd13646,17'd11274,17'd19532,17'd10024,17'd9340,17'd9189,17'd15684,17'd9039,17'd15944,17'd24361,17'd9039,17'd9045,17'd10177,17'd30217,17'd11966,17'd29920,17'd24361,17'd16549,17'd12116,17'd9883,17'd10741,17'd25675,17'd24040,17'd8247,17'd34829,17'd34830,17'd34831,17'd34832,17'd29779,17'd33096,17'd34833,17'd33729,17'd34834,17'd34834,17'd34556,17'd31590,17'd34835,17'd29482,17'd27234,17'd12415,17'd13518,17'd34836,17'd34837,17'd34215,17'd33579,17'd33736,17'd31140,17'd34393,17'd30380,17'd34049,17'd34838,17'd34710,17'd10322,17'd34712,17'd34218,17'd30552,17'd30705,17'd30859,17'd34839,17'd31309,17'd30855,17'd34840,17'd34565,17'd34714,17'd34568,17'd31152,17'd31164,17'd34841,17'd34842,17'd34843,17'd34844,17'd34845,17'd34846,17'd34847,17'd34848,17'd34849,17'd34850,17'd34851,17'd34852,17'd34853,17'd34854,17'd34855,17'd34856,17'd34731,17'd34857,17'd34425,17'd34247,17'd34428,17'd34425,17'd34080,17'd34425,17'd34858,17'd34247,17'd34593,17'd34735,17'd34593,17'd34247,17'd34594,17'd34594,17'd34859,17'd34860,17'd34861,17'd34862,17'd34863,17'd34864,17'd34865,17'd34866,17'd34867,17'd34868,17'd34869,17'd34870,17'd34871,17'd34442,17'd34267,17'd34872,17'd33936,17'd33783,17'd34873,17'd33470,17'd34271,17'd34874,17'd34101,17'd34875,17'd34613,17'd34449,17'd34876,17'd34877,17'd34104,17'd33790,17'd32185,17'd33478,17'd28253,17'd25317,17'd32007,17'd24087,17'd30128,17'd22327,17'd22159,17'd22009,17'd34878,17'd34879,17'd34880,17'd34881,17'd31660,17'd34882,17'd34620,17'd31495,17'd23569,17'd34883,17'd34884,17'd28129,17'd32007,17'd28484,17'd25708,17'd28853,17'd31035,17'd29977,17'd32354,17'd32017,17'd32017,17'd33654,17'd32355,17'd28372,17'd29537,17'd29833,17'd31037,17'd33167,17'd32508,17'd34114,17'd30435,17'd34760,17'd34761,17'd34885,17'd30887,17'd34886,17'd34887,17'd30753,17'd34888,17'd34889,17'd34890,17'd34891,17'd34892,17'd34893,17'd34894,17'd34895,17'd23563,17'd24418,17'd24894,17'd25173,17'd24242,17'd25948,17'd25945,17'd28727,17'd34896,17'd34897,17'd30290,17'd27535,17'd28623,17'd29555,17'd31517,17'd34898,17'd34899,17'd30450,17'd25458,17'd25199,17'd34900,17'd25333,17'd34901,17'd34902,17'd34903,17'd34904,17'd25835,17'd25567,17'd24408,17'd25699,17'd26055,17'd27372,17'd26174,17'd28723,17'd25320,17'd23919,17'd30425,17'd34905,17'd34906,17'd34907,17'd24596,17'd34908,17'd34909,17'd34910,17'd34911,17'd34912,17'd34913,17'd34914,17'd34915,17'd31712,17'd4984,17'd34916,17'd34917,17'd34918,17'd4666,17'd34919,17'd34920,17'd4836,17'd34921,17'd27697,17'd4846,17'd4687,17'd5330,17'd6392,17'd12307,17'd34922,17'd30933,17'd27933,17'd27815,17'd28058,17'd28058,17'd27696,17'd29593,17'd30933,17'd31551,17'd10642,17'd28184,17'd6391,17'd7499,17'd27696,17'd29592,17'd29592,17'd9933,17'd7499,17'd6554,17'd28185,17'd30638,17'd6554,17'd7668,17'd10515,17'd27933,17'd31551,17'd31551,17'd31551,17'd31551,17'd27933,17'd27815,17'd7500,17'd7011,17'd8630,17'd34923,17'd34794,17'd34924,17'd34659,17'd34796,17'd34925,17'd4699,17'd34926,17'd34927,17'd34928,17'd24664,17'd34929,17'd34930,17'd784,17'd1678,17'd1243,17'd2740,17'd14178,17'd5631,17'd34000,17'd29169,17'd34001,17'd5777,17'd11335,17'd11335,17'd11336,17'd11061,17'd33051,17'd33051,17'd31729,17'd31101,17'd29170,17'd29170,17'd31409,17'd31409,17'd31900,17'd29039,17'd30649,17'd28545,17'd29610,17'd29037,17'd27094,17'd15233,17'd2393,17'd6868,17'd5957,17'd1396,17'd608,17'd1091,17'd18515,17'd31103,17'd34931,17'd34668
},
'{
17'd4890,17'd4890,17'd4890,17'd29756,17'd4892,17'd4246,17'd7711,17'd4886,17'd10535,17'd3252,17'd3101,17'd3428,17'd3428,17'd3101,17'd2422,17'd1688,17'd2597,17'd2425,17'd1416,17'd4089,17'd1278,17'd27,17'd28,17'd2424,17'd7061,17'd7728,17'd7388,17'd6599,17'd27592,17'd27445,17'd13067,17'd4432,17'd3597,17'd4583,17'd2786,17'd1978,17'd34167,17'd34347,17'd3109,17'd2952,17'd34008,17'd34932,17'd29177,17'd22617,17'd26242,17'd34933,17'd34934,17'd32095,17'd34935,17'd34519,17'd34807,17'd34936,17'd34937,17'd34177,17'd15767,17'd15384,17'd14768,17'd17320,17'd16986,17'd19006,17'd16658,17'd13211,17'd12954,17'd12678,17'd13968,17'd12357,17'd12679,17'd34938,17'd34939,17'd34940,17'd18298,17'd34941,17'd34942,17'd34943,17'd34944,17'd33066,17'd34364,17'd34945,17'd34946,17'd34814,17'd34367,17'd33864,17'd16778,17'd18667,17'd10291,17'd9310,17'd12370,17'd12071,17'd12371,17'd14640,17'd14231,17'd13611,17'd13611,17'd14231,17'd14640,17'd12686,17'd34816,17'd34368,17'd8391,17'd34947,17'd34948,17'd34949,17'd34950,17'd34951,17'd34952,17'd34822,17'd34953,17'd34954,17'd33876,17'd9884,17'd10479,17'd16796,17'd22812,17'd22812,17'd16554,17'd9478,17'd14811,17'd24712,17'd34040,17'd7954,17'd34955,17'd9350,17'd24545,17'd26631,17'd27744,17'd34956,17'd23337,17'd29488,17'd31443,17'd30370,17'd30833,17'd34957,17'd34828,17'd34697,17'd31590,17'd31288,17'd31767,17'd29067,17'd30222,17'd25672,17'd23515,17'd24995,17'd15185,17'd10854,17'd26152,17'd10992,17'd23679,17'd9190,17'd10336,17'd17123,17'd15944,17'd17123,17'd9194,17'd10338,17'd18201,17'd12587,17'd8572,17'd29920,17'd24361,17'd16549,17'd12116,17'd11671,17'd9739,17'd15048,17'd9194,17'd34958,17'd34959,17'd34960,17'd34961,17'd34962,17'd31295,17'd32932,17'd32930,17'd33728,17'd34963,17'd34964,17'd31590,17'd34037,17'd30677,17'd34390,17'd16556,17'd14525,17'd21506,17'd34965,17'd34215,17'd30236,17'd33582,17'd34966,17'd34393,17'd34967,17'd34968,17'd32610,17'd34969,17'd34710,17'd11272,17'd34970,17'd29496,17'd34971,17'd34972,17'd31000,17'd32305,17'd30699,17'd34973,17'd34565,17'd34714,17'd34974,17'd34975,17'd34976,17'd34977,17'd34978,17'd34979,17'd34980,17'd34981,17'd34982,17'd34983,17'd34984,17'd34985,17'd34986,17'd34987,17'd34988,17'd34989,17'd34990,17'd34991,17'd34992,17'd34586,17'd34993,17'd34080,17'd34425,17'd34428,17'd34735,17'd34593,17'd34247,17'd34428,17'd34428,17'd34428,17'd34428,17'd34247,17'd34735,17'd34735,17'd34592,17'd34592,17'd34247,17'd34994,17'd34995,17'd34996,17'd34997,17'd34998,17'd34999,17'd35000,17'd35001,17'd35002,17'd35003,17'd35004,17'd35005,17'd35006,17'd34747,17'd35007,17'd34748,17'd34096,17'd34610,17'd34097,17'd33470,17'd34874,17'd35008,17'd35009,17'd34754,17'd35010,17'd35010,17'd34450,17'd34451,17'd33790,17'd35011,17'd32006,17'd35012,17'd28600,17'd25180,17'd30431,17'd23387,17'd22502,17'd22681,17'd23222,17'd35013,17'd33947,17'd35014,17'd35015,17'd33648,17'd35016,17'd35017,17'd35018,17'd33158,17'd30424,17'd28975,17'd23563,17'd24895,17'd28369,17'd27766,17'd28978,17'd28486,17'd29379,17'd32354,17'd32017,17'd33654,17'd33654,17'd32355,17'd28372,17'd28857,17'd32508,17'd31037,17'd33167,17'd34286,17'd32508,17'd30435,17'd34760,17'd34761,17'd34885,17'd30743,17'd34886,17'd34887,17'd30753,17'd34888,17'd32042,17'd34763,17'd34764,17'd35019,17'd35020,17'd24421,17'd35021,17'd35022,17'd24252,17'd24894,17'd25173,17'd24584,17'd25561,17'd35023,17'd35024,17'd35025,17'd35026,17'd35027,17'd27152,17'd35028,17'd35029,17'd31517,17'd31517,17'd34899,17'd27661,17'd26411,17'd25199,17'd35030,17'd35031,17'd35032,17'd35033,17'd34635,17'd33017,17'd35034,17'd35035,17'd25708,17'd25699,17'd25696,17'd35011,17'd27259,17'd27766,17'd28850,17'd35036,17'd23217,17'd35037,17'd35038,17'd23744,17'd35039,17'd35040,17'd35041,17'd35042,17'd35043,17'd35044,17'd35045,17'd35046,17'd35047,17'd17250,17'd8286,17'd33530,17'd3829,17'd5140,17'd35048,17'd35049,17'd33531,17'd34156,17'd27697,17'd35050,17'd27697,17'd29739,17'd5333,17'd25084,17'd14050,17'd35051,17'd31715,17'd30933,17'd10515,17'd28058,17'd28058,17'd9933,17'd35052,17'd30933,17'd30933,17'd10642,17'd28184,17'd7499,17'd32073,17'd29740,17'd29592,17'd29592,17'd27815,17'd7499,17'd6390,17'd28185,17'd30333,17'd31891,17'd9091,17'd27815,17'd27933,17'd31551,17'd31551,17'd31551,17'd31551,17'd27933,17'd29592,17'd9934,17'd7011,17'd34336,17'd34923,17'd6396,17'd8938,17'd34795,17'd35053,17'd34925,17'd35054,17'd35055,17'd35056,17'd35057,17'd34342,17'd34929,17'd35058,17'd35059,17'd627,17'd954,17'd6407,17'd5940,17'd14586,17'd35060,17'd28916,17'd34001,17'd5777,17'd11335,17'd11335,17'd11336,17'd11061,17'd33051,17'd33051,17'd31729,17'd31101,17'd29170,17'd29170,17'd31409,17'd31409,17'd31900,17'd31900,17'd29039,17'd35061,17'd28315,17'd32082,17'd28916,17'd15233,17'd2393,17'd12026,17'd5371,17'd1262,17'd609,17'd1091,17'd18515,17'd218,17'd35062,17'd34668
},
'{
17'd4890,17'd4890,17'd32728,17'd35063,17'd4892,17'd4246,17'd7711,17'd7214,17'd3252,17'd3252,17'd3101,17'd3428,17'd3428,17'd3101,17'd2422,17'd1688,17'd2596,17'd2425,17'd1416,17'd4089,17'd1278,17'd27,17'd28,17'd2424,17'd7061,17'd7556,17'd6600,17'd6599,17'd26971,17'd6110,17'd5055,17'd4253,17'd3261,17'd24967,17'd2786,17'd3917,17'd33851,17'd32254,17'd24181,17'd32255,17'd34008,17'd34932,17'd35064,17'd27717,17'd26132,17'd35065,17'd26134,17'd35066,17'd35067,17'd34673,17'd34807,17'd34936,17'd31917,17'd16029,17'd15641,17'd14767,17'd16033,17'd17319,17'd18774,17'd12681,17'd12361,17'd13211,17'd12954,17'd13092,17'd13968,17'd13597,17'd13209,17'd34180,17'd35068,17'd18536,17'd35069,17'd35070,17'd15265,17'd34943,17'd33554,17'd33555,17'd35071,17'd35072,17'd35073,17'd34814,17'd34367,17'd35074,17'd14781,17'd9992,17'd35075,17'd11239,17'd19521,17'd12685,17'd12371,17'd14640,17'd14231,17'd14231,17'd14231,17'd14231,17'd14640,17'd25261,17'd35076,17'd35077,17'd35078,17'd35079,17'd35080,17'd35081,17'd35082,17'd35083,17'd35084,17'd35085,17'd35086,17'd35087,17'd18325,17'd11671,17'd12863,17'd10169,17'd35088,17'd9743,17'd15187,17'd18080,17'd23859,17'd9744,17'd35089,17'd35090,17'd35091,17'd14527,17'd12425,17'd16552,17'd17606,17'd20046,17'd13367,17'd24362,17'd26873,17'd29924,17'd32919,17'd35092,17'd35093,17'd34697,17'd31590,17'd31288,17'd33884,17'd28461,17'd28103,17'd24537,17'd22819,17'd14261,17'd13762,17'd14263,17'd21503,17'd10857,17'd9191,17'd9190,17'd17480,17'd16795,17'd17123,17'd15684,17'd17237,17'd32921,17'd35094,17'd12867,17'd8572,17'd23861,17'd24361,17'd11809,17'd9885,17'd11277,17'd15048,17'd9345,17'd9621,17'd35095,17'd35096,17'd35097,17'd35098,17'd28692,17'd35099,17'd32770,17'd34387,17'd34046,17'd35100,17'd34545,17'd34037,17'd33576,17'd29330,17'd35101,17'd21504,17'd13760,17'd29653,17'd33737,17'd31450,17'd35102,17'd31954,17'd34966,17'd35103,17'd35104,17'd35105,17'd35106,17'd10598,17'd10321,17'd29810,17'd29496,17'd29799,17'd35107,17'd30542,17'd30096,17'd35108,17'd35109,17'd35110,17'd34565,17'd35111,17'd31152,17'd35112,17'd35113,17'd35114,17'd35115,17'd35116,17'd35117,17'd35118,17'd35119,17'd35120,17'd35121,17'd35122,17'd35123,17'd35124,17'd35125,17'd35126,17'd35127,17'd35128,17'd35129,17'd35130,17'd35131,17'd34254,17'd34425,17'd34858,17'd34247,17'd34735,17'd34735,17'd34593,17'd34593,17'd34247,17'd34247,17'd34593,17'd35132,17'd35133,17'd35134,17'd35135,17'd35136,17'd34076,17'd35137,17'd35138,17'd35139,17'd35140,17'd35141,17'd35142,17'd35143,17'd35144,17'd35145,17'd35146,17'd35147,17'd35006,17'd34608,17'd33634,17'd34748,17'd34096,17'd34610,17'd33784,17'd34097,17'd35148,17'd34101,17'd34875,17'd34613,17'd34754,17'd35149,17'd35150,17'd35151,17'd35152,17'd34637,17'd31827,17'd28252,17'd28723,17'd25178,17'd32659,17'd29376,17'd33158,17'd33311,17'd35153,17'd22003,17'd33947,17'd35154,17'd35155,17'd35156,17'd35157,17'd35158,17'd22858,17'd22502,17'd30578,17'd28975,17'd29243,17'd35159,17'd29244,17'd28720,17'd28252,17'd27027,17'd29246,17'd30279,17'd28373,17'd28134,17'd28134,17'd32355,17'd28372,17'd28728,17'd34114,17'd31037,17'd33167,17'd32508,17'd29831,17'd29381,17'd34760,17'd34761,17'd34885,17'd30887,17'd34886,17'd35160,17'd35161,17'd35162,17'd32042,17'd35163,17'd34628,17'd35164,17'd35165,17'd34894,17'd35166,17'd23563,17'd24418,17'd33340,17'd27882,17'd28602,17'd25172,17'd27145,17'd28979,17'd34468,17'd35167,17'd35168,17'd32838,17'd35169,17'd35170,17'd34471,17'd32519,17'd31848,17'd27904,17'd25731,17'd25845,17'd35171,17'd35172,17'd23060,17'd23060,17'd35173,17'd35174,17'd30595,17'd31855,17'd32364,17'd28853,17'd25696,17'd26525,17'd25429,17'd25949,17'd25317,17'd30126,17'd23923,17'd35175,17'd35176,17'd35177,17'd35178,17'd35179,17'd35180,17'd35181,17'd35182,17'd35183,17'd35184,17'd20224,17'd35185,17'd35186,17'd35187,17'd35188,17'd35048,17'd5140,17'd35189,17'd35190,17'd4987,17'd35191,17'd35192,17'd35193,17'd35193,17'd30794,17'd26828,17'd35194,17'd12468,17'd35195,17'd35196,17'd28057,17'd10642,17'd8780,17'd8780,17'd27815,17'd35052,17'd31243,17'd30933,17'd10642,17'd10514,17'd7499,17'd32073,17'd32074,17'd9933,17'd9933,17'd27815,17'd7668,17'd6219,17'd27935,17'd30333,17'd33369,17'd32073,17'd9933,17'd10515,17'd28183,17'd28183,17'd31551,17'd31551,17'd30933,17'd29592,17'd9934,17'd6223,17'd35197,17'd35198,17'd6396,17'd5341,17'd6859,17'd6860,17'd35199,17'd35200,17'd35201,17'd35202,17'd35203,17'd35204,17'd35205,17'd35206,17'd24496,17'd226,17'd607,17'd1667,17'd5630,17'd14586,17'd35060,17'd5030,17'd34001,17'd5631,17'd11335,17'd11335,17'd7537,17'd7705,17'd34002,17'd34002,17'd27949,17'd35207,17'd31251,17'd31251,17'd31409,17'd31409,17'd31900,17'd31900,17'd29039,17'd27708,17'd27707,17'd29169,17'd5777,17'd14586,17'd2393,17'd6868,17'd5957,17'd1396,17'd1539,17'd430,17'd35208,17'd218,17'd35062,17'd35209
},
'{
17'd4890,17'd5200,17'd32728,17'd35063,17'd4243,17'd4246,17'd7711,17'd7214,17'd3252,17'd2935,17'd2934,17'd3428,17'd3428,17'd3101,17'd2422,17'd1688,17'd2596,17'd2257,17'd1416,17'd4089,17'd1278,17'd27,17'd28,17'd2424,17'd7061,17'd7556,17'd6600,17'd6599,17'd26971,17'd12931,17'd5055,17'd4253,17'd2608,17'd24967,17'd2786,17'd1978,17'd34167,17'd34347,17'd1147,17'd32255,17'd33544,17'd34932,17'd2445,17'd22112,17'd21029,17'd18524,17'd35210,17'd15753,17'd35211,17'd34520,17'd34936,17'd34937,17'd31918,17'd16029,17'd15641,17'd14767,17'd15902,17'd17319,17'd17689,17'd16658,17'd14470,17'd13093,17'd13092,17'd13092,17'd13968,17'd13092,17'd12813,17'd9836,17'd35212,17'd21040,17'd35213,17'd34942,17'd32572,17'd33065,17'd33703,17'd34187,17'd35214,17'd35215,17'd34814,17'd35216,17'd33228,17'd35217,17'd14358,17'd9992,17'd12070,17'd11095,17'd12685,17'd14640,17'd35218,17'd12371,17'd12685,17'd14231,17'd14231,17'd14640,17'd7264,17'd35219,17'd35076,17'd35220,17'd35221,17'd34532,17'd35222,17'd35223,17'd35224,17'd35225,17'd35226,17'd35227,17'd10147,17'd35228,17'd18196,17'd11671,17'd11527,17'd10169,17'd35088,17'd22813,17'd15187,17'd18080,17'd29637,17'd24213,17'd35229,17'd35090,17'd7952,17'd8250,17'd16205,17'd17728,17'd33725,17'd35230,17'd14382,17'd26496,17'd29197,17'd31940,17'd34543,17'd35092,17'd35093,17'd31589,17'd34037,17'd33568,17'd30972,17'd28571,17'd28816,17'd24537,17'd24362,17'd14259,17'd11397,17'd24996,17'd10992,17'd9346,17'd9190,17'd9190,17'd17480,17'd16795,17'd23859,17'd8886,17'd14675,17'd12725,17'd33715,17'd8248,17'd8573,17'd23861,17'd24361,17'd9345,17'd9341,17'd15048,17'd23857,17'd8874,17'd24367,17'd35231,17'd35232,17'd35233,17'd35234,17'd35235,17'd35236,17'd35237,17'd35238,17'd34044,17'd35239,17'd31589,17'd33576,17'd31129,17'd28571,17'd35240,17'd14525,17'd29339,17'd31777,17'd31140,17'd35102,17'd31954,17'd34966,17'd35103,17'd35241,17'd35242,17'd35243,17'd35244,17'd35245,17'd31283,17'd29658,17'd29349,17'd29799,17'd30542,17'd30096,17'd35246,17'd31154,17'd35247,17'd35248,17'd33894,17'd31152,17'd35249,17'd35250,17'd35251,17'd35115,17'd35252,17'd35253,17'd35254,17'd35255,17'd35256,17'd35257,17'd35258,17'd35259,17'd35260,17'd35261,17'd35262,17'd35263,17'd35264,17'd35265,17'd35266,17'd35267,17'd35268,17'd34254,17'd34247,17'd34592,17'd34735,17'd34593,17'd34735,17'd34592,17'd34592,17'd35132,17'd35132,17'd35132,17'd35136,17'd35269,17'd35270,17'd35271,17'd35272,17'd35273,17'd35274,17'd35275,17'd35276,17'd35277,17'd35278,17'd35279,17'd35280,17'd35281,17'd35282,17'd35283,17'd35284,17'd35006,17'd34747,17'd35285,17'd34748,17'd34444,17'd34096,17'd33784,17'd34097,17'd35286,17'd34874,17'd34875,17'd35287,17'd35288,17'd35149,17'd35289,17'd35290,17'd35291,17'd30735,17'd27146,17'd26903,17'd27766,17'd25438,17'd28851,17'd23918,17'd29829,17'd22500,17'd35292,17'd22336,17'd33647,17'd35293,17'd35294,17'd35295,17'd23394,17'd33645,17'd35296,17'd22502,17'd33801,17'd28722,17'd23564,17'd32659,17'd25178,17'd28130,17'd25707,17'd27258,17'd29245,17'd30279,17'd28373,17'd28134,17'd28134,17'd32355,17'd28372,17'd28728,17'd34114,17'd29981,17'd33167,17'd32833,17'd29831,17'd29381,17'd35297,17'd34288,17'd33805,17'd35298,17'd35299,17'd35160,17'd35300,17'd35301,17'd32042,17'd34627,17'd35302,17'd35303,17'd33331,17'd24421,17'd23921,17'd35022,17'd24743,17'd33340,17'd25709,17'd26064,17'd25704,17'd35304,17'd35305,17'd34632,17'd35306,17'd29835,17'd35307,17'd35308,17'd28506,17'd35309,17'd35310,17'd31848,17'd32207,17'd25731,17'd25845,17'd25200,17'd35311,17'd35312,17'd35313,17'd35314,17'd35315,17'd35316,17'd35317,17'd35318,17'd28853,17'd25554,17'd25697,17'd25698,17'd27514,17'd28600,17'd32007,17'd23565,17'd30729,17'd35319,17'd35320,17'd35321,17'd24426,17'd35322,17'd35323,17'd35324,17'd35325,17'd35326,17'd20667,17'd35327,17'd35328,17'd35329,17'd35188,17'd35189,17'd35330,17'd35330,17'd35331,17'd35332,17'd35333,17'd35334,17'd35335,17'd35336,17'd35337,17'd30935,17'd25361,17'd14050,17'd35338,17'd35339,17'd35340,17'd11037,17'd28184,17'd8780,17'd27815,17'd35052,17'd31243,17'd31243,17'd28183,17'd10515,17'd7668,17'd32073,17'd32074,17'd27696,17'd27696,17'd28184,17'd28058,17'd6219,17'd27935,17'd30333,17'd33369,17'd6554,17'd7668,17'd27815,17'd28183,17'd28183,17'd31551,17'd29158,17'd30933,17'd29593,17'd9934,17'd7011,17'd34336,17'd35198,17'd6070,17'd5341,17'd6859,17'd6860,17'd35199,17'd6714,17'd35341,17'd35342,17'd35343,17'd35344,17'd35345,17'd35346,17'd1665,17'd8014,17'd233,17'd1262,17'd4729,17'd9123,17'd35060,17'd28657,17'd5777,17'd5631,17'd11335,17'd5029,17'd8507,17'd7705,17'd34002,17'd34002,17'd33051,17'd27949,17'd31251,17'd31251,17'd31409,17'd31409,17'd31900,17'd31900,17'd29039,17'd29441,17'd28315,17'd32082,17'd5030,17'd14586,17'd2393,17'd12026,17'd5371,17'd1262,17'd428,17'd430,17'd35208,17'd218,17'd35347,17'd35209
},
'{
17'd29756,17'd29756,17'd32728,17'd35063,17'd4892,17'd4887,17'd3250,17'd1831,17'd3252,17'd2935,17'd2934,17'd3592,17'd3428,17'd3101,17'd2422,17'd1688,17'd2596,17'd2257,17'd1416,17'd4089,17'd1278,17'd27,17'd6744,17'd9275,17'd7225,17'd7556,17'd6600,17'd6599,17'd26971,17'd12931,17'd4742,17'd3911,17'd2608,17'd24967,17'd2786,17'd33850,17'd33851,17'd3437,17'd1147,17'd32255,17'd33544,17'd34932,17'd27957,17'd14197,17'd3930,17'd18398,17'd35348,17'd35349,17'd35350,17'd35351,17'd34936,17'd34177,17'd33548,17'd16029,17'd14892,17'd16881,17'd24348,17'd17206,17'd19006,17'd12361,17'd13211,17'd12954,17'd15762,17'd13462,17'd14469,17'd13092,17'd35352,17'd34939,17'd35353,17'd35354,17'd16292,17'd32741,17'd35355,17'd33224,17'd34810,17'd34187,17'd35356,17'd35357,17'd34683,17'd35358,17'd15535,17'd16778,17'd35359,17'd9849,17'd9310,17'd18542,17'd12685,17'd8702,17'd35218,17'd14640,17'd14231,17'd14231,17'd14359,17'd14640,17'd7264,17'd7104,17'd8549,17'd35360,17'd35361,17'd35362,17'd35363,17'd35364,17'd35365,17'd35366,17'd35367,17'd35368,17'd35369,17'd35370,17'd9618,17'd11671,17'd19155,17'd10333,17'd16682,17'd10175,17'd9345,17'd17716,17'd29920,17'd14812,17'd35229,17'd35371,17'd16566,17'd25679,17'd25677,17'd10334,17'd19779,17'd13368,17'd29783,17'd24208,17'd28343,17'd34827,17'd30834,17'd31442,17'd31590,17'd31590,17'd34380,17'd34381,17'd31587,17'd35372,17'd26370,17'd24707,17'd15055,17'd14264,17'd11275,17'd10328,17'd9341,17'd9339,17'd9190,17'd9190,17'd26153,17'd14811,17'd16317,17'd24368,17'd18808,17'd13005,17'd13005,17'd8249,17'd8573,17'd23861,17'd15944,17'd9346,17'd9341,17'd15048,17'd25525,17'd9044,17'd24367,17'd16439,17'd35373,17'd35374,17'd32286,17'd32596,17'd35375,17'd32929,17'd34211,17'd34044,17'd35239,17'd31943,17'd31588,17'd31940,17'd35376,17'd16556,17'd14525,17'd29490,17'd31140,17'd35102,17'd35102,17'd34966,17'd35103,17'd35377,17'd34561,17'd30090,17'd35378,17'd10468,17'd30093,17'd29810,17'd29496,17'd34972,17'd30542,17'd35379,17'd35246,17'd30395,17'd35380,17'd33893,17'd35381,17'd35382,17'd35383,17'd34977,17'd35384,17'd35385,17'd35386,17'd35387,17'd35388,17'd35389,17'd35390,17'd35391,17'd35392,17'd35393,17'd35394,17'd35395,17'd35396,17'd35397,17'd35398,17'd35399,17'd35400,17'd35267,17'd35401,17'd35401,17'd34253,17'd34858,17'd34247,17'd34428,17'd34428,17'd34593,17'd34592,17'd35132,17'd35402,17'd35402,17'd35403,17'd35403,17'd35404,17'd35270,17'd35405,17'd35271,17'd35406,17'd35407,17'd35408,17'd35409,17'd35410,17'd35411,17'd35412,17'd35413,17'd35414,17'd35415,17'd35416,17'd35417,17'd35418,17'd35419,17'd35420,17'd35007,17'd34444,17'd34096,17'd35421,17'd33784,17'd35422,17'd35148,17'd34752,17'd35009,17'd35423,17'd35149,17'd35424,17'd35424,17'd35425,17'd35426,17'd30586,17'd26903,17'd25565,17'd28369,17'd25032,17'd24086,17'd23736,17'd22502,17'd22334,17'd22005,17'd35427,17'd35428,17'd35294,17'd32499,17'd33480,17'd33944,17'd35429,17'd22503,17'd35430,17'd24902,17'd23564,17'd29534,17'd25030,17'd25317,17'd25565,17'd28853,17'd28727,17'd30279,17'd28373,17'd28134,17'd28134,17'd33485,17'd28371,17'd28728,17'd34114,17'd29833,17'd29979,17'd29690,17'd29536,17'd29381,17'd35431,17'd34288,17'd35432,17'd30284,17'd29696,17'd35433,17'd30893,17'd35434,17'd35435,17'd34627,17'd35302,17'd35436,17'd35437,17'd31350,17'd35438,17'd35439,17'd24743,17'd25180,17'd25709,17'd30606,17'd24735,17'd35440,17'd34767,17'd35441,17'd35442,17'd35443,17'd35444,17'd31508,17'd35445,17'd35446,17'd27162,17'd25967,17'd27904,17'd28024,17'd35447,17'd35448,17'd35449,17'd22703,17'd35450,17'd35451,17'd35452,17'd34293,17'd35161,17'd35453,17'd34311,17'd25696,17'd35454,17'd24578,17'd25561,17'd23554,17'd25320,17'd23731,17'd35455,17'd32503,17'd35456,17'd35457,17'd24425,17'd35458,17'd35459,17'd35460,17'd35325,17'd35461,17'd35462,17'd35463,17'd35464,17'd35465,17'd9499,17'd35330,17'd35466,17'd35467,17'd35468,17'd7654,17'd35469,17'd35470,17'd35471,17'd35472,17'd35473,17'd35474,17'd35475,17'd12468,17'd35476,17'd35477,17'd35478,17'd11316,17'd30332,17'd8780,17'd27815,17'd31888,17'd31243,17'd29592,17'd10515,17'd10642,17'd8780,17'd32073,17'd32073,17'd7499,17'd7668,17'd8780,17'd28058,17'd6220,17'd5614,17'd30333,17'd30333,17'd6554,17'd7499,17'd27815,17'd28183,17'd27933,17'd31551,17'd29158,17'd31551,17'd29593,17'd9934,17'd6223,17'd35197,17'd35479,17'd35480,17'd5923,17'd5485,17'd35481,17'd6073,17'd6399,17'd35482,17'd35483,17'd35484,17'd35485,17'd35486,17'd1807,17'd1809,17'd30342,17'd210,17'd953,17'd4085,17'd9123,17'd35060,17'd5030,17'd2906,17'd5183,17'd9123,17'd9123,17'd8507,17'd7537,17'd9124,17'd34002,17'd33051,17'd35487,17'd31101,17'd31251,17'd31101,17'd31101,17'd31900,17'd31900,17'd29039,17'd27708,17'd27949,17'd33050,17'd5777,17'd14586,17'd12496,17'd6868,17'd5957,17'd1396,17'd1539,17'd430,17'd35208,17'd218,17'd35347,17'd34345
},
'{
17'd10533,17'd10533,17'd29756,17'd35063,17'd4892,17'd4887,17'd2781,17'd1831,17'd3252,17'd2935,17'd2934,17'd3592,17'd3428,17'd3101,17'd2422,17'd1688,17'd2596,17'd2257,17'd17,17'd4089,17'd1278,17'd27,17'd6744,17'd9275,17'd7225,17'd7556,17'd6600,17'd6599,17'd26971,17'd12931,17'd4742,17'd3911,17'd2608,17'd35488,17'd2786,17'd33850,17'd33851,17'd3437,17'd1147,17'd32255,17'd34008,17'd29177,17'd15749,17'd2627,17'd31736,17'd35489,17'd35490,17'd35491,17'd35492,17'd34937,17'd34937,17'd34177,17'd33548,17'd15384,17'd14768,17'd16411,17'd17319,17'd16986,17'd19006,17'd12361,17'd17096,17'd12678,17'd13597,17'd13462,17'd12357,17'd12527,17'd9836,17'd35493,17'd20295,17'd35494,17'd35495,17'd35496,17'd34944,17'd32742,17'd35497,17'd33555,17'd35498,17'd35357,17'd34683,17'd35499,17'd17213,17'd14781,17'd9992,17'd9583,17'd9310,17'd14231,17'd12371,17'd7923,17'd7921,17'd7264,17'd14640,17'd14231,17'd14359,17'd7763,17'd25914,17'd35500,17'd35501,17'd8550,17'd35502,17'd35503,17'd35504,17'd35505,17'd35506,17'd35507,17'd35508,17'd35509,17'd35510,17'd27983,17'd15048,17'd11671,17'd19155,17'd13370,17'd10336,17'd10175,17'd10173,17'd24361,17'd23861,17'd12867,17'd35511,17'd35512,17'd8581,17'd24862,17'd24999,17'd9480,17'd10331,17'd23166,17'd33572,17'd35513,17'd30369,17'd34827,17'd32283,17'd31442,17'd31590,17'd31590,17'd34380,17'd34704,17'd30072,17'd28460,17'd26370,17'd28231,17'd29488,17'd13367,17'd11669,17'd21503,17'd9346,17'd9347,17'd9043,17'd9481,17'd26153,17'd17848,17'd26154,17'd35514,17'd12867,17'd8102,17'd8101,17'd8418,17'd8573,17'd23861,17'd14811,17'd9743,17'd9479,17'd33083,17'd15944,17'd8883,17'd35515,17'd35516,17'd35517,17'd35518,17'd33573,17'd32597,17'd32769,17'd34209,17'd34386,17'd34047,17'd31590,17'd31442,17'd32436,17'd29066,17'd35519,17'd21504,17'd14523,17'd35520,17'd33583,17'd35521,17'd35102,17'd34966,17'd35103,17'd35104,17'd29938,17'd29795,17'd10731,17'd11272,17'd27344,17'd30692,17'd30705,17'd35522,17'd35379,17'd35523,17'd32148,17'd35524,17'd35525,17'd35526,17'd35527,17'd35528,17'd35529,17'd35530,17'd35531,17'd35532,17'd33269,17'd35533,17'd35534,17'd35535,17'd35536,17'd35537,17'd35538,17'd35539,17'd35540,17'd35541,17'd34074,17'd35542,17'd35543,17'd35544,17'd33921,17'd35267,17'd35267,17'd35545,17'd34594,17'd34858,17'd34594,17'd34247,17'd34593,17'd34592,17'd34428,17'd34735,17'd35136,17'd35132,17'd35546,17'd35547,17'd35548,17'd35549,17'd35271,17'd35550,17'd35551,17'd35552,17'd35553,17'd35554,17'd35555,17'd35556,17'd35557,17'd35558,17'd35559,17'd35560,17'd35561,17'd35562,17'd35563,17'd35564,17'd35565,17'd35285,17'd34444,17'd34096,17'd35421,17'd35421,17'd35566,17'd35286,17'd35008,17'd34752,17'd35009,17'd34754,17'd35567,17'd35568,17'd35569,17'd35570,17'd31035,17'd27259,17'd25707,17'd28594,17'd27637,17'd24415,17'd30127,17'd23569,17'd22856,17'd21847,17'd35571,17'd22001,17'd35294,17'd34456,17'd23220,17'd33944,17'd35429,17'd22503,17'd35430,17'd24902,17'd23564,17'd30431,17'd24898,17'd28369,17'd25565,17'd28853,17'd28727,17'd29977,17'd28134,17'd28134,17'd28134,17'd32355,17'd28372,17'd28728,17'd34114,17'd29833,17'd29979,17'd29690,17'd29536,17'd29381,17'd35431,17'd32024,17'd32359,17'd35572,17'd28860,17'd35433,17'd35573,17'd35574,17'd35575,17'd29388,17'd31369,17'd35576,17'd35437,17'd33673,17'd35577,17'd35439,17'd24743,17'd25180,17'd25709,17'd28594,17'd24736,17'd35578,17'd33500,17'd35441,17'd35579,17'd35580,17'd31665,17'd35581,17'd35582,17'd29395,17'd26540,17'd26913,17'd28617,17'd28505,17'd26798,17'd35583,17'd35584,17'd35311,17'd35585,17'd35586,17'd35587,17'd24752,17'd35588,17'd35589,17'd33509,17'd33163,17'd35590,17'd25826,17'd25699,17'd24408,17'd25438,17'd23916,17'd31836,17'd33479,17'd33480,17'd35591,17'd35592,17'd35593,17'd35594,17'd35595,17'd35596,17'd35597,17'd35598,17'd35599,17'd35600,17'd35601,17'd8603,17'd35602,17'd9367,17'd35603,17'd35468,17'd7654,17'd35604,17'd35605,17'd35606,17'd35607,17'd35608,17'd25361,17'd35609,17'd12162,17'd35610,17'd35610,17'd35051,17'd27934,17'd11037,17'd9933,17'd29593,17'd29593,17'd31243,17'd29593,17'd10515,17'd10642,17'd28184,17'd9091,17'd32073,17'd7499,17'd7499,17'd8780,17'd28058,17'd6220,17'd6390,17'd30333,17'd31553,17'd31717,17'd7499,17'd27815,17'd27933,17'd27933,17'd31551,17'd29158,17'd31551,17'd29593,17'd9934,17'd6223,17'd35197,17'd35479,17'd35480,17'd5923,17'd5485,17'd6228,17'd4380,17'd6399,17'd35200,17'd35611,17'd35612,17'd35613,17'd35614,17'd35615,17'd35616,17'd1379,17'd1681,17'd623,17'd3391,17'd4714,17'd35060,17'd5030,17'd2906,17'd5183,17'd9123,17'd9123,17'd8507,17'd7537,17'd9124,17'd9124,17'd33051,17'd35487,17'd31101,17'd31251,17'd31101,17'd31101,17'd31900,17'd31900,17'd29039,17'd29441,17'd31729,17'd28066,17'd5030,17'd16256,17'd12496,17'd11600,17'd5371,17'd1262,17'd428,17'd430,17'd18515,17'd35617,17'd35618,17'd34345
},
'{
17'd29756,17'd29756,17'd4087,17'd4425,17'd4428,17'd4577,17'd3252,17'd2422,17'd14070,17'd3101,17'd2593,17'd15496,17'd35619,17'd3101,17'd1831,17'd1127,17'd2597,17'd2257,17'd22965,17'd4089,17'd980,17'd286,17'd7061,17'd7728,17'd7556,17'd7225,17'd7226,17'd7062,17'd27445,17'd13067,17'd4896,17'd3260,17'd1705,17'd3599,17'd1707,17'd3917,17'd35620,17'd3436,17'd24510,17'd32255,17'd2796,17'd35621,17'd27102,17'd35622,17'd4108,17'd35623,17'd15886,17'd35624,17'd35625,17'd32260,17'd33548,17'd33548,17'd15384,17'd15384,17'd16168,17'd16169,17'd16986,17'd18774,17'd12681,17'd13211,17'd12954,17'd13092,17'd13462,17'd13462,17'd13092,17'd12813,17'd34181,17'd35626,17'd20429,17'd16884,17'd32741,17'd35627,17'd33224,17'd32742,17'd33386,17'd35356,17'd35628,17'd35629,17'd35630,17'd33390,17'd15782,17'd18178,17'd9992,17'd9583,17'd13611,17'd12685,17'd12686,17'd26856,17'd35631,17'd7921,17'd13612,17'd8701,17'd14640,17'd7763,17'd25514,17'd35632,17'd35633,17'd8705,17'd35634,17'd35635,17'd35636,17'd35637,17'd35638,17'd35639,17'd35640,17'd35641,17'd35642,17'd35643,17'd15048,17'd14928,17'd27490,17'd26875,17'd10336,17'd9041,17'd24361,17'd24040,17'd26039,17'd16916,17'd16917,17'd8421,17'd8419,17'd8731,17'd15430,17'd9479,17'd10331,17'd23166,17'd33572,17'd26493,17'd30831,17'd30833,17'd31287,17'd32920,17'd35644,17'd34380,17'd34203,17'd30221,17'd29645,17'd28103,17'd24537,17'd24208,17'd28112,17'd11668,17'd10328,17'd19918,17'd9347,17'd8720,17'd9189,17'd10174,17'd17480,17'd16317,17'd24368,17'd14812,17'd33715,17'd7947,17'd35645,17'd35646,17'd11137,17'd9046,17'd10336,17'd10335,17'd15569,17'd18080,17'd9041,17'd24367,17'd26631,17'd35647,17'd35648,17'd34208,17'd33092,17'd35649,17'd35650,17'd35651,17'd35652,17'd33882,17'd32592,17'd35653,17'd29329,17'd29778,17'd24991,17'd14672,17'd29339,17'd31777,17'd33736,17'd31954,17'd34966,17'd34966,17'd35103,17'd35654,17'd35655,17'd10598,17'd10322,17'd34051,17'd29661,17'd29799,17'd35656,17'd35379,17'd35657,17'd31968,17'd35658,17'd35659,17'd35660,17'd35661,17'd35662,17'd35663,17'd35664,17'd35665,17'd33120,17'd35666,17'd35667,17'd35668,17'd35669,17'd35670,17'd35671,17'd35672,17'd35673,17'd35674,17'd34854,17'd35675,17'd35676,17'd35677,17'd34430,17'd35678,17'd35679,17'd34247,17'd34247,17'd34429,17'd35680,17'd34079,17'd34079,17'd34079,17'd34428,17'd34593,17'd34735,17'd34735,17'd35546,17'd35546,17'd35403,17'd35681,17'd35403,17'd35133,17'd35682,17'd35683,17'd35684,17'd35552,17'd35685,17'd35686,17'd35687,17'd35688,17'd35689,17'd35690,17'd35691,17'd35692,17'd35693,17'd35694,17'd35695,17'd35696,17'd35697,17'd35698,17'd35699,17'd34444,17'd35700,17'd35701,17'd35566,17'd35702,17'd35008,17'd35703,17'd35009,17'd35423,17'd35704,17'd35705,17'd35706,17'd35707,17'd31035,17'd27027,17'd26903,17'd28723,17'd25178,17'd24416,17'd24086,17'd23567,17'd22680,17'd22507,17'd35708,17'd35709,17'd35710,17'd32664,17'd23220,17'd23393,17'd35711,17'd22329,17'd33794,17'd24086,17'd23385,17'd30431,17'd25180,17'd28369,17'd27766,17'd28725,17'd28727,17'd29977,17'd28134,17'd33654,17'd33654,17'd32017,17'd28372,17'd28728,17'd34285,17'd29833,17'd30130,17'd30884,17'd29106,17'd30740,17'd35712,17'd35713,17'd32197,17'd35572,17'd35714,17'd31049,17'd28868,17'd35715,17'd35716,17'd35717,17'd35718,17'd35719,17'd35720,17'd31195,17'd35721,17'd35722,17'd24252,17'd24898,17'd25568,17'd28598,17'd24736,17'd27025,17'd35723,17'd34632,17'd35724,17'd35725,17'd35726,17'd35727,17'd27152,17'd27535,17'd35728,17'd26540,17'd27168,17'd31363,17'd26798,17'd35729,17'd24757,17'd23941,17'd22883,17'd35730,17'd35731,17'd35732,17'd28261,17'd35733,17'd30001,17'd35734,17'd28980,17'd25557,17'd26055,17'd24242,17'd28600,17'd35735,17'd34298,17'd35736,17'd22158,17'd35737,17'd35738,17'd35739,17'd35740,17'd35741,17'd35742,17'd35743,17'd35744,17'd35745,17'd35746,17'd35747,17'd33832,17'd9213,17'd5475,17'd35748,17'd4353,17'd35749,17'd35750,17'd35751,17'd35752,17'd35753,17'd35754,17'd35755,17'd17536,17'd12161,17'd35756,17'd35757,17'd35758,17'd35759,17'd10642,17'd10514,17'd9933,17'd29592,17'd29593,17'd29593,17'd10515,17'd10515,17'd8780,17'd9091,17'd6219,17'd6220,17'd7499,17'd7668,17'd8780,17'd6391,17'd31717,17'd30638,17'd30638,17'd30333,17'd6390,17'd27696,17'd27933,17'd27933,17'd30933,17'd31551,17'd31551,17'd27933,17'd9934,17'd35760,17'd35197,17'd35479,17'd35480,17'd35761,17'd35762,17'd8636,17'd6073,17'd35763,17'd8311,17'd35764,17'd35765,17'd35766,17'd2551,17'd35767,17'd35768,17'd23814,17'd622,17'd443,17'd3895,17'd5630,17'd14586,17'd28657,17'd12495,17'd4714,17'd8186,17'd6416,17'd35769,17'd8507,17'd7705,17'd7705,17'd34002,17'd35487,17'd31101,17'd31101,17'd31101,17'd31101,17'd31900,17'd31900,17'd35770,17'd31101,17'd27949,17'd33050,17'd5777,17'd14586,17'd5630,17'd5371,17'd5050,17'd1262,17'd609,17'd1091,17'd786,17'd218,17'd35618,17'd35771
},
'{
17'd29756,17'd10533,17'd4087,17'd4425,17'd4428,17'd27591,17'd2935,17'd2422,17'd14070,17'd3101,17'd2593,17'd15496,17'd35619,17'd3101,17'd1831,17'd1127,17'd2596,17'd2257,17'd1416,17'd3905,17'd980,17'd286,17'd7061,17'd7728,17'd7556,17'd7225,17'd7226,17'd7062,17'd27445,17'd13067,17'd4896,17'd3260,17'd1705,17'd35772,17'd1707,17'd3917,17'd35620,17'd3436,17'd24510,17'd32255,17'd2796,17'd35621,17'd2626,17'd4752,17'd18159,17'd35773,17'd35774,17'd35775,17'd35776,17'd32099,17'd33548,17'd33548,17'd15384,17'd14767,17'd16411,17'd18657,17'd16986,17'd20422,17'd16658,17'd13211,17'd12954,17'd13092,17'd13462,17'd14469,17'd13092,17'd35352,17'd35777,17'd35778,17'd14349,17'd35779,17'd32263,17'd33065,17'd33224,17'd34678,17'd35780,17'd35356,17'd35781,17'd35629,17'd35782,17'd35783,17'd35784,17'd35359,17'd9849,17'd9583,17'd13611,17'd14640,17'd35631,17'd35785,17'd7104,17'd26742,17'd8077,17'd8701,17'd13612,17'd7921,17'd25514,17'd35786,17'd35787,17'd8705,17'd35788,17'd35789,17'd35790,17'd35791,17'd35792,17'd35793,17'd35794,17'd35795,17'd35796,17'd24037,17'd9619,17'd11277,17'd19531,17'd16328,17'd10175,17'd9041,17'd24361,17'd24040,17'd35797,17'd35798,17'd16917,17'd34036,17'd12119,17'd8729,17'd15944,17'd9885,17'd19280,17'd35799,17'd35800,17'd26493,17'd30071,17'd32919,17'd31127,17'd32920,17'd31590,17'd34037,17'd34835,17'd30073,17'd35372,17'd28816,17'd26493,17'd27985,17'd35801,17'd12423,17'd16796,17'd18332,17'd8873,17'd8720,17'd9189,17'd17480,17'd26498,17'd26259,17'd35514,17'd12426,17'd8252,17'd7947,17'd35645,17'd24043,17'd11137,17'd9046,17'd10336,17'd26153,17'd15807,17'd17716,17'd8884,17'd10337,17'd27988,17'd35802,17'd35803,17'd34542,17'd30974,17'd35804,17'd32929,17'd35805,17'd34211,17'd33882,17'd31127,17'd33718,17'd30831,17'd28347,17'd16556,17'd14525,17'd35806,17'd31777,17'd33736,17'd31954,17'd34966,17'd35103,17'd35241,17'd35242,17'd35807,17'd10323,17'd29796,17'd35808,17'd35809,17'd35810,17'd35379,17'd35811,17'd32307,17'd35812,17'd33743,17'd35813,17'd35814,17'd35815,17'd35816,17'd35817,17'd35818,17'd35819,17'd35820,17'd35821,17'd35822,17'd35823,17'd35670,17'd35824,17'd35825,17'd35826,17'd35827,17'd35828,17'd35829,17'd35830,17'd35831,17'd35832,17'd35833,17'd35834,17'd35835,17'd35836,17'd34078,17'd34078,17'd35837,17'd34429,17'd35680,17'd35680,17'd34594,17'd34428,17'd34593,17'd34593,17'd35546,17'd35681,17'd35681,17'd35547,17'd35546,17'd35548,17'd35838,17'd35839,17'd35406,17'd35684,17'd35840,17'd35686,17'd35841,17'd35842,17'd35843,17'd35844,17'd35845,17'd35846,17'd35847,17'd35848,17'd35147,17'd35849,17'd35850,17'd35285,17'd35699,17'd33936,17'd35700,17'd35701,17'd35566,17'd35702,17'd35851,17'd34752,17'd35852,17'd35423,17'd35704,17'd35705,17'd35853,17'd35854,17'd30735,17'd30586,17'd28725,17'd27766,17'd25709,17'd24745,17'd23731,17'd29099,17'd23389,17'd22159,17'd22003,17'd21699,17'd35855,17'd35856,17'd32829,17'd30728,17'd35429,17'd22328,17'd33950,17'd30879,17'd29377,17'd30431,17'd25030,17'd27882,17'd27766,17'd28725,17'd28727,17'd33001,17'd33654,17'd33654,17'd33654,17'd32017,17'd28372,17'd28372,17'd29249,17'd29833,17'd29978,17'd30884,17'd29106,17'd29833,17'd35712,17'd34623,17'd35857,17'd35168,17'd35858,17'd35859,17'd35860,17'd35861,17'd35862,17'd35863,17'd35718,17'd35864,17'd35720,17'd35865,17'd35577,17'd35722,17'd24252,17'd24898,17'd25568,17'd25567,17'd24891,17'd33815,17'd34301,17'd35866,17'd35724,17'd35725,17'd35867,17'd35307,17'd27380,17'd27265,17'd26296,17'd27664,17'd27276,17'd34471,17'd35868,17'd35869,17'd35870,17'd35871,17'd35872,17'd31859,17'd23584,17'd32377,17'd35873,17'd35874,17'd35875,17'd35876,17'd35866,17'd25944,17'd25559,17'd25707,17'd26402,17'd29386,17'd35877,17'd23572,17'd30426,17'd23743,17'd35878,17'd24426,17'd35879,17'd35880,17'd35881,17'd35882,17'd35883,17'd35884,17'd35885,17'd35886,17'd35887,17'd35467,17'd35888,17'd35889,17'd4353,17'd3830,17'd33204,17'd35890,17'd35891,17'd35754,17'd29298,17'd35755,17'd15728,17'd12307,17'd35892,17'd35757,17'd35477,17'd35893,17'd10515,17'd10515,17'd29593,17'd29592,17'd29593,17'd29593,17'd10515,17'd10515,17'd27815,17'd7499,17'd6390,17'd6219,17'd9091,17'd7499,17'd8780,17'd7668,17'd6554,17'd30638,17'd5160,17'd30333,17'd6390,17'd7668,17'd10515,17'd28183,17'd31551,17'd31551,17'd31551,17'd27933,17'd9934,17'd6223,17'd35197,17'd35479,17'd35894,17'd35895,17'd35896,17'd35897,17'd35898,17'd35899,17'd35900,17'd35901,17'd35902,17'd35903,17'd35904,17'd35905,17'd35906,17'd24496,17'd244,17'd428,17'd445,17'd8185,17'd14586,17'd35060,17'd12495,17'd9123,17'd8186,17'd8186,17'd35769,17'd8507,17'd7537,17'd7537,17'd34002,17'd35487,17'd31101,17'd31251,17'd31101,17'd31101,17'd31900,17'd31900,17'd35770,17'd31101,17'd27949,17'd28066,17'd5030,17'd14586,17'd5630,17'd35907,17'd5371,17'd1262,17'd609,17'd35908,17'd18515,17'd585,17'd35909,17'd35910
},
'{
17'd4891,17'd3902,17'd3902,17'd4425,17'd4428,17'd4577,17'd3252,17'd2422,17'd3101,17'd3101,17'd2934,17'd15877,17'd35619,17'd3101,17'd1831,17'd4247,17'd2596,17'd1414,17'd1416,17'd3905,17'd980,17'd286,17'd7061,17'd7061,17'd7225,17'd7225,17'd6599,17'd5972,17'd27445,17'd34004,17'd4253,17'd3107,17'd1706,17'd1707,17'd4095,17'd3917,17'd35620,17'd3436,17'd3264,17'd32090,17'd30050,17'd27830,17'd35911,17'd4592,17'd18524,17'd35912,17'd35913,17'd35914,17'd35915,17'd32099,17'd33548,17'd33548,17'd14893,17'd16881,17'd16169,17'd19383,17'd18774,17'd20423,17'd13969,17'd13211,17'd12954,17'd13092,17'd14469,17'd12357,17'd13092,17'd9836,17'd19623,17'd18416,17'd35916,17'd35917,17'd32572,17'd34944,17'd33224,17'd33703,17'd33555,17'd35072,17'd35629,17'd34367,17'd35918,17'd35919,17'd35920,17'd14230,17'd9849,17'd9310,17'd14231,17'd35218,17'd7104,17'd7104,17'd7104,17'd35631,17'd13612,17'd8701,17'd13612,17'd7921,17'd7104,17'd35786,17'd35921,17'd35078,17'd35922,17'd35923,17'd35924,17'd35925,17'd35926,17'd35927,17'd35928,17'd35929,17'd28702,17'd15569,17'd9619,17'd17011,17'd11809,17'd10335,17'd9041,17'd9041,17'd17716,17'd33238,17'd35930,17'd10340,17'd16917,17'd33874,17'd9887,17'd25677,17'd15180,17'd9741,17'd11400,17'd18326,17'd26258,17'd29196,17'd35931,17'd30834,17'd31127,17'd32920,17'd34037,17'd31288,17'd31767,17'd29930,17'd28460,17'd27121,17'd24030,17'd29928,17'd13367,17'd19280,17'd17012,17'd9338,17'd8720,17'd9040,17'd9038,17'd10174,17'd9041,17'd24368,17'd24213,17'd17849,17'd14527,17'd14527,17'd10608,17'd14135,17'd10607,17'd9040,17'd15684,17'd10336,17'd10335,17'd10174,17'd8880,17'd17848,17'd35932,17'd32764,17'd34962,17'd29924,17'd34381,17'd35933,17'd35238,17'd35934,17'd34387,17'd33096,17'd31128,17'd30072,17'd35376,17'd28107,17'd21504,17'd29208,17'd35520,17'd33416,17'd33736,17'd34966,17'd33250,17'd33103,17'd35935,17'd35655,17'd10468,17'd35936,17'd34396,17'd29501,17'd35937,17'd35938,17'd35523,17'd35939,17'd31786,17'd34974,17'd35940,17'd35941,17'd35942,17'd35943,17'd35944,17'd35945,17'd35946,17'd35947,17'd35948,17'd35949,17'd35950,17'd35951,17'd35952,17'd35953,17'd35954,17'd35955,17'd35956,17'd35957,17'd35958,17'd34736,17'd35959,17'd35960,17'd35961,17'd35683,17'd35962,17'd35963,17'd34077,17'd35964,17'd34077,17'd35965,17'd35966,17'd35966,17'd35837,17'd35967,17'd34247,17'd34593,17'd34735,17'd34592,17'd35681,17'd35547,17'd35547,17'd35968,17'd35969,17'd35970,17'd35971,17'd35972,17'd35973,17'd35974,17'd35975,17'd35976,17'd35977,17'd35978,17'd35979,17'd35980,17'd35981,17'd35982,17'd35983,17'd35984,17'd35850,17'd35985,17'd35699,17'd33936,17'd35986,17'd35700,17'd35566,17'd35702,17'd35148,17'd35008,17'd35987,17'd35988,17'd35704,17'd35705,17'd35989,17'd35990,17'd35426,17'd33163,17'd27258,17'd26174,17'd28597,17'd25029,17'd24252,17'd23733,17'd32351,17'd22333,17'd22004,17'd22494,17'd35991,17'd35992,17'd30727,17'd22682,17'd35296,17'd22503,17'd33950,17'd23732,17'd23385,17'd30431,17'd25030,17'd25709,17'd28602,17'd28725,17'd28979,17'd29977,17'd28134,17'd33654,17'd33654,17'd32355,17'd29380,17'd28372,17'd29249,17'd34114,17'd29978,17'd30884,17'd29691,17'd29833,17'd35712,17'd35297,17'd31355,17'd35026,17'd30000,17'd35993,17'd26066,17'd35994,17'd35995,17'd35996,17'd35997,17'd35998,17'd24746,17'd29530,17'd35999,17'd24089,17'd24743,17'd24745,17'd27637,17'd28597,17'd24891,17'd36000,17'd27883,17'd35866,17'd35724,17'd36001,17'd36002,17'd31199,17'd30745,17'd31041,17'd29543,17'd34771,17'd36003,17'd32034,17'd31848,17'd34473,17'd28624,17'd35871,17'd36004,17'd36005,17'd23584,17'd36006,17'd36007,17'd27890,17'd35433,17'd32515,17'd36008,17'd28486,17'd25559,17'd25831,17'd26064,17'd25318,17'd35577,17'd31836,17'd36009,17'd32009,17'd36010,17'd36011,17'd36012,17'd36013,17'd36014,17'd36015,17'd36016,17'd36017,17'd36018,17'd36019,17'd30932,17'd6377,17'd36020,17'd35889,17'd36021,17'd36021,17'd36022,17'd36023,17'd36024,17'd36025,17'd36026,17'd36027,17'd35755,17'd17536,17'd36028,17'd36029,17'd36030,17'd36031,17'd10515,17'd10515,17'd29592,17'd29592,17'd9933,17'd9933,17'd27933,17'd10642,17'd27815,17'd7499,17'd6390,17'd6390,17'd6219,17'd6220,17'd8780,17'd8780,17'd6390,17'd28185,17'd5160,17'd25627,17'd27935,17'd7499,17'd27815,17'd28183,17'd31551,17'd31551,17'd31551,17'd27933,17'd9934,17'd6223,17'd35197,17'd36032,17'd36033,17'd35895,17'd36034,17'd36035,17'd36036,17'd36037,17'd36038,17'd36039,17'd36040,17'd36041,17'd36042,17'd36043,17'd36044,17'd1665,17'd784,17'd233,17'd1261,17'd35907,17'd16256,17'd15233,17'd5777,17'd9123,17'd7365,17'd8186,17'd36045,17'd6417,17'd7537,17'd7537,17'd34002,17'd35487,17'd31101,17'd31251,17'd31101,17'd31101,17'd31251,17'd31251,17'd28793,17'd27708,17'd27949,17'd33050,17'd5777,17'd14586,17'd5940,17'd5371,17'd2392,17'd1262,17'd609,17'd29749,17'd18515,17'd36046,17'd36047,17'd36048
},
'{
17'd4891,17'd3902,17'd3902,17'd4891,17'd4428,17'd27591,17'd2935,17'd3252,17'd3101,17'd2934,17'd3751,17'd15877,17'd35619,17'd2935,17'd1831,17'd4247,17'd2596,17'd1414,17'd1416,17'd3905,17'd980,17'd286,17'd7061,17'd7061,17'd7225,17'd7225,17'd6599,17'd26971,17'd5810,17'd34004,17'd4253,17'd2607,17'd1706,17'd35772,17'd2786,17'd4095,17'd2609,17'd3436,17'd3264,17'd32090,17'd31106,17'd27957,17'd3767,17'd4908,17'd28198,17'd36049,17'd36050,17'd36051,17'd35915,17'd32099,17'd33548,17'd15384,17'd14767,17'd16411,17'd17690,17'd18656,17'd17689,17'd22630,17'd14622,17'd17096,17'd12954,17'd13092,17'd14469,17'd12357,17'd35352,17'd36052,17'd35212,17'd36053,17'd35779,17'd32263,17'd33224,17'd34184,17'd33224,17'd35497,17'd34187,17'd35072,17'd36054,17'd34367,17'd36055,17'd36056,17'd14782,17'd12822,17'd9583,17'd9165,17'd14640,17'd35631,17'd36057,17'd35632,17'd7104,17'd25514,17'd8077,17'd13612,17'd13612,17'd7921,17'd7104,17'd36058,17'd36059,17'd35078,17'd36060,17'd36061,17'd36062,17'd36063,17'd36064,17'd36065,17'd36066,17'd36067,17'd36068,17'd15807,17'd11809,17'd15187,17'd14674,17'd10336,17'd8885,17'd16317,17'd36069,17'd33238,17'd23342,17'd36070,17'd34040,17'd25289,17'd24545,17'd24212,17'd9345,17'd12116,17'd11400,17'd36071,17'd35800,17'd29065,17'd30675,17'd32283,17'd31442,17'd32920,17'd33875,17'd34203,17'd30677,17'd29198,17'd30222,17'd26370,17'd24538,17'd24363,17'd36072,17'd17847,17'd10857,17'd9192,17'd9044,17'd9194,17'd10174,17'd9038,17'd9348,17'd11404,17'd12867,17'd8581,17'd17128,17'd17850,17'd8580,17'd9349,17'd8725,17'd9040,17'd9194,17'd10336,17'd10335,17'd22645,17'd36073,17'd26632,17'd36074,17'd36075,17'd31594,17'd29067,17'd34704,17'd34833,17'd34044,17'd36076,17'd33095,17'd31591,17'd30677,17'd31286,17'd28347,17'd16557,17'd14525,17'd36077,17'd34708,17'd33736,17'd34966,17'd33102,17'd33250,17'd34214,17'd36078,17'd36079,17'd27001,17'd36080,17'd29809,17'd36081,17'd36082,17'd29945,17'd30391,17'd30851,17'd36083,17'd31624,17'd36084,17'd36085,17'd35816,17'd36086,17'd36087,17'd36088,17'd36089,17'd36090,17'd36091,17'd36092,17'd36093,17'd36094,17'd36095,17'd36096,17'd36097,17'd36098,17'd36099,17'd34734,17'd36100,17'd36101,17'd36102,17'd36103,17'd36104,17'd36105,17'd35971,17'd35684,17'd36106,17'd35839,17'd35970,17'd36107,17'd36108,17'd35964,17'd36109,17'd35966,17'd34593,17'd34593,17'd34735,17'd34592,17'd35403,17'd35546,17'd35546,17'd35546,17'd36110,17'd36111,17'd36105,17'd35971,17'd36112,17'd35974,17'd36113,17'd36114,17'd36115,17'd35557,17'd36116,17'd36117,17'd36118,17'd36119,17'd36120,17'd36121,17'd36122,17'd35985,17'd35699,17'd33936,17'd35986,17'd35700,17'd35702,17'd36123,17'd35286,17'd34101,17'd35008,17'd36124,17'd35704,17'd35568,17'd36125,17'd36126,17'd36127,17'd30735,17'd30586,17'd26903,17'd27638,17'd27512,17'd24417,17'd30879,17'd23923,17'd22678,17'd36128,17'd36129,17'd21692,17'd36130,17'd30727,17'd36131,17'd35296,17'd22502,17'd33950,17'd30275,17'd23385,17'd30431,17'd24898,17'd25709,17'd27766,17'd28725,17'd28979,17'd33952,17'd28134,17'd33654,17'd33654,17'd32355,17'd29380,17'd29248,17'd29249,17'd34114,17'd29981,17'd30884,17'd30884,17'd36132,17'd29107,17'd35431,17'd36133,17'd35026,17'd36134,17'd36135,17'd26066,17'd36136,17'd27030,17'd30150,17'd36137,17'd36138,17'd36139,17'd29530,17'd23921,17'd24088,17'd24743,17'd24745,17'd27637,17'd27882,17'd23909,17'd25832,17'd33815,17'd34128,17'd36140,17'd36141,17'd36142,17'd35572,17'd36143,17'd33004,17'd27380,17'd27270,17'd29558,17'd36144,17'd27162,17'd26084,17'd36145,17'd26672,17'd36146,17'd36147,17'd36148,17'd36149,17'd36150,17'd35873,17'd36151,17'd32849,17'd27517,17'd34479,17'd34637,17'd28365,17'd28481,17'd25436,17'd24250,17'd36152,17'd35018,17'd32346,17'd36153,17'd36154,17'd36155,17'd36156,17'd36157,17'd36158,17'd36159,17'd21740,17'd36160,17'd36161,17'd36162,17'd36163,17'd36164,17'd36165,17'd33990,17'd34649,17'd36166,17'd36167,17'd36168,17'd35753,17'd36169,17'd36027,17'd35755,17'd17536,17'd17535,17'd19222,17'd36170,17'd36171,17'd10642,17'd10515,17'd29592,17'd29592,17'd9933,17'd9933,17'd27933,17'd28183,17'd10515,17'd7668,17'd6390,17'd31717,17'd6390,17'd6390,17'd7668,17'd8780,17'd6219,17'd28185,17'd5160,17'd25627,17'd28185,17'd6219,17'd8780,17'd10642,17'd28057,17'd31551,17'd30933,17'd27933,17'd9934,17'd6223,17'd35197,17'd36172,17'd36173,17'd35895,17'd36034,17'd36035,17'd36174,17'd36175,17'd36176,17'd36177,17'd36178,17'd36179,17'd23298,17'd36180,17'd19730,17'd36181,17'd35059,17'd793,17'd625,17'd3391,17'd14178,17'd5631,17'd2906,17'd8186,17'd7365,17'd8186,17'd36045,17'd6417,17'd7537,17'd7537,17'd34002,17'd33051,17'd31101,17'd31251,17'd31251,17'd31101,17'd31251,17'd31251,17'd29170,17'd27708,17'd27949,17'd33050,17'd5777,17'd14586,17'd5940,17'd5371,17'd2392,17'd625,17'd1122,17'd29749,17'd18515,17'd31730,17'd36182,17'd34668
},
'{
17'd4891,17'd3902,17'd3902,17'd27713,17'd3427,17'd2592,17'd3252,17'd3252,17'd3101,17'd3251,17'd2934,17'd15877,17'd35619,17'd2935,17'd1831,17'd4247,17'd2596,17'd1414,17'd1416,17'd3905,17'd27,17'd285,17'd7061,17'd7061,17'd7225,17'd7225,17'd6599,17'd26971,17'd5810,17'd4895,17'd4253,17'd2607,17'd1706,17'd1707,17'd4095,17'd4095,17'd2609,17'd36183,17'd3264,17'd32886,17'd31106,17'd2958,17'd36184,17'd31107,17'd36185,17'd36186,17'd36187,17'd36188,17'd34937,17'd32099,17'd33548,17'd15384,17'd14768,17'd24520,17'd18657,17'd18655,17'd19382,17'd16658,17'd17940,17'd13599,17'd13092,17'd12678,17'd12357,17'd12357,17'd11475,17'd34939,17'd36189,17'd17211,17'd36190,17'd34678,17'd34944,17'd36191,17'd36192,17'd33386,17'd35356,17'd35073,17'd35358,17'd33706,17'd35919,17'd36193,17'd15150,17'd9444,17'd9310,17'd12370,17'd12371,17'd35631,17'd36057,17'd36194,17'd36195,17'd25514,17'd7921,17'd13612,17'd13612,17'd35631,17'd35500,17'd36058,17'd36059,17'd36196,17'd36197,17'd36061,17'd36198,17'd36199,17'd36200,17'd36201,17'd36202,17'd36203,17'd16441,17'd14811,17'd15187,17'd27856,17'd13887,17'd8873,17'd15297,17'd9194,17'd25408,17'd17472,17'd15945,17'd36070,17'd12427,17'd36204,17'd36205,17'd10336,17'd27856,17'd9740,17'd11400,17'd36206,17'd26151,17'd32435,17'd34827,17'd31941,17'd31127,17'd31442,17'd33875,17'd34203,17'd30073,17'd29201,17'd28104,17'd25927,17'd24992,17'd14259,17'd28821,17'd13522,17'd9342,17'd24039,17'd9044,17'd9194,17'd10174,17'd8873,17'd15297,17'd15568,17'd8419,17'd17241,17'd17017,17'd17850,17'd8580,17'd17481,17'd8724,17'd9041,17'd9194,17'd10336,17'd16552,17'd36207,17'd26633,17'd36208,17'd36209,17'd36210,17'd26873,17'd36211,17'd34704,17'd33574,17'd36212,17'd36213,17'd31591,17'd36214,17'd29482,17'd29336,17'd35240,17'd16913,17'd13643,17'd36215,17'd31602,17'd33736,17'd32939,17'd31451,17'd36216,17'd35935,17'd36217,17'd36218,17'd11272,17'd29495,17'd36219,17'd36220,17'd36221,17'd29946,17'd36222,17'd31150,17'd36223,17'd36224,17'd31797,17'd36225,17'd36226,17'd36227,17'd36228,17'd36229,17'd36230,17'd36231,17'd36232,17'd36233,17'd36234,17'd36235,17'd35672,17'd36236,17'd36237,17'd36238,17'd36239,17'd36240,17'd34250,17'd36241,17'd35965,17'd35682,17'd36106,17'd36242,17'd35683,17'd35683,17'd36105,17'd36243,17'd36244,17'd35972,17'd36245,17'd36246,17'd36247,17'd35274,17'd35132,17'd34735,17'd34593,17'd34735,17'd35403,17'd35403,17'd35546,17'd35547,17'd35968,17'd36248,17'd35405,17'd35550,17'd35679,17'd36249,17'd36250,17'd36251,17'd36252,17'd36253,17'd36254,17'd36255,17'd36256,17'd36257,17'd36258,17'd36259,17'd36122,17'd35985,17'd35699,17'd35699,17'd36260,17'd35700,17'd35702,17'd35702,17'd36261,17'd34101,17'd35008,17'd36262,17'd36263,17'd35705,17'd36125,17'd35706,17'd36264,17'd35011,17'd27146,17'd28724,17'd28594,17'd25568,17'd24896,17'd23917,17'd35865,17'd22331,17'd22165,17'd22011,17'd21698,17'd22003,17'd22156,17'd32999,17'd31343,17'd22503,17'd31029,17'd23564,17'd23385,17'd29375,17'd24745,17'd25438,17'd25566,17'd28724,17'd28486,17'd33952,17'd32354,17'd32354,17'd32192,17'd32017,17'd29248,17'd29249,17'd29249,17'd34114,17'd29981,17'd29690,17'd30884,17'd36132,17'd29107,17'd35431,17'd36265,17'd36266,17'd31210,17'd36267,17'd36268,17'd36269,17'd36270,17'd36271,17'd36272,17'd36273,17'd36274,17'd29530,17'd23921,17'd25439,17'd24090,17'd24745,17'd28254,17'd25709,17'd24892,17'd25434,17'd28482,17'd27027,17'd29379,17'd35579,17'd28859,17'd29383,17'd31199,17'd30592,17'd33004,17'd36275,17'd36276,17'd27529,17'd26920,17'd25720,17'd36145,17'd24432,17'd36277,17'd36278,17'd36279,17'd36280,17'd36281,17'd36282,17'd28021,17'd36283,17'd36284,17'd36285,17'd35011,17'd36286,17'd27514,17'd28600,17'd36287,17'd35877,17'd36288,17'd36289,17'd36290,17'd36291,17'd36292,17'd36293,17'd34320,17'd36294,17'd36295,17'd36296,17'd36297,17'd36298,17'd36299,17'd35887,17'd36300,17'd35748,17'd36301,17'd36302,17'd36303,17'd36304,17'd36305,17'd36306,17'd36026,17'd35754,17'd36307,17'd36308,17'd24802,17'd36309,17'd36170,17'd36310,17'd10642,17'd10515,17'd27933,17'd29592,17'd9933,17'd9933,17'd27933,17'd27933,17'd10515,17'd8780,17'd6390,17'd28185,17'd27935,17'd6554,17'd7499,17'd8780,17'd6220,17'd27935,17'd5160,17'd25627,17'd30638,17'd6554,17'd7668,17'd10515,17'd28057,17'd28183,17'd30933,17'd27933,17'd9934,17'd6223,17'd36311,17'd36032,17'd36312,17'd35895,17'd35896,17'd36313,17'd36314,17'd36315,17'd36316,17'd36317,17'd36318,17'd36319,17'd36320,17'd36321,17'd19863,17'd36322,17'd36323,17'd630,17'd446,17'd3895,17'd14178,17'd6721,17'd2906,17'd8186,17'd7365,17'd6258,17'd6417,17'd6418,17'd7537,17'd7537,17'd34002,17'd33051,17'd31101,17'd31251,17'd31101,17'd31101,17'd31101,17'd31251,17'd29170,17'd27708,17'd27949,17'd33050,17'd5777,17'd2098,17'd6415,17'd5371,17'd2392,17'd1262,17'd609,17'd29749,17'd767,17'd36324,17'd34667,17'd36325
},
'{
17'd4891,17'd3902,17'd4244,17'd4891,17'd3901,17'd6424,17'd2935,17'd3252,17'd3101,17'd3427,17'd3901,17'd15877,17'd15358,17'd2935,17'd1831,17'd1127,17'd2597,17'd1414,17'd1416,17'd3905,17'd27,17'd285,17'd7061,17'd7061,17'd7225,17'd7225,17'd6599,17'd26971,17'd5810,17'd4741,17'd4253,17'd2607,17'd1706,17'd35772,17'd4095,17'd4095,17'd2609,17'd36183,17'd3266,17'd32886,17'd31106,17'd2958,17'd36184,17'd5070,17'd36326,17'd15633,17'd36327,17'd35625,17'd34937,17'd31918,17'd15519,17'd14892,17'd16768,17'd17690,17'd19008,17'd18774,17'd19382,17'd12361,17'd17096,17'd12954,17'd13092,17'd12678,17'd12357,17'd15516,17'd36328,17'd36329,17'd36330,17'd17944,17'd36331,17'd33224,17'd33861,17'd33861,17'd36332,17'd36333,17'd35214,17'd36334,17'd35358,17'd33228,17'd36335,17'd15914,17'd15150,17'd9445,17'd11095,17'd12370,17'd12371,17'd25126,17'd36336,17'd36336,17'd35632,17'd25514,17'd7921,17'd13612,17'd35218,17'd35631,17'd35500,17'd7107,17'd36337,17'd36338,17'd36197,17'd36339,17'd36340,17'd36341,17'd36342,17'd36343,17'd36344,17'd36345,17'd8876,17'd17480,17'd15187,17'd13887,17'd9038,17'd9040,17'd8881,17'd9194,17'd22814,17'd17123,17'd8414,17'd36070,17'd8734,17'd23866,17'd26259,17'd22813,17'd9341,17'd17719,17'd12423,17'd36071,17'd36346,17'd29197,17'd34827,17'd32283,17'd31442,17'd32920,17'd33875,17'd33568,17'd29785,17'd36347,17'd28103,17'd25927,17'd24992,17'd36348,17'd36349,17'd16912,17'd9339,17'd8720,17'd9045,17'd15684,17'd8874,17'd8720,17'd12118,17'd8246,17'd17483,17'd17016,17'd16333,17'd17352,17'd12119,17'd15429,17'd8878,17'd9045,17'd9194,17'd10336,17'd26153,17'd32924,17'd28113,17'd36350,17'd36351,17'd36352,17'd28103,17'd36353,17'd34835,17'd36354,17'd36355,17'd32920,17'd33568,17'd30371,17'd36347,17'd27235,17'd27486,17'd14524,17'd29340,17'd34708,17'd32447,17'd34966,17'd36356,17'd31451,17'd34214,17'd36078,17'd36357,17'd36358,17'd36080,17'd36359,17'd30860,17'd29801,17'd29947,17'd36360,17'd30852,17'd36361,17'd36362,17'd36363,17'd36225,17'd36364,17'd36365,17'd36366,17'd36367,17'd36368,17'd36369,17'd36370,17'd36371,17'd36372,17'd36373,17'd36374,17'd36375,17'd36376,17'd36377,17'd34733,17'd36378,17'd36379,17'd33769,17'd34593,17'd36380,17'd35838,17'd36381,17'd36382,17'd35970,17'd35839,17'd35683,17'd36383,17'd36384,17'd36385,17'd36385,17'd36385,17'd35971,17'd36246,17'd36386,17'd35136,17'd34735,17'd34735,17'd35681,17'd35403,17'd35403,17'd35546,17'd35968,17'd35404,17'd36387,17'd35405,17'd36388,17'd36249,17'd36389,17'd36390,17'd36391,17'd36392,17'd36393,17'd36394,17'd36395,17'd36396,17'd36397,17'd36259,17'd36122,17'd35420,17'd35985,17'd35699,17'd36260,17'd35700,17'd35566,17'd35702,17'd36398,17'd36399,17'd34874,17'd36400,17'd36401,17'd35705,17'd36125,17'd36402,17'd36403,17'd35426,17'd33163,17'd28978,17'd28723,17'd28717,17'd28596,17'd34467,17'd30127,17'd22503,17'd30727,17'd22010,17'd22169,17'd36404,17'd32345,17'd22324,17'd31343,17'd22328,17'd30127,17'd23384,17'd23385,17'd24087,17'd24417,17'd25177,17'd25566,17'd28724,17'd28486,17'd29379,17'd27885,17'd32354,17'd32192,17'd32017,17'd29248,17'd29249,17'd36405,17'd36406,17'd32508,17'd32833,17'd29690,17'd29978,17'd34114,17'd36407,17'd36408,17'd29695,17'd31210,17'd31361,17'd25836,17'd36409,17'd36410,17'd36411,17'd36412,17'd36413,17'd36414,17'd35865,17'd23921,17'd24088,17'd28601,17'd24744,17'd28254,17'd28717,17'd27257,17'd25564,17'd27639,17'd26902,17'd26780,17'd30279,17'd28011,17'd36415,17'd35572,17'd35307,17'd36416,17'd36417,17'd36418,17'd30145,17'd26410,17'd27160,17'd26420,17'd28747,17'd36419,17'd36420,17'd32216,17'd30761,17'd36421,17'd36422,17'd36423,17'd28380,17'd36424,17'd36425,17'd34637,17'd27369,17'd28725,17'd28723,17'd33969,17'd35577,17'd36426,17'd36427,17'd36428,17'd34907,17'd36429,17'd36430,17'd36431,17'd36432,17'd36433,17'd36434,17'd20983,17'd36435,17'd36436,17'd21588,17'd36437,17'd36438,17'd36301,17'd36302,17'd36303,17'd36439,17'd36440,17'd36441,17'd36025,17'd36026,17'd36442,17'd36443,17'd29297,17'd36028,17'd36170,17'd36444,17'd11316,17'd10642,17'd27933,17'd27933,17'd9933,17'd9933,17'd29592,17'd27933,17'd10515,17'd28184,17'd6219,17'd30638,17'd28185,17'd31717,17'd9091,17'd8780,17'd7499,17'd27935,17'd5160,17'd25627,17'd30333,17'd31717,17'd7499,17'd27815,17'd28183,17'd28183,17'd30933,17'd27933,17'd9934,17'd6558,17'd36311,17'd36172,17'd36173,17'd35895,17'd35896,17'd36445,17'd36446,17'd36447,17'd36448,17'd36449,17'd36450,17'd36451,17'd36452,17'd36321,17'd36453,17'd36454,17'd36455,17'd18144,17'd1825,17'd1119,17'd2097,17'd4559,17'd9544,17'd7365,17'd6095,17'd6258,17'd6417,17'd6418,17'd7537,17'd7537,17'd34002,17'd33051,17'd31101,17'd31251,17'd31101,17'd31101,17'd31101,17'd31251,17'd27708,17'd27708,17'd27949,17'd33050,17'd5777,17'd2098,17'd6415,17'd5371,17'd2392,17'd625,17'd1122,17'd29749,17'd787,17'd36456,17'd35209,17'd36457
},
'{
17'd4891,17'd3902,17'd4244,17'd27713,17'd3427,17'd2592,17'd14070,17'd3252,17'd3101,17'd3251,17'd3427,17'd15877,17'd15358,17'd2784,17'd1831,17'd1127,17'd2597,17'd2257,17'd1416,17'd1128,17'd26,17'd285,17'd7061,17'd7061,17'd7225,17'd6599,17'd6440,17'd26971,17'd26605,17'd4740,17'd36458,17'd2608,17'd1841,17'd35772,17'd4095,17'd3918,17'd2609,17'd3600,17'd3436,17'd32731,17'd31106,17'd2958,17'd4591,17'd36459,17'd26134,17'd36460,17'd36461,17'd36462,17'd34937,17'd31918,17'd14893,17'd14768,17'd16411,17'd17690,17'd19255,17'd17689,17'd19006,17'd14470,17'd17809,17'd12954,17'd13092,17'd12678,17'd15763,17'd15516,17'd36463,17'd36464,17'd20430,17'd16414,17'd36465,17'd34944,17'd36191,17'd36466,17'd36467,17'd33555,17'd36468,17'd36469,17'd35216,17'd32268,17'd35217,17'd14782,17'd15023,17'd9583,17'd11631,17'd14231,17'd36470,17'd25126,17'd36471,17'd36472,17'd35632,17'd25126,17'd24980,17'd27835,17'd36473,17'd35631,17'd35500,17'd7107,17'd36337,17'd35221,17'd36197,17'd36339,17'd36474,17'd36475,17'd36342,17'd36476,17'd36477,17'd9184,17'd8876,17'd10336,17'd9345,17'd9347,17'd11402,17'd15297,17'd8882,17'd9041,17'd14674,17'd15684,17'd8416,17'd36478,17'd18203,17'd26262,17'd26154,17'd26153,17'd9341,17'd9740,17'd15176,17'd36071,17'd36479,17'd36480,17'd32919,17'd31287,17'd34037,17'd34037,17'd34203,17'd34835,17'd30220,17'd34390,17'd26629,17'd25925,17'd24362,17'd36481,17'd36482,17'd13255,17'd9192,17'd8720,17'd9041,17'd10336,17'd9189,17'd19033,17'd11403,17'd36483,17'd17483,17'd16333,17'd17016,17'd25411,17'd24213,17'd11966,17'd8885,17'd29334,17'd9041,17'd17480,17'd22813,17'd36484,17'd36485,17'd27865,17'd36486,17'd36487,17'd36488,17'd30678,17'd33409,17'd36354,17'd36489,17'd35092,17'd36490,17'd36491,17'd31136,17'd17726,17'd14524,17'd16799,17'd29792,17'd31602,17'd33583,17'd36492,17'd36356,17'd33103,17'd36493,17'd29938,17'd11394,17'd26033,17'd34396,17'd31609,17'd29800,17'd29801,17'd29946,17'd36494,17'd36495,17'd36496,17'd36362,17'd36497,17'd36498,17'd36499,17'd36500,17'd36501,17'd36502,17'd36503,17'd36504,17'd36505,17'd36506,17'd36507,17'd36508,17'd36509,17'd36510,17'd36511,17'd34249,17'd35970,17'd36512,17'd36513,17'd36513,17'd36514,17'd36515,17'd36516,17'd36516,17'd36517,17'd35839,17'd35970,17'd35972,17'd35972,17'd35972,17'd35972,17'd36385,17'd36384,17'd36384,17'd36384,17'd35271,17'd35272,17'd36518,17'd35136,17'd35403,17'd36519,17'd35548,17'd36519,17'd36520,17'd35404,17'd35272,17'd36521,17'd36522,17'd36523,17'd34082,17'd36524,17'd36525,17'd36526,17'd36527,17'd36528,17'd36529,17'd36530,17'd36531,17'd36532,17'd36533,17'd35850,17'd35420,17'd35985,17'd36260,17'd35700,17'd35566,17'd35566,17'd36534,17'd36535,17'd34874,17'd36536,17'd36537,17'd36538,17'd36539,17'd36540,17'd36541,17'd36542,17'd27372,17'd29535,17'd27766,17'd25709,17'd28254,17'd24416,17'd23920,17'd36543,17'd22683,17'd36544,17'd36545,17'd22004,17'd31829,17'd22325,17'd30427,17'd22329,17'd31502,17'd23384,17'd23385,17'd24086,17'd28601,17'd25178,17'd25435,17'd25707,17'd27027,17'd29246,17'd30279,17'd27885,17'd32354,17'd32017,17'd29248,17'd29249,17'd36405,17'd36406,17'd32508,17'd29690,17'd36546,17'd29979,17'd34114,17'd36547,17'd36408,17'd36548,17'd31210,17'd36549,17'd36268,17'd36550,17'd36551,17'd36552,17'd36553,17'd36413,17'd24592,17'd23212,17'd30275,17'd25439,17'd24415,17'd24745,17'd25030,17'd25177,17'd24078,17'd27257,17'd27767,17'd25948,17'd36554,17'd26277,17'd36555,17'd36556,17'd36557,17'd36558,17'd36559,17'd36416,17'd30603,17'd36560,17'd25849,17'd25961,17'd27385,17'd28747,17'd26672,17'd36561,17'd36562,17'd36563,17'd23053,17'd31684,17'd28606,17'd30448,17'd29398,17'd36564,17'd30586,17'd27369,17'd27146,17'd28602,17'd33345,17'd36565,17'd23215,17'd36566,17'd36567,17'd36568,17'd36569,17'd36570,17'd36571,17'd36572,17'd36573,17'd36574,17'd36575,17'd36576,17'd36161,17'd21587,17'd36577,17'd36578,17'd5140,17'd36302,17'd36579,17'd36580,17'd36581,17'd36582,17'd36025,17'd36583,17'd36584,17'd36585,17'd24802,17'd18500,17'd19222,17'd36170,17'd29161,17'd11181,17'd27933,17'd10515,17'd8780,17'd8780,17'd27815,17'd29592,17'd10515,17'd28184,17'd6219,17'd30638,17'd28185,17'd33369,17'd36586,17'd7668,17'd7499,17'd6554,17'd5334,17'd5329,17'd25627,17'd31891,17'd9091,17'd28184,17'd10642,17'd28183,17'd27933,17'd27933,17'd10238,17'd6558,17'd36311,17'd36587,17'd36588,17'd35895,17'd35896,17'd36589,17'd36590,17'd36591,17'd36592,17'd36593,17'd36594,17'd36595,17'd36596,17'd36597,17'd36598,17'd36599,17'd36600,17'd6867,17'd795,17'd228,17'd1946,17'd6889,17'd8187,17'd7365,17'd4868,17'd6095,17'd36045,17'd6417,17'd6418,17'd8507,17'd36601,17'd33051,17'd31101,17'd31101,17'd31101,17'd31101,17'd31101,17'd31101,17'd27708,17'd29610,17'd36602,17'd34001,17'd6721,17'd14178,17'd6415,17'd5371,17'd445,17'd1962,17'd771,17'd224,17'd32405,17'd36603,17'd33377,17'd36604
},
'{
17'd4891,17'd3902,17'd4244,17'd27713,17'd3427,17'd2592,17'd3101,17'd3101,17'd3101,17'd3427,17'd3901,17'd15877,17'd15358,17'd2784,17'd1688,17'd1127,17'd2257,17'd2257,17'd1416,17'd18,17'd27,17'd285,17'd7061,17'd7061,17'd7225,17'd7225,17'd6599,17'd27445,17'd34004,17'd4581,17'd3912,17'd2608,17'd1706,17'd1707,17'd4095,17'd31732,17'd31732,17'd3600,17'd3436,17'd36605,17'd27829,17'd36606,17'd36607,17'd20137,17'd35773,17'd36608,17'd36609,17'd36610,17'd31917,17'd33549,17'd14893,17'd14768,17'd16033,17'd17690,17'd19255,17'd19128,17'd20292,17'd14470,17'd12954,17'd13092,17'd13092,17'd12357,17'd15763,17'd10941,17'd36329,17'd36611,17'd36612,17'd16172,17'd35627,17'd33553,17'd36191,17'd36466,17'd36613,17'd36614,17'd35072,17'd36615,17'd35216,17'd36616,17'd32111,17'd35359,17'd9583,17'd9309,17'd16042,17'd13612,17'd35631,17'd36057,17'd36617,17'd36472,17'd36194,17'd25126,17'd24980,17'd36473,17'd36473,17'd35631,17'd35500,17'd7107,17'd36618,17'd36619,17'd7273,17'd36620,17'd36621,17'd36622,17'd36342,17'd36476,17'd36623,17'd36624,17'd8723,17'd15684,17'd24361,17'd24039,17'd8566,17'd20176,17'd20176,17'd9348,17'd16795,17'd16067,17'd24043,17'd36070,17'd8252,17'd32121,17'd36625,17'd26153,17'd9344,17'd9740,17'd12584,17'd36626,17'd36627,17'd36628,17'd32919,17'd31287,17'd34037,17'd34037,17'd34203,17'd34381,17'd29646,17'd36629,17'd27121,17'd25925,17'd29488,17'd18326,17'd13369,17'd36630,17'd9043,17'd8720,17'd9194,17'd15684,17'd8720,17'd11810,17'd36631,17'd8099,17'd16691,17'd17016,17'd15056,17'd17353,17'd24213,17'd24368,17'd8885,17'd29334,17'd9042,17'd17480,17'd22645,17'd36208,17'd35232,17'd36632,17'd36633,17'd24031,17'd36634,17'd36635,17'd36636,17'd31441,17'd36637,17'd36638,17'd31763,17'd36211,17'd31447,17'd16327,17'd14672,17'd29205,17'd32294,17'd33249,17'd33583,17'd36356,17'd31141,17'd35654,17'd33251,17'd36357,17'd24854,17'd36639,17'd29669,17'd29216,17'd31149,17'd36640,17'd36360,17'd36641,17'd34570,17'd36642,17'd36643,17'd36644,17'd36645,17'd36646,17'd36647,17'd36648,17'd36649,17'd36650,17'd36651,17'd36652,17'd36653,17'd36654,17'd36655,17'd36656,17'd36657,17'd36658,17'd36659,17'd36660,17'd36661,17'd36514,17'd36662,17'd36663,17'd36664,17'd36665,17'd36666,17'd36667,17'd36668,17'd36668,17'd36669,17'd36670,17'd36384,17'd35972,17'd35972,17'd35972,17'd35972,17'd36385,17'd36671,17'd35550,17'd36387,17'd36386,17'd35136,17'd35402,17'd35135,17'd35134,17'd35403,17'd35133,17'd36672,17'd36672,17'd36522,17'd36673,17'd36674,17'd36675,17'd36676,17'd36677,17'd36678,17'd36679,17'd36680,17'd36681,17'd36531,17'd36682,17'd36121,17'd36122,17'd35420,17'd35285,17'd36683,17'd35700,17'd35422,17'd35422,17'd36684,17'd36685,17'd36535,17'd36536,17'd36686,17'd36687,17'd36688,17'd36689,17'd35291,17'd36690,17'd34637,17'd27146,17'd26174,17'd28597,17'd27637,17'd28851,17'd23733,17'd29974,17'd22334,17'd36691,17'd36692,17'd22166,17'd32345,17'd34111,17'd30426,17'd22329,17'd23736,17'd34137,17'd23386,17'd23733,17'd28975,17'd25178,17'd28600,17'd25833,17'd26902,17'd29245,17'd31503,17'd27885,17'd28134,17'd32355,17'd33486,17'd29249,17'd29249,17'd29249,17'd34285,17'd29690,17'd30884,17'd29979,17'd34285,17'd36547,17'd30589,17'd36693,17'd36694,17'd30149,17'd29116,17'd36695,17'd36696,17'd36697,17'd36698,17'd36699,17'd36700,17'd29376,17'd30275,17'd36701,17'd24415,17'd28851,17'd25030,17'd25177,17'd24078,17'd33342,17'd30606,17'd25948,17'd36702,17'd25826,17'd32356,17'd28859,17'd36703,17'd36704,17'd36705,17'd36558,17'd36706,17'd30758,17'd31854,17'd36707,17'd25448,17'd24432,17'd36708,17'd36147,17'd36709,17'd36710,17'd36711,17'd36712,17'd29399,17'd36713,17'd36714,17'd36715,17'd36008,17'd35426,17'd36542,17'd26174,17'd36716,17'd30126,17'd23567,17'd22677,17'd36717,17'd36718,17'd36719,17'd36720,17'd36721,17'd36722,17'd36723,17'd36724,17'd36725,17'd36726,17'd36727,17'd30178,17'd36728,17'd36729,17'd3829,17'd36302,17'd5321,17'd36730,17'd36731,17'd36168,17'd36732,17'd36583,17'd36442,17'd36733,17'd17905,17'd18500,17'd18970,17'd36734,17'd36735,17'd28305,17'd27933,17'd27933,17'd9933,17'd9933,17'd9933,17'd27815,17'd10515,17'd10514,17'd6220,17'd30638,17'd30638,17'd30333,17'd6554,17'd7499,17'd7499,17'd6554,17'd5335,17'd5330,17'd25627,17'd30638,17'd6390,17'd8780,17'd28183,17'd30933,17'd27933,17'd28183,17'd10238,17'd6558,17'd8630,17'd36736,17'd36588,17'd36737,17'd36034,17'd36738,17'd36590,17'd36739,17'd36740,17'd36741,17'd36742,17'd36743,17'd36744,17'd36745,17'd36746,17'd36747,17'd36322,17'd36748,17'd628,17'd446,17'd4423,17'd6889,17'd6581,17'd4869,17'd4868,17'd6095,17'd36045,17'd6417,17'd6418,17'd8507,17'd36601,17'd33051,17'd31729,17'd31101,17'd31101,17'd31101,17'd31101,17'd31101,17'd31101,17'd31101,17'd27949,17'd33050,17'd5631,17'd14178,17'd5372,17'd5371,17'd445,17'd2249,17'd1959,17'd224,17'd766,17'd36749,17'd36750,17'd36604
},
'{
17'd3902,17'd3902,17'd4243,17'd27951,17'd15746,17'd4887,17'd2784,17'd3101,17'd2934,17'd3751,17'd3592,17'd15877,17'd15358,17'd14070,17'd1688,17'd1127,17'd1414,17'd1416,17'd17,17'd18,17'd27,17'd286,17'd7555,17'd7555,17'd7386,17'd6599,17'd26971,17'd26731,17'd34004,17'd4581,17'd3912,17'd2608,17'd3598,17'd4258,17'd2609,17'd2609,17'd2435,17'd1708,17'd3436,17'd36751,17'd3765,17'd13192,17'd36752,17'd4109,17'd36753,17'd36754,17'd36755,17'd34937,17'd15385,17'd32739,17'd14767,17'd14768,17'd16033,17'd27833,17'd36756,17'd19128,17'd16765,17'd14621,17'd13092,17'd12357,17'd14469,17'd12357,17'd11762,17'd36757,17'd36189,17'd36053,17'd36758,17'd36759,17'd36760,17'd34525,17'd36191,17'd36192,17'd36761,17'd36762,17'd35781,17'd35358,17'd35499,17'd32424,17'd14639,17'd18306,17'd9849,17'd9309,17'd13611,17'd7921,17'd25126,17'd36617,17'd36763,17'd36472,17'd36194,17'd25126,17'd24980,17'd24980,17'd36764,17'd25126,17'd36336,17'd7107,17'd36765,17'd36766,17'd36767,17'd36768,17'd36769,17'd36770,17'd36771,17'd36772,17'd36773,17'd36774,17'd8728,17'd29920,17'd29637,17'd8566,17'd12118,17'd17237,17'd8410,17'd9046,17'd17231,17'd26038,17'd12867,17'd36775,17'd12867,17'd8571,17'd17607,17'd10336,17'd17716,17'd11277,17'd11669,17'd25143,17'd36776,17'd32760,17'd33718,17'd31442,17'd31442,17'd31442,17'd31288,17'd34704,17'd36777,17'd29480,17'd26629,17'd25671,17'd23167,17'd11669,17'd10169,17'd23679,17'd9189,17'd8720,17'd8873,17'd8721,17'd15297,17'd8726,17'd9349,17'd12588,17'd17353,17'd16691,17'd8581,17'd19780,17'd21987,17'd8572,17'd8886,17'd17607,17'd10175,17'd26153,17'd36778,17'd34695,17'd36779,17'd36780,17'd24363,17'd28817,17'd29642,17'd36781,17'd36782,17'd34545,17'd34380,17'd31941,17'd29482,17'd28466,17'd36783,17'd28232,17'd16915,17'd30983,17'd36784,17'd36785,17'd32939,17'd31451,17'd36786,17'd36787,17'd29634,17'd36788,17'd35936,17'd34396,17'd29501,17'd30994,17'd36789,17'd36790,17'd36791,17'd36792,17'd36793,17'd36497,17'd36794,17'd36795,17'd36796,17'd36797,17'd36798,17'd36799,17'd36800,17'd36801,17'd36802,17'd36803,17'd36804,17'd36805,17'd36806,17'd36807,17'd36808,17'd36809,17'd36810,17'd36811,17'd36243,17'd36512,17'd36812,17'd36813,17'd36814,17'd36814,17'd36515,17'd36815,17'd36816,17'd36664,17'd36817,17'd36818,17'd36819,17'd36820,17'd36383,17'd36105,17'd36105,17'd36383,17'd36383,17'd36383,17'd36105,17'd35838,17'd36108,17'd36108,17'd36821,17'd35135,17'd36822,17'd36823,17'd35135,17'd35271,17'd36824,17'd34424,17'd36825,17'd36524,17'd33453,17'd36826,17'd36827,17'd36828,17'd36829,17'd36830,17'd36831,17'd36832,17'd36833,17'd36121,17'd35565,17'd36834,17'd36835,17'd36836,17'd35700,17'd36837,17'd36838,17'd36839,17'd36840,17'd34874,17'd36841,17'd36842,17'd36843,17'd36842,17'd34877,17'd33791,17'd34637,17'd27146,17'd26174,17'd28598,17'd27512,17'd24416,17'd31033,17'd29829,17'd22330,17'd30580,17'd36844,17'd22164,17'd36845,17'd36846,17'd23573,17'd32827,17'd30579,17'd23923,17'd29975,17'd29376,17'd28849,17'd25032,17'd25317,17'd25565,17'd28853,17'd31035,17'd31353,17'd31354,17'd32354,17'd32193,17'd36847,17'd33166,17'd29249,17'd28728,17'd36848,17'd29536,17'd29536,17'd29831,17'd34114,17'd35712,17'd36849,17'd36850,17'd36851,17'd36852,17'd36853,17'd36854,17'd29843,17'd36550,17'd36855,17'd36856,17'd35999,17'd29242,17'd29242,17'd29241,17'd23917,17'd28851,17'd25030,17'd28717,17'd28599,17'd27513,17'd30734,17'd26903,17'd25698,17'd26277,17'd36857,17'd36858,17'd36859,17'd36703,17'd36860,17'd36861,17'd34130,17'd36862,17'd30146,17'd28384,17'd32205,17'd27159,17'd24916,17'd35173,17'd36863,17'd36864,17'd32529,17'd34890,17'd36865,17'd36866,17'd33658,17'd33808,17'd36867,17'd36868,17'd27516,17'd36869,17'd28723,17'd29976,17'd23211,17'd36870,17'd30727,17'd36871,17'd24749,17'd36872,17'd36873,17'd36874,17'd36875,17'd36876,17'd36877,17'd36878,17'd22233,17'd36879,17'd36880,17'd36881,17'd36882,17'd35190,17'd9213,17'd10195,17'd36883,17'd36884,17'd36885,17'd36583,17'd36733,17'd36443,17'd24802,17'd18500,17'd19222,17'd36734,17'd36886,17'd28183,17'd27933,17'd28057,17'd29592,17'd9933,17'd27815,17'd27815,17'd27815,17'd10515,17'd7668,17'd33369,17'd5004,17'd25627,17'd5160,17'd5614,17'd6220,17'd6390,17'd5160,17'd5160,17'd5008,17'd5164,17'd36887,17'd7669,17'd30933,17'd36888,17'd31551,17'd10515,17'd6555,17'd5920,17'd8473,17'd36889,17'd36890,17'd36737,17'd36891,17'd36892,17'd36893,17'd36894,17'd36895,17'd36896,17'd36897,17'd36898,17'd36899,17'd36900,17'd36901,17'd22099,17'd36181,17'd36902,17'd1121,17'd625,17'd4085,17'd6889,17'd6889,17'd5630,17'd4713,17'd4713,17'd4868,17'd6258,17'd7537,17'd8507,17'd11336,17'd11061,17'd36903,17'd36904,17'd36905,17'd36905,17'd36905,17'd36905,17'd36906,17'd36905,17'd35487,17'd11061,17'd4714,17'd3073,17'd5372,17'd5050,17'd2559,17'd953,17'd771,17'd224,17'd36907,17'd36603,17'd36908,17'd36909
},
'{
17'd3902,17'd3902,17'd4243,17'd27951,17'd15746,17'd7545,17'd2784,17'd2934,17'd3751,17'd3751,17'd3592,17'd15877,17'd15358,17'd3252,17'd1688,17'd1127,17'd1416,17'd1416,17'd17,17'd16,17'd28,17'd286,17'd7555,17'd7555,17'd7386,17'd7225,17'd5972,17'd12931,17'd32729,17'd4432,17'd3912,17'd2608,17'd3598,17'd2435,17'd2609,17'd35620,17'd1842,17'd1561,17'd3266,17'd36910,17'd36911,17'd26131,17'd20578,17'd36912,17'd36913,17'd36914,17'd36915,17'd34521,17'd15385,17'd32739,17'd14767,17'd14768,17'd16033,17'd27833,17'd36756,17'd19128,17'd16765,17'd13211,17'd13092,17'd14469,17'd14763,17'd12357,17'd10687,17'd36916,17'd36917,17'd16292,17'd36918,17'd35355,17'd34944,17'd33553,17'd36191,17'd36332,17'd36333,17'd36762,17'd35781,17'd35358,17'd33706,17'd35074,17'd16665,17'd14230,17'd9849,17'd11631,17'd8701,17'd25514,17'd36194,17'd36763,17'd36919,17'd36920,17'd36921,17'd36922,17'd36923,17'd36764,17'd25126,17'd36057,17'd36924,17'd35921,17'd36925,17'd36926,17'd36927,17'd36928,17'd36929,17'd36770,17'd36771,17'd36930,17'd36931,17'd36932,17'd8728,17'd23861,17'd24999,17'd8881,17'd12118,17'd8724,17'd15429,17'd8729,17'd23860,17'd23861,17'd12867,17'd23685,17'd18808,17'd8724,17'd9194,17'd17480,17'd17716,17'd19531,17'd28463,17'd20608,17'd32759,17'd32918,17'd33567,17'd31442,17'd32920,17'd32920,17'd34203,17'd31773,17'd36777,17'd28460,17'd25927,17'd30229,17'd17478,17'd19280,17'd10992,17'd9339,17'd9043,17'd8720,17'd8875,17'd9348,17'd8725,17'd15429,17'd24213,17'd12588,17'd25680,17'd25680,17'd9888,17'd8579,17'd21987,17'd8572,17'd8886,17'd16317,17'd10336,17'd16552,17'd36778,17'd34695,17'd36933,17'd36934,17'd26035,17'd36935,17'd31295,17'd33575,17'd34047,17'd36936,17'd33568,17'd36937,17'd29201,17'd28465,17'd36783,17'd28232,17'd17015,17'd30086,17'd33249,17'd36785,17'd33102,17'd31451,17'd33251,17'd36079,17'd11273,17'd27001,17'd31783,17'd36938,17'd29350,17'd36939,17'd36940,17'd36941,17'd30696,17'd33262,17'd31796,17'd36942,17'd36943,17'd36944,17'd36945,17'd36946,17'd36947,17'd36948,17'd36949,17'd36950,17'd36951,17'd36952,17'd36953,17'd36954,17'd36955,17'd36956,17'd36957,17'd36958,17'd36959,17'd36960,17'd36819,17'd36817,17'd36961,17'd36961,17'd36962,17'd36962,17'd36961,17'd36664,17'd36815,17'd36515,17'd36819,17'd36963,17'd36817,17'd36963,17'd36964,17'd36383,17'd36105,17'd36105,17'd36105,17'd35683,17'd36105,17'd35683,17'd36965,17'd35273,17'd36247,17'd36966,17'd36967,17'd36967,17'd36108,17'd36521,17'd36824,17'd36968,17'd36969,17'd36970,17'd35137,17'd36971,17'd36972,17'd36973,17'd36974,17'd36975,17'd36976,17'd36832,17'd36832,17'd36121,17'd35565,17'd36977,17'd36978,17'd36836,17'd35700,17'd36979,17'd36980,17'd36981,17'd36839,17'd35148,17'd36982,17'd36842,17'd36843,17'd36687,17'd36983,17'd33941,17'd30735,17'd33163,17'd26903,17'd27513,17'd25568,17'd24745,17'd23917,17'd29530,17'd22329,17'd31343,17'd32497,17'd36984,17'd36845,17'd36985,17'd23573,17'd36986,17'd29974,17'd23388,17'd36987,17'd23566,17'd23384,17'd28977,17'd25317,17'd25708,17'd28853,17'd31035,17'd31353,17'd31354,17'd32192,17'd36988,17'd36847,17'd33166,17'd28857,17'd28728,17'd29537,17'd29537,17'd28857,17'd29831,17'd36989,17'd28982,17'd36990,17'd27516,17'd36991,17'd36992,17'd36993,17'd36994,17'd36995,17'd36695,17'd36996,17'd36997,17'd36701,17'd25033,17'd34137,17'd29528,17'd23917,17'd28851,17'd28254,17'd28717,17'd31055,17'd27513,17'd28599,17'd25833,17'd26167,17'd29379,17'd36998,17'd36999,17'd37000,17'd37001,17'd35867,17'd37002,17'd34897,17'd30743,17'd37003,17'd29987,17'd26302,17'd30295,17'd24915,17'd37004,17'd37005,17'd37006,17'd32840,17'd37007,17'd37008,17'd36282,17'd29128,17'd28022,17'd31362,17'd37009,17'd36868,17'd37010,17'd27766,17'd29103,17'd23919,17'd37011,17'd22157,17'd37012,17'd37013,17'd37014,17'd37015,17'd37016,17'd37017,17'd37018,17'd37019,17'd19691,17'd22075,17'd37020,17'd37021,17'd37022,17'd5907,17'd35190,17'd35467,17'd37023,17'd37024,17'd37025,17'd36732,17'd37026,17'd37027,17'd37027,17'd24654,17'd18375,17'd19222,17'd22943,17'd35477,17'd34922,17'd28057,17'd28183,17'd29592,17'd29592,17'd27815,17'd28184,17'd27815,17'd10515,17'd27696,17'd37028,17'd30637,17'd5002,17'd5329,17'd5336,17'd5919,17'd6390,17'd30638,17'd5160,17'd37029,17'd5008,17'd37030,17'd7669,17'd30933,17'd36888,17'd31551,17'd10515,17'd37031,17'd36311,17'd8474,17'd37032,17'd36890,17'd37033,17'd37034,17'd36892,17'd36448,17'd37035,17'd37036,17'd37037,17'd37038,17'd37039,17'd37040,17'd37041,17'd36901,17'd37042,17'd23300,17'd37043,17'd235,17'd626,17'd4085,17'd3073,17'd3073,17'd5630,17'd4713,17'd4713,17'd4868,17'd6258,17'd7537,17'd8507,17'd11336,17'd11061,17'd36903,17'd36903,17'd36905,17'd36905,17'd36905,17'd36905,17'd36906,17'd36905,17'd35487,17'd34002,17'd11335,17'd9123,17'd8185,17'd4880,17'd2392,17'd2249,17'd1959,17'd224,17'd36907,17'd37044,17'd37045,17'd37046
},
'{
17'd4244,17'd4243,17'd27951,17'd15876,17'd13428,17'd7545,17'd2935,17'd3101,17'd3427,17'd3751,17'd3592,17'd35619,17'd37047,17'd3252,17'd1689,17'd1127,17'd1416,17'd1416,17'd17,17'd18,17'd27,17'd286,17'd7555,17'd7555,17'd7386,17'd6599,17'd26971,17'd12931,17'd4741,17'd4253,17'd3912,17'd4433,17'd4258,17'd2435,17'd2609,17'd35620,17'd1842,17'd3439,17'd24674,17'd36910,17'd12934,17'd37048,17'd37049,17'd37050,17'd37051,17'd37052,17'd37053,17'd34521,17'd15385,17'd32739,17'd14767,17'd16768,17'd17448,17'd19255,17'd19007,17'd20292,17'd14622,17'd13093,17'd13092,17'd14469,17'd12062,17'd12062,17'd10687,17'd37054,17'd14224,17'd14771,17'd36759,17'd15526,17'd33065,17'd34184,17'd33861,17'd36467,17'd36333,17'd37055,17'd35781,17'd35358,17'd33228,17'd32111,17'd35359,17'd13104,17'd9849,17'd9016,17'd8701,17'd25514,17'd37056,17'd37057,17'd37058,17'd36763,17'd37056,17'd25126,17'd36764,17'd36764,17'd25126,17'd36057,17'd36924,17'd35921,17'd37059,17'd37060,17'd7274,17'd36928,17'd37061,17'd36770,17'd37062,17'd37063,17'd37064,17'd10858,17'd8728,17'd9046,17'd9040,17'd8882,17'd12118,17'd12118,17'd9482,17'd8569,17'd25531,17'd9046,17'd8100,17'd13004,17'd9349,17'd9046,17'd15684,17'd10174,17'd14674,17'd11277,17'd11275,17'd21362,17'd29327,17'd37065,17'd32283,17'd31442,17'd32920,17'd32920,17'd34203,17'd36937,17'd29645,17'd28460,17'd24856,17'd15055,17'd11397,17'd22820,17'd11136,17'd9191,17'd9043,17'd9041,17'd16067,17'd15297,17'd8410,17'd9744,17'd24213,17'd12426,17'd25680,17'd25680,17'd8580,17'd19923,17'd17481,17'd15429,17'd8886,17'd16317,17'd17480,17'd16552,17'd27988,17'd35932,17'd37066,17'd37067,17'd37068,17'd28103,17'd37069,17'd33575,17'd33882,17'd33243,17'd31773,17'd29646,17'd28945,17'd28348,17'd27235,17'd17726,17'd29205,17'd30087,17'd37070,17'd37071,17'd32773,17'd36493,17'd35242,17'd35655,17'd36788,17'd35936,17'd37072,17'd29500,17'd30994,17'd37073,17'd37074,17'd36641,17'd37075,17'd34569,17'd37076,17'd35528,17'd37077,17'd37078,17'd37079,17'd37080,17'd37081,17'd37082,17'd37083,17'd37084,17'd37085,17'd37086,17'd37087,17'd37088,17'd37089,17'd37090,17'd37091,17'd37091,17'd36108,17'd35970,17'd35839,17'd36964,17'd36661,17'd37092,17'd37093,17'd37094,17'd37094,17'd37094,17'd37095,17'd37096,17'd36819,17'd36668,17'd36963,17'd36963,17'd36668,17'd37097,17'd36820,17'd36243,17'd36383,17'd35839,17'd36105,17'd36243,17'd35683,17'd35838,17'd36821,17'd35135,17'd37098,17'd36967,17'd36108,17'd36107,17'd37099,17'd37100,17'd35678,17'd35137,17'd37101,17'd37102,17'd37103,17'd37104,17'd37105,17'd36118,17'd37106,17'd37107,17'd37108,17'd37109,17'd35565,17'd36977,17'd36978,17'd36836,17'd35986,17'd36979,17'd37110,17'd37111,17'd37112,17'd35286,17'd36982,17'd36843,17'd36843,17'd37113,17'd37114,17'd32005,17'd34637,17'd34637,17'd28853,17'd26064,17'd25568,17'd24895,17'd24249,17'd29376,17'd22501,17'd30426,17'd22157,17'd22163,17'd36845,17'd37115,17'd23573,17'd36986,17'd37116,17'd23569,17'd37117,17'd29686,17'd29242,17'd30126,17'd28369,17'd27766,17'd28853,17'd30586,17'd35426,17'd31503,17'd32354,17'd32193,17'd37118,17'd33166,17'd28857,17'd28857,17'd29537,17'd29537,17'd28857,17'd29536,17'd36989,17'd28982,17'd32832,17'd30735,17'd37119,17'd25835,17'd37120,17'd37121,17'd37122,17'd37123,17'd36996,17'd37124,17'd36565,17'd35021,17'd34137,17'd29528,17'd23917,17'd28851,17'd28254,17'd28717,17'd31055,17'd30734,17'd31055,17'd26174,17'd26279,17'd29379,17'd37125,17'd36858,17'd37126,17'd37001,17'd35867,17'd35168,17'd37127,17'd30743,17'd37003,17'd30146,17'd26189,17'd25453,17'd25049,17'd37128,17'd37129,17'd37130,17'd37131,17'd37132,17'd37133,17'd35315,17'd37134,17'd28022,17'd29542,17'd30594,17'd37135,17'd34480,17'd25833,17'd29101,17'd30431,17'd32008,17'd22158,17'd35737,17'd24906,17'd37136,17'd37137,17'd37138,17'd37139,17'd37140,17'd37141,17'd37142,17'd21914,17'd37143,17'd37144,17'd37145,17'd10357,17'd37146,17'd37147,17'd5141,17'd36304,17'd36440,17'd36025,17'd37148,17'd37149,17'd37150,17'd18135,17'd20115,17'd19480,17'd19087,17'd36170,17'd37151,17'd30488,17'd28305,17'd29592,17'd27815,17'd28184,17'd28184,17'd27815,17'd10515,17'd9933,17'd37152,17'd32553,17'd30637,17'd5004,17'd5335,17'd5919,17'd5615,17'd5335,17'd5160,17'd29024,17'd37153,17'd5009,17'd6222,17'd27933,17'd31243,17'd28183,17'd37154,17'd37155,17'd36311,17'd8474,17'd37032,17'd37156,17'd37157,17'd37158,17'd36892,17'd37159,17'd37160,17'd37161,17'd37162,17'd37163,17'd37039,17'd37164,17'd37165,17'd37166,17'd37042,17'd36454,17'd37167,17'd630,17'd623,17'd3391,17'd5958,17'd3073,17'd5630,17'd4729,17'd4713,17'd4868,17'd6258,17'd6418,17'd8507,17'd11336,17'd11061,17'd35487,17'd36903,17'd36905,17'd36905,17'd37168,17'd36905,17'd36905,17'd36905,17'd35487,17'd11061,17'd4714,17'd3073,17'd5372,17'd5050,17'd2417,17'd953,17'd771,17'd224,17'd36907,17'd31104,17'd37169,17'd37170
},
'{
17'd4244,17'd3902,17'd4243,17'd25384,17'd14743,17'd5508,17'd2935,17'd2934,17'd3901,17'd3901,17'd3592,17'd15877,17'd15358,17'd3252,17'd1689,17'd1127,17'd1416,17'd1416,17'd17,17'd18,17'd27,17'd286,17'd7385,17'd7385,17'd7386,17'd6745,17'd5972,17'd26469,17'd4741,17'd4253,17'd3261,17'd37171,17'd24967,17'd2435,17'd35620,17'd35620,17'd1561,17'd3437,17'd32731,17'd27829,17'd37172,17'd37173,17'd5070,17'd4110,17'd3454,17'd37174,17'd37175,17'd34521,17'd15385,17'd32739,17'd14768,17'd16033,17'd17445,17'd19255,17'd17689,17'd28667,17'd14622,17'd35352,17'd14469,17'd16284,17'd12062,17'd11625,17'd10424,17'd37176,17'd37177,17'd37178,17'd37179,17'd34943,17'd37180,17'd37181,17'd33861,17'd36613,17'd37182,17'd36762,17'd37183,17'd35358,17'd33864,17'd15399,17'd14230,17'd9707,17'd9309,17'd16042,17'd13612,17'd25126,17'd36471,17'd37057,17'd37184,17'd36919,17'd36617,17'd37056,17'd25126,17'd37185,17'd37186,17'd37187,17'd36924,17'd36059,17'd7271,17'd37188,17'd37189,17'd37190,17'd37191,17'd37192,17'd37193,17'd37194,17'd37195,17'd36932,17'd8728,17'd9046,17'd9348,17'd8882,17'd17237,17'd8725,17'd9482,17'd8886,17'd17123,17'd8886,17'd12724,17'd13139,17'd8413,17'd9046,17'd15684,17'd10335,17'd14674,17'd17718,17'd37196,17'd23170,17'd33402,17'd37065,17'd32283,17'd31442,17'd32920,17'd32920,17'd33568,17'd36491,17'd31286,17'd28343,17'd26149,17'd29488,17'd11668,17'd17842,17'd13255,17'd9190,17'd9042,17'd9041,17'd9040,17'd8726,17'd9744,17'd11967,17'd13257,17'd12426,17'd25680,17'd25680,17'd10028,17'd8578,17'd17481,17'd8412,17'd8886,17'd26498,17'd26153,17'd17728,17'd37197,17'd37198,17'd37199,17'd37200,17'd37201,17'd37202,17'd37203,17'd33575,17'd33096,17'd31591,17'd37204,17'd37205,17'd28572,17'd37206,17'd27235,17'd16327,17'd29340,17'd31140,17'd32448,17'd31778,17'd31603,17'd34214,17'd37207,17'd35655,17'd29939,17'd29796,17'd37208,17'd37209,17'd28959,17'd30102,17'd37210,17'd37211,17'd31467,17'd35528,17'd31004,17'd37212,17'd37213,17'd37214,17'd37215,17'd31978,17'd37216,17'd37217,17'd37218,17'd37219,17'd37220,17'd37221,17'd37222,17'd37223,17'd37224,17'd35961,17'd36103,17'd37225,17'd36383,17'd37226,17'd37226,17'd36668,17'd37227,17'd37228,17'd36661,17'd37092,17'd37229,17'd37093,17'd37230,17'd37231,17'd37095,17'd36963,17'd36819,17'd36819,17'd36668,17'd36963,17'd36819,17'd36660,17'd37226,17'd36105,17'd36105,17'd36383,17'd35683,17'd35970,17'd35838,17'd36821,17'd35135,17'd36518,17'd35964,17'd35964,17'd37232,17'd37233,17'd35678,17'd37234,17'd37235,17'd33923,17'd37236,17'd37237,17'd37238,17'd37239,17'd37240,17'd36531,17'd37241,17'd37109,17'd35565,17'd36977,17'd36978,17'd37242,17'd35986,17'd37243,17'd37244,17'd37245,17'd37246,17'd35286,17'd36982,17'd36843,17'd37247,17'd37113,17'd37248,17'd33790,17'd31035,17'd34637,17'd27146,17'd28602,17'd28717,17'd25030,17'd23916,17'd29376,17'd33158,17'd23573,17'd22158,17'd32497,17'd37249,17'd36131,17'd23573,17'd36986,17'd36543,17'd23569,17'd37117,17'd29975,17'd23385,17'd32659,17'd25438,17'd28602,17'd28725,17'd28486,17'd31352,17'd31503,17'd32354,17'd32193,17'd37118,17'd33166,17'd28857,17'd28857,17'd29537,17'd28728,17'd28857,17'd29536,17'd36989,17'd37250,17'd32832,17'd30735,17'd37251,17'd33008,17'd37252,17'd37121,17'd37253,17'd31046,17'd37254,17'd37255,17'd30731,17'd37256,17'd23384,17'd31033,17'd23917,17'd28851,17'd28254,17'd28717,17'd31055,17'd30734,17'd31055,17'd26174,17'd26279,17'd29246,17'd37125,17'd36999,17'd37257,17'd29984,17'd36002,17'd36557,17'd35168,17'd37127,17'd37258,17'd30438,17'd25848,17'd26188,17'd25191,17'd29389,17'd37259,17'd37260,17'd37261,17'd37262,17'd37263,17'd31357,17'd37264,17'd28022,17'd33005,17'd33327,17'd37265,17'd27517,17'd37266,17'd29970,17'd37267,17'd34452,17'd23573,17'd37268,17'd37269,17'd37270,17'd37271,17'd37272,17'd37273,17'd37274,17'd37275,17'd37276,17'd23779,17'd22729,17'd37277,17'd37278,17'd37279,17'd37280,17'd6206,17'd33038,17'd37281,17'd37282,17'd37283,17'd37284,17'd37285,17'd37285,17'd18261,17'd18852,17'd19222,17'd22767,17'd37286,17'd37287,17'd36735,17'd28534,17'd27933,17'd29592,17'd27815,17'd28184,17'd27815,17'd10515,17'd9933,17'd32073,17'd31553,17'd5004,17'd30637,17'd30333,17'd6219,17'd6219,17'd28185,17'd25627,17'd37153,17'd4685,17'd37288,17'd6708,17'd29592,17'd31243,17'd28183,17'd10514,17'd37289,17'd35197,17'd37290,17'd37291,17'd37156,17'd37292,17'd37293,17'd37294,17'd37295,17'd37296,17'd37297,17'd37298,17'd37299,17'd37300,17'd37301,17'd37302,17'd37303,17'd37042,17'd36599,17'd36455,17'd242,17'd2587,17'd2586,17'd4882,17'd5940,17'd4729,17'd4729,17'd4713,17'd4868,17'd6095,17'd6418,17'd6417,17'd7537,17'd11061,17'd35487,17'd36903,17'd36905,17'd37168,17'd37168,17'd36905,17'd36905,17'd36905,17'd35487,17'd11061,17'd4714,17'd3073,17'd5372,17'd4880,17'd1261,17'd623,17'd1961,17'd29891,17'd36907,17'd36603,17'd37304,17'd37305
},
'{
17'd4244,17'd4243,17'd27951,17'd25384,17'd14743,17'd4246,17'd2935,17'd3101,17'd3428,17'd3901,17'd3592,17'd35619,17'd34512,17'd3252,17'd1689,17'd1127,17'd1416,17'd1416,17'd3905,17'd18,17'd27,17'd286,17'd7385,17'd7385,17'd6745,17'd7062,17'd26846,17'd26469,17'd4581,17'd4252,17'd3261,17'd4583,17'd4257,17'd2435,17'd35620,17'd35620,17'd1561,17'd3266,17'd37306,17'd27829,17'd37307,17'd37308,17'd20137,17'd37309,17'd37310,17'd37311,17'd36462,17'd32098,17'd15008,17'd14767,17'd16768,17'd16033,17'd17320,17'd17206,17'd17204,17'd12361,17'd14890,17'd12678,17'd14469,17'd16284,17'd11762,17'd11625,17'd37312,17'd37313,17'd16524,17'd37314,17'd37315,17'd33553,17'd37316,17'd37181,17'd33861,17'd37317,17'd36333,17'd37318,17'd37319,17'd35358,17'd32424,17'd35784,17'd14230,17'd14109,17'd11631,17'd13733,17'd36473,17'd36057,17'd36763,17'd37320,17'd37184,17'd36763,17'd37321,17'd37322,17'd7103,17'd7103,17'd37323,17'd37187,17'd37324,17'd36337,17'd37325,17'd37326,17'd37327,17'd37328,17'd37329,17'd37330,17'd37331,17'd37332,17'd37333,17'd37334,17'd8728,17'd9046,17'd8886,17'd10027,17'd8569,17'd8725,17'd8410,17'd9195,17'd17123,17'd8886,17'd18808,17'd8100,17'd11137,17'd8877,17'd9189,17'd10335,17'd15807,17'd11671,17'd24029,17'd24209,17'd32591,17'd32919,17'd31287,17'd33875,17'd34037,17'd31288,17'd34381,17'd37335,17'd35372,17'd28104,17'd25671,17'd14259,17'd28463,17'd10168,17'd10857,17'd9191,17'd9189,17'd9194,17'd9040,17'd11403,17'd15568,17'd9349,17'd21208,17'd12426,17'd9888,17'd8580,17'd19923,17'd8578,17'd17481,17'd8410,17'd9041,17'd17480,17'd16552,17'd37336,17'd37337,17'd37338,17'd37339,17'd37340,17'd37341,17'd33092,17'd33727,17'd33730,17'd33093,17'd32597,17'd37205,17'd34390,17'd29336,17'd37206,17'd28233,17'd13642,17'd30087,17'd33250,17'd31603,17'd33578,17'd37342,17'd33886,17'd35242,17'd10730,17'd10845,17'd34051,17'd37343,17'd29665,17'd37344,17'd37345,17'd36495,17'd37346,17'd36643,17'd37347,17'd35528,17'd37348,17'd37349,17'd37350,17'd37351,17'd37352,17'd37353,17'd37354,17'd37355,17'd37356,17'd37357,17'd37358,17'd37359,17'd37360,17'd35833,17'd37231,17'd37361,17'd37362,17'd37363,17'd37362,17'd37363,17'd37230,17'd37363,17'd37231,17'd37364,17'd37364,17'd37364,17'd37364,17'd37365,17'd37231,17'd37363,17'd37363,17'd37230,17'd37096,17'd37366,17'd37367,17'd37368,17'd37368,17'd36820,17'd36243,17'd36383,17'd36105,17'd35683,17'd36105,17'd35839,17'd35838,17'd35272,17'd36386,17'd34077,17'd34077,17'd35135,17'd37369,17'd36969,17'd37370,17'd34076,17'd37371,17'd37372,17'd37373,17'd37374,17'd37375,17'd37376,17'd37377,17'd37378,17'd36682,17'd37379,17'd37380,17'd37381,17'd36683,17'd36260,17'd37382,17'd37244,17'd37245,17'd37383,17'd36398,17'd36686,17'd36843,17'd37384,17'd37247,17'd35567,17'd33790,17'd31035,17'd30735,17'd27372,17'd27766,17'd28717,17'd29976,17'd23916,17'd34137,17'd32008,17'd22332,17'd22161,17'd30580,17'd37385,17'd22505,17'd22677,17'd22329,17'd36543,17'd29974,17'd23217,17'd37386,17'd29687,17'd23916,17'd25177,17'd28602,17'd28725,17'd30586,17'd32016,17'd31503,17'd32354,17'd32193,17'd33656,17'd29249,17'd28857,17'd28857,17'd29536,17'd28857,17'd28857,17'd29536,17'd29831,17'd28728,17'd27885,17'd30735,17'd32995,17'd28717,17'd37387,17'd30446,17'd24089,17'd37388,17'd37389,17'd37390,17'd35159,17'd28722,17'd29689,17'd23732,17'd23917,17'd28851,17'd27637,17'd25709,17'd28597,17'd28598,17'd31055,17'd25833,17'd26279,17'd29246,17'd37125,17'd36849,17'd36858,17'd37391,17'd37392,17'd36002,17'd37393,17'd37127,17'd37258,17'd37394,17'd37395,17'd37396,17'd25453,17'd37397,17'd37398,17'd37399,17'd37400,17'd37401,17'd37402,17'd37403,17'd32213,17'd37404,17'd29705,17'd28382,17'd28610,17'd37405,17'd37406,17'd26402,17'd31360,17'd37407,17'd34278,17'd37408,17'd37409,17'd37410,17'd37411,17'd37412,17'd37413,17'd37414,17'd36015,17'd37415,17'd20500,17'd37416,17'd37417,17'd37418,17'd37419,17'd37420,17'd9499,17'd37421,17'd37422,17'd37423,17'd37424,17'd37425,17'd37426,17'd37426,17'd18135,17'd18852,17'd18970,17'd37427,17'd37428,17'd37429,17'd37430,17'd37431,17'd30933,17'd29592,17'd27815,17'd10514,17'd27815,17'd27933,17'd29592,17'd32074,17'd30333,17'd25627,17'd30637,17'd25627,17'd5614,17'd5615,17'd5335,17'd25627,17'd37153,17'd37432,17'd37433,17'd37434,17'd9933,17'd31243,17'd28183,17'd37154,17'd37155,17'd37435,17'd37290,17'd37436,17'd37156,17'd37437,17'd37293,17'd37438,17'd37439,17'd37296,17'd37440,17'd37441,17'd37299,17'd37442,17'd37443,17'd37444,17'd37303,17'd19600,17'd2556,17'd36600,17'd6867,17'd447,17'd228,17'd4423,17'd4713,17'd4729,17'd4729,17'd3896,17'd37445,17'd6095,17'd6094,17'd6258,17'd7537,17'd7705,17'd35487,17'd36903,17'd36905,17'd37168,17'd37168,17'd36905,17'd36905,17'd36905,17'd35487,17'd11061,17'd4714,17'd3073,17'd5372,17'd5050,17'd1680,17'd953,17'd771,17'd29891,17'd767,17'd37446,17'd175,17'd37447
},
'{
17'd3903,17'd3902,17'd4243,17'd6420,17'd4246,17'd4246,17'd3101,17'd2934,17'd3592,17'd3901,17'd3592,17'd15496,17'd3428,17'd2422,17'd1689,17'd1127,17'd1416,17'd1416,17'd3905,17'd18,17'd27,17'd286,17'd7385,17'd7385,17'd6745,17'd5972,17'd26731,17'd26469,17'd4581,17'd2948,17'd3261,17'd1706,17'd37448,17'd1708,17'd35620,17'd34168,17'd1561,17'd3266,17'd2953,17'd28077,17'd37449,17'd36607,17'd35065,17'd37450,17'd37451,17'd37452,17'd36462,17'd31917,17'd15008,17'd14767,17'd16987,17'd15902,17'd17207,17'd27461,17'd19006,17'd12361,17'd13093,17'd12357,17'd14468,17'd14469,17'd15516,17'd36757,17'd37453,17'd19263,17'd15014,17'd37454,17'd37455,17'd36191,17'd36191,17'd37181,17'd37456,17'd37457,17'd36333,17'd37458,17'd37459,17'd34367,17'd35074,17'd35920,17'd14230,17'd14109,17'd11631,17'd15151,17'd36764,17'd37186,17'd37057,17'd37320,17'd37320,17'd36919,17'd37460,17'd37056,17'd37323,17'd37323,17'd37186,17'd36471,17'd37461,17'd36337,17'd37462,17'd37463,17'd37464,17'd37465,17'd37466,17'd7602,17'd7603,17'd37467,17'd37468,17'd37334,17'd8731,17'd9046,17'd8886,17'd10338,17'd8569,17'd8725,17'd8410,17'd25677,17'd17472,17'd17607,17'd8247,17'd18808,17'd10607,17'd8877,17'd9189,17'd10335,17'd10334,17'd17847,17'd21985,17'd24538,17'd30526,17'd32761,17'd31287,17'd33875,17'd34037,17'd31288,17'd34704,17'd36211,17'd35372,17'd26872,17'd30229,17'd14264,17'd28352,17'd37469,17'd9340,17'd9743,17'd10175,17'd9194,17'd9348,17'd8410,17'd9744,17'd25147,17'd23343,17'd12426,17'd8419,17'd19780,17'd8578,17'd21987,17'd11404,17'd8410,17'd9194,17'd16552,17'd17728,17'd37470,17'd37471,17'd37472,17'd37473,17'd37474,17'd32591,17'd31588,17'd34203,17'd33730,17'd32933,17'd29786,17'd34390,17'd29336,17'd36783,17'd37206,17'd17726,17'd31774,17'd31602,17'd33102,17'd37342,17'd33411,17'd30841,17'd33886,17'd35105,17'd30240,17'd10844,17'd35808,17'd37209,17'd37475,17'd37476,17'd37477,17'd33596,17'd36496,17'd37478,17'd37479,17'd37480,17'd37481,17'd37482,17'd37483,17'd37484,17'd37485,17'd37486,17'd37487,17'd37488,17'd37489,17'd37490,17'd37491,17'd37492,17'd37493,17'd37096,17'd37494,17'd37096,17'd37096,17'd37095,17'd37231,17'd37363,17'd37230,17'd37363,17'd37363,17'd37365,17'd37365,17'd37365,17'd37365,17'd37365,17'd37365,17'd37363,17'd37363,17'd37363,17'd37231,17'd37231,17'd37095,17'd37495,17'd37366,17'd36964,17'd36820,17'd37226,17'd36383,17'd36105,17'd36243,17'd36383,17'd35970,17'd36387,17'd36821,17'd37496,17'd35964,17'd35135,17'd35135,17'd37235,17'd35273,17'd36522,17'd37371,17'd37497,17'd37498,17'd37499,17'd37500,17'd36830,17'd37501,17'd37502,17'd36682,17'd37379,17'd37503,17'd37504,17'd37505,17'd37505,17'd37382,17'd37506,17'd37507,17'd37383,17'd36398,17'd37508,17'd37509,17'd37384,17'd37384,17'd35567,17'd34104,17'd31035,17'd31035,17'd27372,17'd26174,17'd28597,17'd25320,17'd28851,17'd34137,17'd32008,17'd22678,17'd32344,17'd37510,17'd31657,17'd22324,17'd22678,17'd22328,17'd36543,17'd37511,17'd23215,17'd37117,17'd29529,17'd24415,17'd25177,17'd26064,17'd28725,17'd28486,17'd31352,17'd27642,17'd33319,17'd33654,17'd32507,17'd29249,17'd29536,17'd28857,17'd29536,17'd28857,17'd28857,17'd29831,17'd29831,17'd28728,17'd27885,17'd33163,17'd33642,17'd25568,17'd33666,17'd30446,17'd24089,17'd24088,17'd37512,17'd37389,17'd30126,17'd29100,17'd29378,17'd24902,17'd34467,17'd30126,17'd25178,17'd27882,17'd28597,17'd28598,17'd31055,17'd25833,17'd25429,17'd37513,17'd37514,17'd37515,17'd36999,17'd37516,17'd29984,17'd37517,17'd37518,17'd37519,17'd37520,17'd34130,17'd33169,17'd37521,17'd26188,17'd37522,17'd37523,17'd37524,17'd37525,17'd37526,17'd37527,17'd28613,17'd37528,17'd37264,17'd33818,17'd37529,17'd24910,17'd28610,17'd27887,17'd37530,17'd37531,17'd37532,17'd37533,17'd37534,17'd35591,17'd37535,17'd37536,17'd37537,17'd37538,17'd37539,17'd37540,17'd37541,17'd37542,17'd37543,17'd37544,17'd37545,17'd37546,17'd37547,17'd37548,17'd4984,17'd37549,17'd37550,17'd37551,17'd37552,17'd37553,17'd37554,17'd18135,17'd18852,17'd18970,17'd37555,17'd37556,17'd37557,17'd37558,17'd37559,17'd31551,17'd29592,17'd27815,17'd10515,17'd29592,17'd27933,17'd29592,17'd27696,17'd30638,17'd5160,17'd5004,17'd30333,17'd6390,17'd6219,17'd28185,17'd25627,17'd29024,17'd29295,17'd29295,17'd5166,17'd27696,17'd29592,17'd10642,17'd10514,17'd5763,17'd5012,17'd37435,17'd37436,17'd37560,17'd37561,17'd37562,17'd37563,17'd37564,17'd37565,17'd37566,17'd37567,17'd37568,17'd37569,17'd37570,17'd37444,17'd37571,17'd37572,17'd37573,17'd36600,17'd6867,17'd448,17'd625,17'd4085,17'd4729,17'd3425,17'd3425,17'd3896,17'd37445,17'd6095,17'd6094,17'd6258,17'd7537,17'd7705,17'd35487,17'd36903,17'd37168,17'd37168,17'd37168,17'd36905,17'd36905,17'd36905,17'd35487,17'd11061,17'd4714,17'd5940,17'd5372,17'd4881,17'd445,17'd626,17'd1961,17'd224,17'd37574,17'd31730,17'd37575,17'd37170
},
'{
17'd3903,17'd4892,17'd27951,17'd6420,17'd4246,17'd4246,17'd3101,17'd3101,17'd3428,17'd3901,17'd3592,17'd15358,17'd34512,17'd2422,17'd1689,17'd1127,17'd1416,17'd1416,17'd3905,17'd18,17'd27,17'd286,17'd7061,17'd7061,17'd6745,17'd5972,17'd26731,17'd5211,17'd4581,17'd2948,17'd37576,17'd1705,17'd37448,17'd1708,17'd35620,17'd3439,17'd3436,17'd3109,17'd2796,17'd37577,17'd3767,17'd4592,17'd26479,17'd35773,17'd37578,17'd37579,17'd37580,17'd31918,17'd14893,17'd14768,17'd16033,17'd17445,17'd18656,17'd19753,17'd11764,17'd12218,17'd12527,17'd14469,17'd14468,17'd12357,17'd35352,17'd37581,17'd37582,17'd18418,17'd36759,17'd37583,17'd37583,17'd34363,17'd34363,17'd37584,17'd37585,17'd37586,17'd37587,17'd37588,17'd37589,17'd33228,17'd15655,17'd14782,17'd13104,17'd14109,17'd13611,17'd37590,17'd37591,17'd36471,17'd37592,17'd37593,17'd37320,17'd37057,17'd37321,17'd37594,17'd7103,17'd37323,17'd37056,17'd37595,17'd37461,17'd36618,17'd37596,17'd37597,17'd37598,17'd37599,17'd37600,17'd37601,17'd37602,17'd37603,17'd37468,17'd23342,17'd8573,17'd37604,17'd8729,17'd10177,17'd8731,17'd8572,17'd8409,17'd23861,17'd37605,17'd17607,17'd9744,17'd9349,17'd22473,17'd16067,17'd9189,17'd10026,17'd17965,17'd29335,17'd23513,17'd26371,17'd37606,17'd32761,17'd31287,17'd33720,17'd31288,17'd31288,17'd31773,17'd36211,17'd28460,17'd27123,17'd24362,17'd18327,17'd27623,17'd18916,17'd10744,17'd9347,17'd9038,17'd16067,17'd8724,17'd9482,17'd9744,17'd8413,17'd8578,17'd12426,17'd8419,17'd8733,17'd8578,17'd8413,17'd14675,17'd10027,17'd10175,17'd16911,17'd17232,17'd37607,17'd37608,17'd37609,17'd37610,17'd26628,17'd30971,17'd31941,17'd33875,17'd33096,17'd30678,17'd29644,17'd28349,17'd28349,17'd37611,17'd28232,17'd16560,17'd29934,17'd32939,17'd36356,17'd32940,17'd30089,17'd34049,17'd36078,17'd37612,17'd30240,17'd11271,17'd29348,17'd37613,17'd29948,17'd37614,17'd37615,17'd37616,17'd37617,17'd37618,17'd37619,17'd37620,17'd37621,17'd37622,17'd35821,17'd37623,17'd37624,17'd37625,17'd37626,17'd37627,17'd37628,17'd37629,17'd37630,17'd37631,17'd37632,17'd37633,17'd37230,17'd37634,17'd37366,17'd37367,17'd37634,17'd37367,17'd37096,17'd37368,17'd37368,17'd37366,17'd37495,17'd37635,17'd37635,17'd37636,17'd37636,17'd37230,17'd37095,17'd37095,17'd37230,17'd37363,17'd37363,17'd37230,17'd37096,17'd36963,17'd37097,17'd36964,17'd36820,17'd36243,17'd36383,17'd36383,17'd35839,17'd35271,17'd36521,17'd36108,17'd36821,17'd35135,17'd36672,17'd35407,17'd36247,17'd37637,17'd37638,17'd37639,17'd37640,17'd37641,17'd37642,17'd37643,17'd37644,17'd37645,17'd37646,17'd37647,17'd37648,17'd37649,17'd37650,17'd37651,17'd37652,17'd37244,17'd37507,17'd37653,17'd37654,17'd37655,17'd37656,17'd37384,17'd37384,17'd37657,17'd37658,17'd30735,17'd28486,17'd30586,17'd25833,17'd25567,17'd29103,17'd28977,17'd30275,17'd23388,17'd22680,17'd22506,17'd22158,17'd37659,17'd22324,17'd22680,17'd22328,17'd33158,17'd31828,17'd33158,17'd23217,17'd29830,17'd24090,17'd25568,17'd28720,17'd28724,17'd30586,17'd32016,17'd27642,17'd33319,17'd33654,17'd32507,17'd29249,17'd29536,17'd30884,17'd29536,17'd28857,17'd28857,17'd29831,17'd29536,17'd28372,17'd26276,17'd25560,17'd28366,17'd28254,17'd24417,17'd24742,17'd35722,17'd35722,17'd30126,17'd29533,17'd32007,17'd24252,17'd29102,17'd28852,17'd34467,17'd24895,17'd25178,17'd27882,17'd28597,17'd28598,17'd31055,17'd26174,17'd25429,17'd26780,17'd27885,17'd37515,17'd36999,17'd37257,17'd37660,17'd37661,17'd37662,17'd37663,17'd37520,17'd37664,17'd30285,17'd29836,17'd24430,17'd37665,17'd35588,17'd37666,17'd37526,17'd36711,17'd37667,17'd37668,17'd37669,17'd37670,17'd33338,17'd29705,17'd37671,17'd37672,17'd32366,17'd32849,17'd30292,17'd29994,17'd37673,17'd33479,17'd37674,17'd37675,17'd37676,17'd37015,17'd37677,17'd37678,17'd37679,17'd37680,17'd37681,17'd37682,17'd35746,17'd37683,17'd37684,17'd37685,17'd37686,17'd37687,17'd37688,17'd37689,17'd37551,17'd37690,17'd37691,17'd37692,17'd18261,17'd19480,17'd18970,17'd37555,17'd37693,17'd37694,17'd37695,17'd37696,17'd31551,17'd29592,17'd27815,17'd10515,17'd29592,17'd27933,17'd27933,17'd9933,17'd31717,17'd28185,17'd25627,17'd25627,17'd27935,17'd5614,17'd5335,17'd25627,17'd4848,17'd28778,17'd29594,17'd5329,17'd7668,17'd29593,17'd10642,17'd37154,17'd5616,17'd37697,17'd37698,17'd36587,17'd37699,17'd37700,17'd37293,17'd37701,17'd37702,17'd37565,17'd37703,17'd37704,17'd37705,17'd37569,17'd24661,17'd37706,17'd37571,17'd37572,17'd37707,17'd36454,17'd8788,17'd448,17'd446,17'd3897,17'd3423,17'd3246,17'd3423,17'd37708,17'd37709,17'd4867,17'd6094,17'd6094,17'd7537,17'd7705,17'd35487,17'd36903,17'd35487,17'd35487,17'd37168,17'd37168,17'd36905,17'd36903,17'd12923,17'd2906,17'd6889,17'd5940,17'd5372,17'd3743,17'd2417,17'd953,17'd771,17'd29891,17'd37574,17'd31904,17'd33377,17'd36604
},
'{
17'd9960,17'd4244,17'd4243,17'd6420,17'd4246,17'd14743,17'd3101,17'd3427,17'd3592,17'd3901,17'd3592,17'd15358,17'd34512,17'd2422,17'd1689,17'd1127,17'd1416,17'd1416,17'd3905,17'd18,17'd27,17'd286,17'd7061,17'd7061,17'd6745,17'd5972,17'd12931,17'd5211,17'd4896,17'd2948,17'd37171,17'd1705,17'd1426,17'd1427,17'd3439,17'd3437,17'd3266,17'd3109,17'd2796,17'd37710,17'd3610,17'd4753,17'd4447,17'd37711,17'd37712,17'd37713,17'd36610,17'd31918,17'd14893,17'd14768,17'd16033,17'd17320,17'd18656,17'd19753,17'd11764,17'd12814,17'd12527,17'd16284,17'd14468,17'd11762,17'd11359,17'd34939,17'd19016,17'd18302,17'd37714,17'd37715,17'd37716,17'd34363,17'd37717,17'd37718,17'd37719,17'd37720,17'd37587,17'd37588,17'd37721,17'd33864,17'd17330,17'd17105,17'd9707,17'd9164,17'd16042,17'd27835,17'd37323,17'd36471,17'd37320,17'd37722,17'd37320,17'd37058,17'd37460,17'd37723,17'd37322,17'd37322,17'd37056,17'd37724,17'd37461,17'd36618,17'd37725,17'd7113,17'd37726,17'd37727,17'd37728,17'd37729,17'd37730,17'd37731,17'd37732,17'd8577,17'd17481,17'd8730,17'd8729,17'd30217,17'd8571,17'd15429,17'd8409,17'd23861,17'd37605,17'd16440,17'd10177,17'd11404,17'd9046,17'd24999,17'd9189,17'd10026,17'd17965,17'd34956,17'd24858,17'd28105,17'd37733,17'd32761,17'd31287,17'd33720,17'd31288,17'd33727,17'd36937,17'd29645,17'd28227,17'd30076,17'd24363,17'd12583,17'd22820,17'd20607,17'd23679,17'd9743,17'd10336,17'd9194,17'd8879,17'd30969,17'd9744,17'd8573,17'd8578,17'd18202,17'd8419,17'd37734,17'd8578,17'd8413,17'd9482,17'd10027,17'd10336,17'd37336,17'd37607,17'd27744,17'd37735,17'd34956,17'd37736,17'd34962,17'd37737,17'd36490,17'd33243,17'd31591,17'd30079,17'd37611,17'd37738,17'd37738,17'd37739,17'd28233,17'd13642,17'd32294,17'd32773,17'd37740,17'd32940,17'd33245,17'd37741,17'd36078,17'd34969,17'd37742,17'd37743,17'd37744,17'd37475,17'd37745,17'd37746,17'd37747,17'd36642,17'd37617,17'd37748,17'd37749,17'd36500,17'd37750,17'd37751,17'd37752,17'd37753,17'd37754,17'd37755,17'd37756,17'd37757,17'd37758,17'd37759,17'd37760,17'd36238,17'd37761,17'd37762,17'd37361,17'd37363,17'd37362,17'd37231,17'd37363,17'd37096,17'd37096,17'd37095,17'd37095,17'd37095,17'd37096,17'd37636,17'd37635,17'd37635,17'd37635,17'd37096,17'd37096,17'd37095,17'd37096,17'd37096,17'd37096,17'd37230,17'd37231,17'd37763,17'd36818,17'd37097,17'd36964,17'd36243,17'd35683,17'd35683,17'd35683,17'd35550,17'd35550,17'd36821,17'd36107,17'd35272,17'd36387,17'd33620,17'd36247,17'd35273,17'd37764,17'd37765,17'd37766,17'd37767,17'd37768,17'd37769,17'd37770,17'd37771,17'd37772,17'd37773,17'd37379,17'd37648,17'd37650,17'd37774,17'd37652,17'd37244,17'd37775,17'd37776,17'd36981,17'd37655,17'd37656,17'd37384,17'd37384,17'd37657,17'd37777,17'd32016,17'd28486,17'd30586,17'd26903,17'd28594,17'd28850,17'd25031,17'd28722,17'd23387,17'd22679,17'd22677,17'd30426,17'd35429,17'd22325,17'd32827,17'd22501,17'd32008,17'd31828,17'd36543,17'd23217,17'd29830,17'd30879,17'd25178,17'd26064,17'd28725,17'd28486,17'd31352,17'd27642,17'd33319,17'd33654,17'd32017,17'd32018,17'd29536,17'd30884,17'd29536,17'd28857,17'd28857,17'd29831,17'd28857,17'd29380,17'd26278,17'd28365,17'd37778,17'd28254,17'd28718,17'd24742,17'd35722,17'd35722,17'd28851,17'd29533,17'd25031,17'd24417,17'd23562,17'd28975,17'd24252,17'd25032,17'd25178,17'd27882,17'd33000,17'd28599,17'd32669,17'd25949,17'd25945,17'd25555,17'd30279,17'd37779,17'd36849,17'd36999,17'd35580,17'd35443,17'd36266,17'd34469,17'd37780,17'd37127,17'd30454,17'd37781,17'd28731,17'd28605,17'd27888,17'd29117,17'd37782,17'd36711,17'd36711,17'd37783,17'd37670,17'd37784,17'd37785,17'd37786,17'd37529,17'd24910,17'd37672,17'd37787,17'd36549,17'd36994,17'd23738,17'd34638,17'd32501,17'd37788,17'd37789,17'd37790,17'd29722,17'd37413,17'd37791,17'd34782,17'd37792,17'd37793,17'd37794,17'd37795,17'd37796,17'd37797,17'd8908,17'd37798,17'd37799,17'd37689,17'd37800,17'd37690,17'd37691,17'd37801,17'd20115,17'd19480,17'd18970,17'd37555,17'd37802,17'd37803,17'd37804,17'd37805,17'd32875,17'd31243,17'd29592,17'd10515,17'd27933,17'd27933,17'd27933,17'd9933,17'd31717,17'd28185,17'd25627,17'd30333,17'd6554,17'd6390,17'd28185,17'd5160,17'd4848,17'd28778,17'd30486,17'd5002,17'd7499,17'd9933,17'd10642,17'd10514,17'd5337,17'd5010,17'd37806,17'd36587,17'd37807,17'd37808,17'd37809,17'd37810,17'd37811,17'd37812,17'd37813,17'd37814,17'd37815,17'd37038,17'd37816,17'd37817,17'd37818,17'd37819,17'd37820,17'd36454,17'd8788,17'd8314,17'd1824,17'd3897,17'd3423,17'd5939,17'd37821,17'd37708,17'd37709,17'd4867,17'd16623,17'd6094,17'd7537,17'd7705,17'd35487,17'd35487,17'd35487,17'd35487,17'd37168,17'd37168,17'd36905,17'd36905,17'd35487,17'd11061,17'd4714,17'd5940,17'd5371,17'd4881,17'd1401,17'd623,17'd799,17'd22264,17'd767,17'd31730,17'd33377,17'd36604
},
'{
17'd4244,17'd4243,17'd25384,17'd6420,17'd4246,17'd4246,17'd2934,17'd3427,17'd3901,17'd3901,17'd3901,17'd3428,17'd3251,17'd1831,17'd1127,17'd466,17'd4089,17'd4089,17'd653,17'd652,17'd286,17'd286,17'd7061,17'd6745,17'd5973,17'd26730,17'd12931,17'd5055,17'd4252,17'd3260,17'd2608,17'd37822,17'd1426,17'd1561,17'd3439,17'd24674,17'd24674,17'd32255,17'd23660,17'd15749,17'd37823,17'd20282,17'd37050,17'd37824,17'd37825,17'd37826,17'd34936,17'd37827,17'd14893,17'd16768,17'd17810,17'd17319,17'd18174,17'd18412,17'd11627,17'd12679,17'd12062,17'd14763,17'd22802,17'd11625,17'd37828,17'd19389,17'd37829,17'd14899,17'd37830,17'd37831,17'd37832,17'd37717,17'd37833,17'd36466,17'd37317,17'd37586,17'd36762,17'd37834,17'd37835,17'd33070,17'd15655,17'd14782,17'd9164,17'd29182,17'd16042,17'd13612,17'd37323,17'd37836,17'd37837,17'd37838,17'd37839,17'd37058,17'd37460,17'd37723,17'd37840,17'd37594,17'd36194,17'd37724,17'd37841,17'd37842,17'd37060,17'd37843,17'd37844,17'd37845,17'd37846,17'd37847,17'd37848,17'd37849,17'd7783,17'd9196,17'd17481,17'd8571,17'd24368,17'd30217,17'd35514,17'd8413,17'd8409,17'd26038,17'd37850,17'd9042,17'd34699,17'd12425,17'd23861,17'd16067,17'd9189,17'd9340,17'd10170,17'd34956,17'd26258,17'd26872,17'd30832,17'd37851,17'd32283,17'd33720,17'd31288,17'd34835,17'd31587,17'd31768,17'd27984,17'd25925,17'd19920,17'd11130,17'd37852,17'd16683,17'd10744,17'd9347,17'd9038,17'd9040,17'd8725,17'd30969,17'd11404,17'd8574,17'd8578,17'd18919,17'd8248,17'd9196,17'd15945,17'd8573,17'd8726,17'd9045,17'd15944,17'd17232,17'd17717,17'd27744,17'd27351,17'd37853,17'd37854,17'd31594,17'd30972,17'd34203,17'd33095,17'd31597,17'd37855,17'd28349,17'd37856,17'd17725,17'd37857,17'd17724,17'd31953,17'd33417,17'd37858,17'd31956,17'd33251,17'd36078,17'd37859,17'd37860,17'd37861,17'd10844,17'd37862,17'd37863,17'd36789,17'd37864,17'd37865,17'd37747,17'd37866,17'd36497,17'd37867,17'd37868,17'd37869,17'd33901,17'd37870,17'd37871,17'd37872,17'd37873,17'd37874,17'd37875,17'd37876,17'd37877,17'd37878,17'd37879,17'd36965,17'd37880,17'd37362,17'd37881,17'd37882,17'd37763,17'd37881,17'd37881,17'd37882,17'd37881,17'd37494,17'd37363,17'd37362,17'd37494,17'd37363,17'd37231,17'd37231,17'd37095,17'd37095,17'd37095,17'd37230,17'd37095,17'd37096,17'd37495,17'd37495,17'd37495,17'd37230,17'd37231,17'd37883,17'd36668,17'd36820,17'd36243,17'd36383,17'd36105,17'd37884,17'd37885,17'd36106,17'd35838,17'd36387,17'd36521,17'd36965,17'd35407,17'd36965,17'd37886,17'd37887,17'd37888,17'd37889,17'd37890,17'd37891,17'd37892,17'd37893,17'd37894,17'd37895,17'd37647,17'd37896,17'd37896,17'd37897,17'd37898,17'd37899,17'd37900,17'd37901,17'd37902,17'd37903,17'd37904,17'd37905,17'd37905,17'd37906,17'd37907,17'd37908,17'd26901,17'd35011,17'd26903,17'd28723,17'd29101,17'd25179,17'd30879,17'd23387,17'd23389,17'd23573,17'd22506,17'd31343,17'd33311,17'd22503,17'd23218,17'd23569,17'd31828,17'd33158,17'd29973,17'd29686,17'd30879,17'd25178,17'd25566,17'd28724,17'd33163,17'd32016,17'd29379,17'd27885,17'd32354,17'd33165,17'd28982,17'd34114,17'd33166,17'd29106,17'd28857,17'd29537,17'd29831,17'd36132,17'd29380,17'd26780,17'd25702,17'd37909,17'd23914,17'd23561,17'd24415,17'd23731,17'd24090,17'd24742,17'd25031,17'd33483,17'd24745,17'd24252,17'd23562,17'd28601,17'd25032,17'd29103,17'd27882,17'd25567,17'd28598,17'd31055,17'd26062,17'd25312,17'd25555,17'd27885,17'd37779,17'd37515,17'd36849,17'd37910,17'd37660,17'd29835,17'd34469,17'd37780,17'd37520,17'd37911,17'd28860,17'd28731,17'd37912,17'd26905,17'd37913,17'd27375,17'd27031,17'd37914,17'd37915,17'd37916,17'd37917,17'd37917,17'd37918,17'd37919,17'd27033,17'd25042,17'd37920,17'd37921,17'd36268,17'd37922,17'd34278,17'd31498,17'd37923,17'd37924,17'd37925,17'd37926,17'd37927,17'd37928,17'd37929,17'd37930,17'd37931,17'd37932,17'd37933,17'd21282,17'd37934,17'd33360,17'd37935,17'd14022,17'd37936,17'd37937,17'd37552,17'd37938,17'd37939,17'd20115,17'd19847,17'd16955,17'd37940,17'd37802,17'd37941,17'd37942,17'd37943,17'd29158,17'd27933,17'd9933,17'd9933,17'd27933,17'd28183,17'd27933,17'd27815,17'd6219,17'd27935,17'd31553,17'd31553,17'd31717,17'd5614,17'd5336,17'd5330,17'd34921,17'd34791,17'd29595,17'd4841,17'd6219,17'd27696,17'd27815,17'd37154,17'd5764,17'd37944,17'd37945,17'd37946,17'd37947,17'd37808,17'd37948,17'd37810,17'd37811,17'd37812,17'd37949,17'd37950,17'd37815,17'd37951,17'd37952,17'd37953,17'd2541,17'd37819,17'd37954,17'd37955,17'd37956,17'd6867,17'd795,17'd5357,17'd4712,17'd6085,17'd5938,17'd37957,17'd37958,17'd4867,17'd37959,17'd6258,17'd7537,17'd7537,17'd33051,17'd36903,17'd35487,17'd33051,17'd33051,17'd35487,17'd36905,17'd35487,17'd12923,17'd2906,17'd6889,17'd5630,17'd4880,17'd3743,17'd1262,17'd954,17'd3100,17'd22264,17'd767,17'd31564,17'd33377,17'd37960
},
'{
17'd4244,17'd4244,17'd4892,17'd6420,17'd4246,17'd4246,17'd2934,17'd3427,17'd3901,17'd3901,17'd3901,17'd3428,17'd3251,17'd1831,17'd1127,17'd2,17'd4089,17'd4089,17'd653,17'd652,17'd286,17'd1833,17'd7061,17'd7060,17'd6438,17'd26468,17'd12507,17'd5055,17'd4252,17'd3107,17'd2268,17'd1139,17'd1141,17'd1561,17'd3437,17'd24674,17'd32731,17'd2952,17'd23660,17'd37961,17'd4105,17'd4593,17'd4110,17'd37962,17'd37963,17'd37964,17'd34936,17'd33549,17'd14768,17'd16411,17'd17445,17'd19255,17'd18774,17'd20423,17'd12530,17'd12679,17'd14469,17'd16284,17'd15763,17'd11359,17'd37965,17'd37966,17'd18302,17'd16174,17'd37967,17'd37831,17'd37968,17'd37833,17'd37833,17'd36466,17'd37317,17'd36333,17'd37969,17'd37834,17'd35358,17'd35217,17'd35920,17'd14230,17'd14109,17'd9015,17'd8852,17'd27962,17'd37322,17'd37970,17'd37971,17'd37838,17'd37839,17'd37972,17'd37973,17'd37974,17'd37975,17'd37974,17'd36472,17'd36919,17'd37976,17'd37977,17'd37188,17'd37978,17'd37979,17'd37980,17'd37981,17'd37982,17'd7281,17'd37849,17'd14005,17'd25148,17'd25147,17'd8731,17'd24368,17'd8247,17'd25147,17'd21987,17'd8409,17'd16067,17'd22814,17'd22645,17'd31438,17'd12425,17'd23861,17'd16067,17'd9189,17'd9340,17'd10170,17'd35230,17'd26150,17'd28343,17'd30832,17'd37851,17'd31287,17'd33875,17'd31288,17'd34835,17'd31587,17'd28461,17'd26873,17'd24208,17'd23167,17'd13521,17'd10167,17'd10992,17'd9340,17'd9346,17'd8874,17'd9041,17'd8879,17'd9482,17'd11966,17'd8731,17'd25147,17'd12867,17'd21208,17'd21987,17'd8573,17'd10607,17'd8881,17'd9041,17'd15807,17'd17232,17'd17717,17'd10332,17'd34826,17'd37983,17'd33572,17'd37984,17'd30972,17'd33568,17'd31591,17'd37985,17'd37986,17'd37738,17'd37738,17'd17725,17'd17724,17'd17013,17'd31138,17'd32295,17'd31141,17'd31956,17'd35935,17'd37987,17'd37988,17'd37860,17'd37861,17'd29810,17'd37744,17'd37613,17'd37989,17'd37990,17'd37865,17'd37991,17'd37992,17'd37992,17'd37993,17'd37994,17'd37995,17'd37996,17'd37997,17'd37998,17'd37999,17'd38000,17'd38001,17'd37357,17'd38002,17'd38003,17'd38004,17'd38005,17'd38006,17'd37231,17'd36660,17'd36660,17'd36964,17'd36660,17'd36963,17'd36818,17'd36963,17'd36963,17'd37096,17'd37495,17'd37095,17'd37231,17'd37230,17'd37231,17'd37363,17'd37230,17'd37231,17'd37231,17'd37230,17'd37095,17'd37096,17'd37495,17'd37366,17'd37366,17'd37366,17'd37095,17'd38007,17'd37883,17'd36668,17'd37226,17'd36383,17'd36383,17'd38008,17'd37884,17'd35970,17'd36106,17'd36387,17'd35682,17'd38009,17'd37234,17'd36965,17'd38010,17'd37887,17'd38011,17'd38012,17'd38013,17'd38014,17'd36257,17'd38015,17'd38016,17'd38017,17'd37773,17'd38018,17'd38019,17'd37897,17'd37652,17'd38020,17'd38021,17'd38022,17'd38023,17'd38024,17'd37904,17'd37905,17'd37905,17'd37906,17'd37907,17'd38025,17'd28979,17'd32016,17'd28725,17'd28602,17'd25317,17'd29244,17'd24090,17'd29827,17'd23216,17'd22859,17'd22506,17'd22858,17'd22331,17'd33158,17'd23215,17'd23569,17'd31828,17'd33158,17'd29973,17'd29686,17'd23731,17'd25178,17'd27766,17'd28725,17'd31035,17'd31352,17'd29379,17'd30279,17'd28134,17'd33320,17'd38026,17'd34114,17'd32833,17'd29106,17'd28857,17'd29537,17'd29536,17'd29979,17'd29380,17'd26780,17'd25831,17'd38027,17'd24412,17'd28601,17'd24415,17'd30879,17'd30879,17'd24742,17'd25031,17'd33483,17'd24897,17'd24417,17'd28008,17'd28601,17'd25032,17'd29103,17'd27882,17'd25567,17'd28598,17'd31055,17'd26062,17'd25312,17'd25555,17'd27885,17'd28134,17'd37779,17'd37515,17'd36858,17'd37910,17'd38028,17'd29695,17'd37780,17'd38029,17'd38030,17'd30147,17'd33657,17'd38031,17'd38032,17'd36552,17'd38033,17'd38034,17'd38035,17'd38036,17'd34119,17'd38037,17'd29252,17'd28497,17'd28985,17'd28501,17'd25584,17'd37920,17'd38038,17'd38039,17'd32852,17'd38040,17'd38041,17'd38042,17'd38043,17'd38044,17'd38045,17'd38046,17'd38047,17'd38048,17'd35597,17'd38049,17'd38050,17'd35885,17'd38051,17'd37934,17'd9212,17'd5907,17'd38052,17'd37936,17'd38053,17'd38054,17'd38055,17'd37939,17'd21310,17'd19847,17'd16955,17'd37940,17'd38056,17'd37693,17'd37694,17'd38057,17'd34502,17'd27933,17'd9933,17'd9933,17'd27933,17'd28183,17'd27933,17'd27815,17'd6219,17'd27935,17'd30333,17'd31553,17'd31717,17'd6390,17'd27935,17'd5160,17'd5162,17'd5155,17'd38058,17'd5328,17'd5615,17'd7668,17'd27815,17'd10514,17'd5763,17'd38059,17'd38060,17'd37946,17'd37947,17'd37808,17'd37562,17'd38061,17'd38062,17'd38063,17'd38064,17'd38065,17'd37704,17'd38066,17'd38067,17'd38068,17'd2374,17'd38069,17'd37954,17'd38070,17'd22263,17'd8788,17'd38071,17'd6085,17'd4558,17'd4558,17'd5938,17'd37957,17'd37958,17'd38072,17'd37959,17'd16492,17'd7364,17'd7537,17'd33051,17'd35487,17'd35487,17'd33051,17'd33051,17'd35487,17'd36905,17'd37168,17'd35487,17'd2906,17'd6889,17'd5630,17'd4880,17'd3743,17'd1262,17'd623,17'd1122,17'd962,17'd786,17'd38073,17'd38074,17'd34668
},
'{
17'd4244,17'd4892,17'd25384,17'd6420,17'd14743,17'd4246,17'd3101,17'd3427,17'd3901,17'd3901,17'd3901,17'd3428,17'd3251,17'd1831,17'd1127,17'd2,17'd4089,17'd4089,17'd653,17'd652,17'd286,17'd1833,17'd7061,17'd6745,17'd5973,17'd5803,17'd13067,17'd4894,17'd2948,17'd3261,17'd1706,17'd1139,17'd1141,17'd1979,17'd3437,17'd24674,17'd32731,17'd38075,17'd13441,17'd38076,17'd3768,17'd38077,17'd37309,17'd15886,17'd38078,17'd38079,17'd38080,17'd15008,17'd16768,17'd16033,17'd17320,17'd17206,17'd18774,17'd12681,17'd12530,17'd12679,17'd14469,17'd16284,17'd11625,17'd38081,17'd38082,17'd14774,17'd38083,17'd38084,17'd38085,17'd38086,17'd38087,17'd38088,17'd37833,17'd38089,17'd33225,17'd37587,17'd38090,17'd38091,17'd33706,17'd15655,17'd14782,17'd13104,17'd14109,17'd9015,17'd24843,17'd24980,17'd37322,17'd38092,17'd37971,17'd38093,17'd6644,17'd38094,17'd38095,17'd38096,17'd38096,17'd37974,17'd37724,17'd38097,17'd38098,17'd38099,17'd38100,17'd38101,17'd38102,17'd38103,17'd38104,17'd38105,17'd38106,17'd38107,17'd14005,17'd8578,17'd17481,17'd8575,17'd8571,17'd12586,17'd25147,17'd25147,17'd8409,17'd8877,17'd25814,17'd22645,17'd10338,17'd8729,17'd12424,17'd8876,17'd21984,17'd9340,17'd10332,17'd13368,17'd23170,17'd28227,17'd30832,17'd30834,17'd34203,17'd33875,17'd31288,17'd34835,17'd29330,17'd28462,17'd27123,17'd24362,17'd21985,17'd14132,17'd15300,17'd17012,17'd9341,17'd9346,17'd8874,17'd8720,17'd8881,17'd20176,17'd8724,17'd8731,17'd25147,17'd14812,17'd9887,17'd24862,17'd8574,17'd10607,17'd8881,17'd9041,17'd14674,17'd17601,17'd17965,17'd10332,17'd29335,17'd22991,17'd24539,17'd28106,17'd30972,17'd34835,17'd36214,17'd30680,17'd38108,17'd37856,17'd28233,17'd17726,17'd18685,17'd16686,17'd35520,17'd38109,17'd38110,17'd30381,17'd35935,17'd29938,17'd38111,17'd38112,17'd34395,17'd36938,17'd29350,17'd37073,17'd36641,17'd38113,17'd37865,17'd37991,17'd38114,17'd37991,17'd35114,17'd38115,17'd38116,17'd38117,17'd38118,17'd38119,17'd38120,17'd38121,17'd38122,17'd38123,17'd38124,17'd38125,17'd38126,17'd36240,17'd38127,17'd38128,17'd37882,17'd38129,17'd36668,17'd36660,17'd37097,17'd36819,17'd36819,17'd36668,17'd36963,17'd36668,17'd36668,17'd36668,17'd36668,17'd36818,17'd38130,17'd38130,17'd37230,17'd37230,17'd37095,17'd37095,17'd37095,17'd37495,17'd37366,17'd37368,17'd37367,17'd37368,17'd37096,17'd37231,17'd37096,17'd36669,17'd36243,17'd38008,17'd38131,17'd38132,17'd35550,17'd35970,17'd36106,17'd35838,17'd38133,17'd38134,17'd36965,17'd38135,17'd38136,17'd38137,17'd38138,17'd38139,17'd38140,17'd38141,17'd38142,17'd37645,17'd38143,17'd38144,17'd38018,17'd38019,17'd38145,17'd38146,17'd38020,17'd38147,17'd38148,17'd38149,17'd37112,17'd38150,17'd38151,17'd38151,17'd38152,17'd38153,17'd35152,17'd31035,17'd35011,17'd28725,17'd28602,17'd28484,17'd29103,17'd24743,17'd29827,17'd23218,17'd22677,17'd22506,17'd22857,17'd22331,17'd36543,17'd32191,17'd29829,17'd31828,17'd33158,17'd29973,17'd23923,17'd23731,17'd25178,17'd25566,17'd28724,17'd33163,17'd32016,17'd29246,17'd30279,17'd32832,17'd38154,17'd38155,17'd34114,17'd32833,17'd29106,17'd29106,17'd28728,17'd28728,17'd29831,17'd30587,17'd29245,17'd28724,17'd38156,17'd28718,17'd28008,17'd24415,17'd30275,17'd28722,17'd24252,17'd32007,17'd33483,17'd25030,17'd24744,17'd28367,17'd29240,17'd24898,17'd29103,17'd27882,17'd25567,17'd28597,17'd33000,17'd26064,17'd26782,17'd28980,17'd27885,17'd28134,17'd38157,17'd38158,17'd38159,17'd38160,17'd38028,17'd36266,17'd37780,17'd38029,17'd38030,17'd33817,17'd37405,17'd38161,17'd32212,17'd38162,17'd32361,17'd26290,17'd36412,17'd38163,17'd38164,17'd28022,17'd38165,17'd29263,17'd38166,17'd29110,17'd32204,17'd38167,17'd38168,17'd38169,17'd38170,17'd38171,17'd38172,17'd38173,17'd38174,17'd38175,17'd38176,17'd36013,17'd38177,17'd38178,17'd38179,17'd38180,17'd38181,17'd38182,17'd38183,17'd38184,17'd38185,17'd5752,17'd38186,17'd38187,17'd38188,17'd38189,17'd38055,17'd37938,17'd37939,17'd19847,17'd16955,17'd37940,17'd38056,17'd37802,17'd38190,17'd38191,17'd28057,17'd27933,17'd9933,17'd9933,17'd27933,17'd27933,17'd27933,17'd9933,17'd6219,17'd28185,17'd30333,17'd31553,17'd31891,17'd5614,17'd5762,17'd5334,17'd34921,17'd5155,17'd38058,17'd4995,17'd5762,17'd7668,17'd9933,17'd8934,17'd5616,17'd38060,17'd38192,17'd38193,17'd38194,17'd38195,17'd37562,17'd38196,17'd37811,17'd3539,17'd38197,17'd3361,17'd37704,17'd38198,17'd3047,17'd38199,17'd2726,17'd3066,17'd19600,17'd21016,17'd38200,17'd8788,17'd4059,17'd4558,17'd5937,17'd5356,17'd38201,17'd38202,17'd37958,17'd38203,17'd37959,17'd6258,17'd7537,17'd7537,17'd33051,17'd35487,17'd35487,17'd33051,17'd33051,17'd35487,17'd36905,17'd35487,17'd12923,17'd2906,17'd3073,17'd6415,17'd445,17'd1401,17'd1262,17'd954,17'd609,17'd962,17'd18515,17'd618,17'd33540,17'd34345
},
'{
17'd4244,17'd4244,17'd4892,17'd6420,17'd14743,17'd4246,17'd3101,17'd3427,17'd3901,17'd3901,17'd3901,17'd3428,17'd3101,17'd1831,17'd1127,17'd2,17'd4089,17'd4089,17'd653,17'd652,17'd286,17'd1833,17'd7061,17'd6437,17'd5803,17'd5804,17'd13067,17'd4894,17'd2948,17'd2608,17'd1706,17'd18150,17'd2949,17'd1979,17'd3437,17'd32731,17'd32090,17'd38204,17'd29899,17'd38205,17'd26132,17'd4594,17'd38206,17'd38207,17'd38208,17'd38209,17'd31917,17'd32739,17'd16411,17'd16169,17'd17207,17'd17206,17'd17689,17'd12681,17'd12218,17'd13093,17'd12678,17'd12527,17'd38210,17'd34939,17'd38211,17'd38212,17'd38213,17'd37830,17'd37831,17'd38086,17'd38087,17'd38214,17'd37717,17'd37456,17'd38215,17'd38216,17'd38217,17'd37589,17'd33228,17'd17330,17'd17105,17'd14109,17'd9164,17'd8699,17'd38218,17'd24979,17'd38219,17'd38220,17'd6643,17'd38093,17'd38221,17'd6644,17'd38222,17'd38223,17'd38223,17'd37973,17'd38097,17'd38224,17'd38225,17'd38226,17'd38227,17'd38228,17'd38229,17'd38230,17'd38231,17'd38232,17'd38233,17'd38234,17'd14136,17'd23343,17'd25147,17'd8575,17'd8571,17'd10339,17'd23343,17'd8578,17'd19535,17'd8877,17'd14674,17'd22645,17'd24367,17'd16205,17'd23517,17'd8723,17'd9043,17'd9340,17'd33725,17'd35799,17'd24031,17'd28344,17'd37065,17'd33718,17'd31287,17'd33875,17'd34203,17'd34381,17'd29330,17'd29328,17'd28105,17'd21505,17'd22817,17'd38235,17'd21503,17'd10992,17'd9620,17'd9344,17'd10174,17'd9043,17'd8883,17'd15297,17'd9195,17'd8724,17'd9744,17'd24213,17'd25147,17'd8572,17'd8728,17'd8725,17'd8881,17'd10175,17'd14674,17'd37607,17'd38236,17'd13522,17'd11526,17'd37196,17'd26496,17'd28106,17'd30972,17'd32933,17'd32444,17'd38237,17'd38108,17'd37856,17'd28233,17'd28232,17'd38238,17'd38239,17'd33249,17'd32609,17'd32940,17'd33251,17'd37987,17'd29938,17'd10598,17'd34711,17'd38240,17'd38241,17'd29950,17'd38242,17'd33744,17'd33264,17'd37747,17'd37867,17'd38243,17'd38244,17'd38245,17'd38246,17'd38247,17'd38248,17'd38249,17'd38250,17'd38251,17'd38252,17'd38253,17'd38254,17'd38255,17'd38256,17'd38257,17'd38258,17'd38259,17'd38260,17'd37763,17'd38129,17'd36817,17'd36668,17'd36819,17'd37097,17'd37097,17'd36819,17'd37097,17'd37097,17'd36819,17'd36819,17'd36819,17'd36819,17'd36819,17'd36819,17'd37366,17'd37366,17'd37495,17'd37095,17'd37095,17'd37096,17'd37366,17'd37367,17'd37368,17'd37634,17'd37634,17'd37366,17'd37495,17'd37368,17'd36964,17'd36243,17'd38261,17'd36671,17'd35683,17'd35683,17'd35839,17'd35970,17'd38262,17'd38263,17'd36246,17'd38264,17'd38265,17'd38266,17'd38267,17'd38268,17'd38269,17'd38270,17'd38142,17'd37771,17'd37894,17'd38017,17'd38271,17'd38272,17'd38273,17'd38274,17'd38020,17'd38275,17'd38276,17'd38277,17'd37654,17'd36536,17'd38278,17'd38151,17'd38279,17'd38153,17'd35291,17'd31035,17'd35011,17'd28853,17'd27766,17'd28600,17'd31034,17'd24742,17'd23385,17'd23217,17'd23038,17'd22677,17'd23573,17'd32827,17'd23569,17'd32191,17'd29829,17'd23567,17'd32351,17'd29973,17'd23923,17'd23731,17'd25178,17'd27766,17'd28853,17'd31035,17'd29245,17'd29246,17'd30279,17'd32832,17'd38280,17'd38281,17'd29107,17'd32833,17'd29106,17'd29106,17'd28372,17'd28728,17'd29536,17'd30587,17'd28727,17'd28252,17'd38282,17'd28601,17'd28975,17'd24249,17'd23564,17'd30275,17'd24252,17'd25032,17'd33483,17'd25178,17'd24897,17'd34622,17'd29240,17'd24898,17'd29103,17'd28369,17'd25567,17'd28597,17'd31366,17'd30606,17'd26782,17'd28980,17'd27885,17'd28134,17'd38157,17'd37779,17'd38283,17'd38160,17'd38284,17'd36266,17'd38285,17'd37780,17'd37520,17'd33817,17'd35858,17'd38161,17'd38286,17'd38287,17'd38288,17'd38289,17'd38290,17'd27647,17'd38291,17'd36713,17'd32366,17'd29263,17'd33657,17'd33807,17'd32366,17'd28497,17'd38292,17'd38293,17'd38294,17'd38295,17'd38296,17'd38297,17'd38298,17'd38299,17'd38300,17'd38301,17'd38302,17'd38303,17'd38304,17'd38305,17'd38306,17'd38307,17'd34492,17'd38308,17'd38309,17'd10194,17'd38310,17'd38311,17'd38312,17'd38189,17'd38055,17'd37801,17'd38313,17'd20384,17'd16955,17'd22942,17'd38314,17'd38056,17'd38315,17'd38316,17'd28057,17'd27933,17'd9933,17'd9933,17'd29592,17'd27933,17'd29592,17'd9933,17'd6219,17'd28185,17'd30333,17'd31553,17'd31891,17'd6390,17'd5614,17'd5335,17'd5161,17'd4526,17'd38317,17'd5153,17'd5336,17'd7499,17'd9933,17'd28184,17'd5337,17'd38318,17'd38319,17'd38320,17'd4200,17'd38321,17'd38322,17'd38061,17'd38323,17'd38324,17'd38325,17'd38326,17'd38327,17'd38198,17'd3047,17'd38328,17'd2726,17'd38329,17'd37572,17'd38330,17'd38331,17'd38332,17'd3390,17'd5937,17'd38333,17'd38333,17'd5356,17'd38201,17'd38334,17'd38203,17'd37959,17'd37959,17'd6418,17'd7537,17'd33051,17'd35487,17'd33051,17'd33051,17'd33051,17'd35487,17'd37168,17'd37168,17'd35487,17'd2906,17'd3073,17'd5372,17'd445,17'd1401,17'd1263,17'd623,17'd1122,17'd621,17'd18515,17'd38335,17'd33848,17'd36182
},
'{
17'd4244,17'd4892,17'd6420,17'd4245,17'd14743,17'd13428,17'd3101,17'd3251,17'd3427,17'd3901,17'd3427,17'd34512,17'd14070,17'd2594,17'd466,17'd13,17'd3905,17'd3905,17'd653,17'd652,17'd287,17'd2424,17'd6902,17'd6437,17'd5803,17'd5804,17'd5211,17'd4896,17'd3912,17'd37171,17'd1705,17'd18150,17'd2949,17'd1979,17'd3437,17'd24674,17'd38336,17'd13307,17'd38337,17'd3115,17'd34351,17'd38338,17'd38339,17'd38340,17'd38341,17'd38342,17'd24194,17'd14767,17'd16411,17'd17690,17'd19008,17'd17206,17'd17689,17'd16658,17'd17940,17'd12813,17'd15516,17'd15516,17'd34180,17'd19389,17'd38343,17'd16415,17'd38344,17'd38345,17'd38346,17'd38086,17'd38087,17'd38214,17'd37717,17'd38347,17'd36761,17'd37458,17'd37834,17'd37835,17'd33864,17'd35784,17'd15023,17'd14109,17'd9164,17'd8852,17'd27962,17'd7103,17'd38096,17'd38348,17'd38349,17'd38350,17'd38350,17'd38351,17'd38094,17'd38220,17'd38220,17'd37058,17'd38352,17'd38353,17'd38354,17'd38355,17'd38356,17'd38357,17'd38358,17'd38359,17'd38360,17'd38361,17'd38362,17'd38363,17'd14136,17'd8733,17'd19923,17'd8574,17'd8573,17'd12725,17'd21208,17'd8578,17'd19535,17'd8877,17'd14674,17'd16682,17'd8884,17'd9046,17'd12722,17'd8565,17'd21984,17'd9340,17'd17847,17'd36072,17'd24538,17'd29328,17'd37065,17'd30834,17'd33568,17'd33720,17'd33568,17'd30221,17'd29067,17'd29328,17'd26371,17'd21362,17'd30532,17'd38235,17'd21503,17'd19918,17'd18332,17'd9344,17'd10335,17'd9189,17'd16910,17'd9348,17'd25677,17'd8569,17'd11404,17'd8247,17'd15429,17'd8572,17'd8728,17'd8725,17'd8881,17'd9189,17'd15569,17'd11809,17'd9742,17'd24709,17'd11400,17'd21985,17'd24031,17'd28345,17'd31295,17'd32926,17'd30531,17'd38364,17'd38108,17'd38365,17'd38366,17'd18448,17'd38367,17'd38368,17'd37071,17'd38110,17'd38369,17'd38370,17'd37987,17'd35655,17'd32452,17'd9880,17'd38371,17'd38372,17'd29081,17'd31312,17'd33896,17'd38373,17'd37747,17'd31468,17'd38374,17'd38375,17'd36647,17'd38376,17'd38377,17'd38378,17'd38379,17'd38380,17'd38381,17'd38382,17'd38383,17'd38384,17'd38385,17'd38386,17'd38387,17'd38388,17'd38389,17'd38390,17'd36105,17'd36383,17'd36243,17'd36964,17'd36668,17'd36818,17'd36963,17'd36963,17'd36668,17'd36963,17'd36668,17'd36819,17'd37634,17'd37634,17'd37367,17'd37368,17'd37367,17'd37367,17'd37368,17'd37366,17'd37096,17'd37096,17'd37495,17'd37368,17'd37368,17'd37634,17'd36669,17'd36669,17'd37368,17'd37495,17'd37367,17'd38391,17'd38261,17'd36671,17'd36105,17'd36105,17'd36104,17'd36103,17'd35972,17'd36246,17'd38392,17'd38393,17'd38394,17'd37103,17'd38395,17'd38396,17'd38397,17'd38398,17'd37770,17'd38399,17'd37894,17'd38017,17'd37244,17'd38400,17'd38273,17'd38274,17'd37899,17'd38275,17'd38401,17'd38402,17'd38403,17'd35148,17'd38278,17'd37905,17'd38279,17'd38153,17'd34275,17'd30735,17'd34637,17'd27258,17'd27766,17'd28600,17'd29101,17'd24416,17'd29529,17'd23217,17'd22678,17'd22332,17'd22332,17'd32827,17'd23569,17'd29686,17'd23387,17'd23567,17'd23215,17'd29973,17'd23388,17'd24086,17'd27637,17'd27766,17'd28853,17'd31035,17'd29245,17'd28727,17'd31503,17'd32506,17'd38404,17'd38405,17'd36848,17'd29690,17'd33486,17'd33486,17'd29248,17'd32018,17'd34285,17'd33321,17'd28727,17'd35012,17'd38406,17'd28975,17'd28852,17'd29534,17'd23565,17'd23565,17'd34467,17'd24895,17'd33483,17'd29244,17'd25030,17'd38407,17'd29240,17'd24897,17'd29103,17'd28850,17'd28369,17'd28597,17'd31366,17'd27513,17'd27259,17'd28727,17'd30279,17'd28134,17'd38408,17'd37514,17'd38283,17'd38160,17'd38409,17'd36266,17'd38285,17'd38029,17'd38030,17'd33817,17'd35858,17'd38161,17'd38286,17'd36552,17'd38410,17'd38411,17'd38412,17'd26404,17'd38413,17'd34625,17'd28605,17'd28731,17'd35714,17'd32682,17'd37405,17'd38414,17'd38415,17'd38416,17'd38417,17'd38418,17'd38419,17'd38420,17'd38421,17'd38422,17'd38423,17'd38424,17'd38425,17'd38426,17'd38427,17'd38428,17'd38429,17'd38430,17'd38431,17'd38184,17'd38432,17'd38433,17'd7001,17'd38434,17'd38435,17'd38436,17'd38055,17'd37938,17'd38437,17'd20384,17'd19222,17'd37427,17'd38438,17'd38439,17'd22943,17'd38440,17'd27934,17'd10515,17'd8780,17'd8780,17'd27815,17'd27933,17'd29592,17'd9933,17'd6219,17'd28185,17'd30333,17'd30333,17'd33369,17'd27935,17'd26949,17'd5335,17'd5161,17'd4684,17'd38441,17'd38442,17'd5335,17'd6220,17'd7668,17'd8934,17'd5616,17'd38443,17'd38444,17'd38445,17'd38446,17'd38447,17'd38448,17'd38449,17'd38450,17'd38451,17'd38452,17'd38453,17'd38454,17'd38455,17'd3047,17'd38328,17'd2726,17'd38456,17'd37572,17'd20560,17'd38457,17'd1665,17'd3390,17'd5937,17'd5496,17'd18142,17'd38458,17'd38201,17'd38334,17'd38203,17'd38459,17'd6095,17'd8507,17'd7537,17'd33051,17'd33051,17'd33051,17'd33051,17'd38460,17'd38460,17'd37168,17'd35487,17'd12923,17'd2906,17'd5958,17'd4085,17'd445,17'd1261,17'd1263,17'd427,17'd609,17'd635,17'd440,17'd35617,17'd35062,17'd38461
},
'{
17'd4244,17'd4892,17'd6420,17'd4245,17'd14743,17'd13428,17'd3101,17'd2934,17'd3901,17'd3901,17'd3427,17'd3251,17'd14070,17'd2594,17'd2,17'd13,17'd3905,17'd3905,17'd653,17'd652,17'd287,17'd2424,17'd6902,17'd6437,17'd5803,17'd5804,17'd5212,17'd4580,17'd2948,17'd37171,17'd1705,17'd38462,17'd2949,17'd1979,17'd3437,17'd32731,17'd32255,17'd13307,17'd38337,17'd38463,17'd34351,17'd38464,17'd37711,17'd38465,17'd38466,17'd38342,17'd24194,17'd14767,17'd16411,17'd17445,17'd19255,17'd17206,17'd17689,17'd12531,17'd24347,17'd33858,17'd12813,17'd11359,17'd35777,17'd19263,17'd38467,17'd38468,17'd38469,17'd38470,17'd38471,17'd38086,17'd38087,17'd38472,17'd37717,17'd38473,17'd38474,17'd38475,17'd37834,17'd35358,17'd38476,17'd17330,17'd14904,17'd14109,17'd9015,17'd38477,17'd38478,17'd38479,17'd38480,17'd38481,17'd38349,17'd38482,17'd38350,17'd38350,17'd38351,17'd38483,17'd38484,17'd37184,17'd38353,17'd38485,17'd38486,17'd38487,17'd38488,17'd37726,17'd38489,17'd38490,17'd38491,17'd38492,17'd38493,17'd38494,17'd11968,17'd19780,17'd21208,17'd8574,17'd8413,17'd13139,17'd19780,17'd25679,17'd25532,17'd8877,17'd15807,17'd38495,17'd8885,17'd9195,17'd17237,17'd38496,17'd21984,17'd13370,17'd29335,17'd38497,17'd26149,17'd30673,17'd37065,17'd33718,17'd31287,17'd38498,17'd33568,17'd30676,17'd31940,17'd27984,17'd26149,17'd24858,17'd38499,17'd38235,17'd21503,17'd9885,17'd9480,17'd9344,17'd10173,17'd9743,17'd15682,17'd9044,17'd9194,17'd8886,17'd9886,17'd9744,17'd15429,17'd8571,17'd8569,17'd8881,17'd16910,17'd9189,17'd15569,17'd18556,17'd38236,17'd13522,17'd15176,17'd18327,17'd24538,17'd28345,17'd31295,17'd38500,17'd31135,17'd38501,17'd29644,17'd38502,17'd38366,17'd18448,17'd38503,17'd30086,17'd32773,17'd38110,17'd30841,17'd38370,17'd37987,17'd35243,17'd34200,17'd9880,17'd38241,17'd29663,17'd38504,17'd38505,17'd38506,17'd31971,17'd37992,17'd37867,17'd38374,17'd38507,17'd38508,17'd38509,17'd38510,17'd38511,17'd38512,17'd38513,17'd38514,17'd38123,17'd38515,17'd38516,17'd38517,17'd38518,17'd38519,17'd38520,17'd37367,17'd36820,17'd36668,17'd36660,17'd36383,17'd36105,17'd36660,17'd36818,17'd38130,17'd37883,17'd37883,17'd38007,17'd38007,17'd38130,17'd37095,17'd37096,17'd37495,17'd37096,17'd37495,17'd37366,17'd37368,17'd37368,17'd37368,17'd37366,17'd37366,17'd37366,17'd37367,17'd37368,17'd37368,17'd37634,17'd37634,17'd37368,17'd37368,17'd37367,17'd38521,17'd36243,17'd36105,17'd36105,17'd36104,17'd36103,17'd35972,17'd36245,17'd35684,17'd38393,17'd38522,17'd38523,17'd38524,17'd38525,17'd38526,17'd38527,17'd38528,17'd38529,17'd38530,17'd38531,17'd38020,17'd38532,17'd38273,17'd38274,17'd37899,17'd38533,17'd38534,17'd38535,17'd38403,17'd35286,17'd38278,17'd37905,17'd38536,17'd38153,17'd34451,17'd30735,17'd33163,17'd27258,17'd27766,17'd28600,17'd28850,17'd24744,17'd29526,17'd29828,17'd22679,17'd22332,17'd22678,17'd32827,17'd23388,17'd29686,17'd23387,17'd23567,17'd23215,17'd29973,17'd23388,17'd24086,17'd27637,17'd27766,17'd27258,17'd31035,17'd28727,17'd38537,17'd29977,17'd32506,17'd38404,17'd38405,17'd29537,17'd29690,17'd33486,17'd33486,17'd29248,17'd36989,17'd34285,17'd33654,17'd31035,17'd38538,17'd33318,17'd23563,17'd23563,17'd29534,17'd34137,17'd34137,17'd34467,17'd24744,17'd32353,17'd31034,17'd25180,17'd27763,17'd29240,17'd24897,17'd29103,17'd25317,17'd28597,17'd33000,17'd31366,17'd30734,17'd27640,17'd28979,17'd30279,17'd32354,17'd38408,17'd37514,17'd38283,17'd38160,17'd38409,17'd36266,17'd38285,17'd37780,17'd38539,17'd37911,17'd35858,17'd33955,17'd38540,17'd27030,17'd38541,17'd38542,17'd38543,17'd38544,17'd28867,17'd35733,17'd33808,17'd29127,17'd35714,17'd38545,17'd32682,17'd38546,17'd38547,17'd38548,17'd35434,17'd38549,17'd38550,17'd38551,17'd38552,17'd38553,17'd38554,17'd38555,17'd19431,17'd38556,17'd38557,17'd38558,17'd38559,17'd38560,17'd38561,17'd38562,17'd38309,17'd8908,17'd8286,17'd38563,17'd38564,17'd38565,17'd38055,17'd37939,17'd38566,17'd20384,17'd19222,17'd37427,17'd38438,17'd38438,17'd22767,17'd36031,17'd27934,17'd28183,17'd27815,17'd9933,17'd29592,17'd27933,17'd29592,17'd9933,17'd6220,17'd28185,17'd30333,17'd30333,17'd32718,17'd27935,17'd26949,17'd5335,17'd5161,17'd4684,17'd38441,17'd33532,17'd5160,17'd6219,17'd7499,17'd8780,17'd5763,17'd38567,17'd38568,17'd38569,17'd38570,17'd38571,17'd38572,17'd38449,17'd38450,17'd3537,17'd38573,17'd3360,17'd38574,17'd38575,17'd38576,17'd38328,17'd2726,17'd38456,17'd37572,17'd38577,17'd38578,17'd1665,17'd3390,17'd38579,17'd5495,17'd18142,17'd11048,17'd38458,17'd38202,17'd38580,17'd38581,17'd37959,17'd6418,17'd7537,17'd33051,17'd33051,17'd34002,17'd33051,17'd38460,17'd38460,17'd37168,17'd35487,17'd11882,17'd5183,17'd4882,17'd4085,17'd445,17'd1261,17'd1263,17'd443,17'd1122,17'd636,17'd28065,17'd35617,17'd35062,17'd38461
},
'{
17'd4892,17'd4892,17'd6420,17'd14743,17'd13428,17'd13428,17'd3101,17'd3101,17'd3427,17'd3901,17'd3427,17'd3251,17'd14070,17'd4247,17'd2,17'd13,17'd20404,17'd20404,17'd653,17'd28,17'd287,17'd9275,17'd6903,17'd6437,17'd5803,17'd5804,17'd5212,17'd38582,17'd3912,17'd37171,17'd1139,17'd38462,17'd2949,17'd1979,17'd3437,17'd24674,17'd38336,17'd38583,17'd38337,17'd38584,17'd26017,17'd38585,17'd38586,17'd38587,17'd38466,17'd38588,17'd32101,17'd14768,17'd16169,17'd17207,17'd18656,17'd27461,17'd19128,17'd30058,17'd38589,17'd38590,17'd11475,17'd36757,17'd38591,17'd38592,17'd38593,17'd38594,17'd38595,17'd38596,17'd38597,17'd38598,17'd38087,17'd38599,17'd38600,17'd38473,17'd38474,17'd38475,17'd38601,17'd35216,17'd33070,17'd35920,17'd12822,17'd14109,17'd9015,17'd38477,17'd38478,17'd38479,17'd38092,17'd38602,17'd38349,17'd38482,17'd38603,17'd38093,17'd38604,17'd38602,17'd38605,17'd37184,17'd38606,17'd38607,17'd38608,17'd38609,17'd38610,17'd38611,17'd38612,17'd38613,17'd38614,17'd38615,17'd38616,17'd38617,17'd10860,17'd10028,17'd8248,17'd15945,17'd8414,17'd35094,17'd8249,17'd11138,17'd14004,17'd8877,17'd15807,17'd35088,17'd17607,17'd9046,17'd20453,17'd38618,17'd21984,17'd9620,17'd10331,17'd38619,17'd28110,17'd28462,17'd32282,17'd31941,17'd33568,17'd33568,17'd31941,17'd30676,17'd29924,17'd27984,17'd24538,17'd20609,17'd29789,17'd27487,17'd16796,17'd10856,17'd10742,17'd9480,17'd9340,17'd9191,17'd9189,17'd8720,17'd9194,17'd9040,17'd8726,17'd9482,17'd8409,17'd10607,17'd8877,17'd17237,17'd26874,17'd8874,17'd15569,17'd11809,17'd17965,17'd19278,17'd10476,17'd17478,17'd26493,17'd28462,17'd30074,17'd30225,17'd30978,17'd38366,17'd29644,17'd29644,17'd38501,17'd18448,17'd17234,17'd35520,17'd38620,17'd31141,17'd33419,17'd38621,17'd36078,17'd38622,17'd34034,17'd27619,17'd29667,17'd30103,17'd31466,17'd38623,17'd38624,17'd38625,17'd37866,17'd36225,17'd38626,17'd38627,17'd38628,17'd37752,17'd38629,17'd38630,17'd38631,17'd38632,17'd38633,17'd38634,17'd38635,17'd38636,17'd38637,17'd38638,17'd38639,17'd38640,17'd38392,17'd34428,17'd34859,17'd38641,17'd38642,17'd38643,17'd38644,17'd33916,17'd33769,17'd35274,17'd36247,17'd38645,17'd36670,17'd37368,17'd37230,17'd37230,17'd37093,17'd38646,17'd37095,17'd37096,17'd37096,17'd37495,17'd37366,17'd37366,17'd37366,17'd37366,17'd37368,17'd37368,17'd37368,17'd37634,17'd36669,17'd37634,17'd37367,17'd37368,17'd37097,17'd36964,17'd36383,17'd38647,17'd38648,17'd36104,17'd36385,17'd35962,17'd38649,17'd35971,17'd38650,17'd38651,17'd38652,17'd38653,17'd38654,17'd38655,17'd37240,17'd36976,17'd38656,17'd38657,17'd38658,17'd38659,17'd38273,17'd38400,17'd37900,17'd38660,17'd38534,17'd38661,17'd38662,17'd36685,17'd38663,17'd38664,17'd38665,17'd38153,17'd36983,17'd30735,17'd30586,17'd28853,17'd26062,17'd28594,17'd28850,17'd24744,17'd29685,17'd23215,17'd22331,17'd22332,17'd22680,17'd32827,17'd23388,17'd29826,17'd29530,17'd23567,17'd32351,17'd23216,17'd23388,17'd24086,17'd28254,17'd27766,17'd27258,17'd31035,17'd28979,17'd28726,17'd27642,17'd32506,17'd38666,17'd38404,17'd29537,17'd29690,17'd33486,17'd32507,17'd32505,17'd32018,17'd34114,17'd33654,17'd31035,17'd38538,17'd38667,17'd29532,17'd29532,17'd29375,17'd38668,17'd38669,17'd24089,17'd38670,17'd33969,17'd33345,17'd29976,17'd28595,17'd29240,17'd24896,17'd31034,17'd29101,17'd27882,17'd33000,17'd31366,17'd38671,17'd27640,17'd28979,17'd30279,17'd32354,17'd38672,17'd37514,17'd38673,17'd38160,17'd38409,17'd36266,17'd38285,17'd38539,17'd38674,17'd37911,17'd35858,17'd38675,17'd38676,17'd28735,17'd38677,17'd38543,17'd35577,17'd38678,17'd33968,17'd38679,17'd38680,17'd29110,17'd38681,17'd31362,17'd38682,17'd38683,17'd29851,17'd32370,17'd26905,17'd36698,17'd38684,17'd38685,17'd38686,17'd38687,17'd38688,17'd38689,17'd19431,17'd38690,17'd38691,17'd38692,17'd28163,17'd37793,17'd38693,17'd21282,17'd38694,17'd11689,17'd38695,17'd38696,17'd38697,17'd38698,17'd38699,17'd37938,17'd38700,17'd20250,17'd18970,17'd37427,17'd38438,17'd38438,17'd37427,17'd38701,17'd27934,17'd10642,17'd28184,17'd8780,17'd10515,17'd27933,17'd29592,17'd9933,17'd6220,17'd30638,17'd25627,17'd30333,17'd32718,17'd28185,17'd5762,17'd5330,17'd5161,17'd4847,17'd38702,17'd38058,17'd5329,17'd6219,17'd7499,17'd7669,17'd5764,17'd38703,17'd38704,17'd4200,17'd38705,17'd38706,17'd38707,17'd38449,17'd38450,17'd38708,17'd38709,17'd38710,17'd38711,17'd38712,17'd36898,17'd38328,17'd38713,17'd38329,17'd2388,17'd19730,17'd38714,17'd38715,17'd38716,17'd38717,17'd38718,17'd5495,17'd11048,17'd38458,17'd38202,17'd37957,17'd37709,17'd4868,17'd35769,17'd7537,17'd33051,17'd34002,17'd34002,17'd33051,17'd38460,17'd38460,17'd38719,17'd33051,17'd11882,17'd5183,17'd4882,17'd3391,17'd445,17'd1261,17'd1262,17'd427,17'd609,17'd636,17'd38720,17'd618,17'd33540,17'd36047
},
'{
17'd4892,17'd4428,17'd6420,17'd4245,17'd14743,17'd14743,17'd3101,17'd2934,17'd3427,17'd3901,17'd3427,17'd3251,17'd14070,17'd4247,17'd2,17'd13,17'd3905,17'd20404,17'd653,17'd28,17'd287,17'd9275,17'd6903,17'd6437,17'd5803,17'd5804,17'd5054,17'd38721,17'd2948,17'd37171,17'd1139,17'd38722,17'd2949,17'd1979,17'd3266,17'd32731,17'd32255,17'd38723,17'd13955,17'd38724,17'd38725,17'd4274,17'd38726,17'd38727,17'd38728,17'd35625,17'd32101,17'd14768,17'd16169,17'd17207,17'd17206,17'd18655,17'd19006,17'd38729,17'd34181,17'd38730,17'd38731,17'd36329,17'd38732,17'd38733,17'd15906,17'd38734,17'd38735,17'd38346,17'd38597,17'd38598,17'd38087,17'd38472,17'd37718,17'd38473,17'd38474,17'd38736,17'd38737,17'd34191,17'd35217,17'd35920,17'd14109,17'd9164,17'd9016,17'd8852,17'd7760,17'd38479,17'd38220,17'd38738,17'd38739,17'd38482,17'd38603,17'd6645,17'd38093,17'd38602,17'd38605,17'd38352,17'd38606,17'd38740,17'd38741,17'd38742,17'd38743,17'd38744,17'd38745,17'd38746,17'd38747,17'd6804,17'd6968,17'd38494,17'd10860,17'd10028,17'd8248,17'd15945,17'd12865,17'd38748,17'd8249,17'd9196,17'd12723,17'd16067,17'd15807,17'd9190,17'd17607,17'd16205,17'd12264,17'd38749,17'd21984,17'd11136,17'd29335,17'd14382,17'd26371,17'd30370,17'd32282,17'd31941,17'd34203,17'd33568,17'd31941,17'd30676,17'd29924,17'd26873,17'd24992,17'd30230,17'd29790,17'd27487,17'd17719,17'd9739,17'd9741,17'd9480,17'd9340,17'd23853,17'd9346,17'd9189,17'd8873,17'd9194,17'd8879,17'd9482,17'd8726,17'd8724,17'd8877,17'd15297,17'd16910,17'd8874,17'd16065,17'd15566,17'd17841,17'd17847,17'd11399,17'd16442,17'd24856,17'd28462,17'd29780,17'd29483,17'd38365,17'd28349,17'd29644,17'd38750,17'd38751,17'd17844,17'd38239,17'd31602,17'd38620,17'd31141,17'd38752,17'd21670,17'd36787,17'd32451,17'd34034,17'd38753,17'd30251,17'd31612,17'd38754,17'd38755,17'd38756,17'd38757,17'd36497,17'd38758,17'd38759,17'd38760,17'd38761,17'd38762,17'd38763,17'd38764,17'd38120,17'd38765,17'd38766,17'd38767,17'd38768,17'd38769,17'd38257,17'd38770,17'd38771,17'd38772,17'd38773,17'd38774,17'd38775,17'd38776,17'd38777,17'd38778,17'd38779,17'd38780,17'd38781,17'd38782,17'd38783,17'd38784,17'd38785,17'd38786,17'd36523,17'd38787,17'd35963,17'd35551,17'd37096,17'd37095,17'd37230,17'd37230,17'd37096,17'd37495,17'd37366,17'd37368,17'd37495,17'd37367,17'd36669,17'd36669,17'd36669,17'd36669,17'd37634,17'd37368,17'd36963,17'd37097,17'd37226,17'd38788,17'd38647,17'd36104,17'd36384,17'd35962,17'd38789,17'd35972,17'd38790,17'd38791,17'd38792,17'd38793,17'd38794,17'd38795,17'd38796,17'd38797,17'd37893,17'd38798,17'd38799,17'd38659,17'd38800,17'd38400,17'd38020,17'd38801,17'd38802,17'd38803,17'd38804,17'd36685,17'd38663,17'd38664,17'd36686,17'd38805,17'd34450,17'd35011,17'd30586,17'd28853,17'd28481,17'd27765,17'd27511,17'd24416,17'd30278,17'd23215,17'd22331,17'd23038,17'd22331,17'd30425,17'd23387,17'd23386,17'd35865,17'd38806,17'd32351,17'd23216,17'd23387,17'd30879,17'd28719,17'd27766,17'd27258,17'd31035,17'd28486,17'd28726,17'd27642,17'd32506,17'd38807,17'd38404,17'd29537,17'd29690,17'd33486,17'd32507,17'd32355,17'd37250,17'd29107,17'd33654,17'd28979,17'd25565,17'd38808,17'd29971,17'd29971,17'd29527,17'd31664,17'd38809,17'd38810,17'd38811,17'd25710,17'd38812,17'd29976,17'd34283,17'd29240,17'd24896,17'd31034,17'd25317,17'd28597,17'd33000,17'd31366,17'd33507,17'd27883,17'd28979,17'd30279,17'd32354,17'd38672,17'd38813,17'd38673,17'd38160,17'd38409,17'd36266,17'd38814,17'd38815,17'd38539,17'd38030,17'd33806,17'd38675,17'd38816,17'd28735,17'd38817,17'd38818,17'd35577,17'd23916,17'd38819,17'd38820,17'd38821,17'd31847,17'd33657,17'd31515,17'd38822,17'd38823,17'd38824,17'd38825,17'd38826,17'd38827,17'd38828,17'd34316,17'd38686,17'd25573,17'd38829,17'd38830,17'd38831,17'd38832,17'd38833,17'd38834,17'd38835,17'd38836,17'd38837,17'd38838,17'd38839,17'd31241,17'd8139,17'd38840,17'd38841,17'd38842,17'd38699,17'd37938,17'd38843,17'd22251,17'd19479,17'd37555,17'd38844,17'd38438,17'd38845,17'd36310,17'd27934,17'd28183,17'd27815,17'd27815,17'd10515,17'd27933,17'd29592,17'd9933,17'd6220,17'd30638,17'd25627,17'd25627,17'd32553,17'd28185,17'd5762,17'd5160,17'd5163,17'd4847,17'd38702,17'd38846,17'd27570,17'd5614,17'd7499,17'd8780,17'd5763,17'd38847,17'd38848,17'd4199,17'd38849,17'd38850,17'd4201,17'd3846,17'd38851,17'd38852,17'd38853,17'd38710,17'd38854,17'd38712,17'd38576,17'd38328,17'd38855,17'd21322,17'd19237,17'd20127,17'd18631,17'd36181,17'd38856,17'd38857,17'd38858,17'd5495,17'd11048,17'd38458,17'd38859,17'd38860,17'd38861,17'd38459,17'd6417,17'd7537,17'd38460,17'd34002,17'd34002,17'd33051,17'd38460,17'd38460,17'd38719,17'd33051,17'd11882,17'd5183,17'd4882,17'd3391,17'd445,17'd1261,17'd1262,17'd232,17'd234,17'd38862,17'd38863,17'd19240,17'd33376,17'd35618
},
'{
17'd25384,17'd6420,17'd4245,17'd4245,17'd4245,17'd4733,17'd4245,17'd25384,17'd6420,17'd6420,17'd3251,17'd38864,17'd27714,17'd4247,17'd17,17'd3905,17'd3905,17'd3905,17'd1278,17'd980,17'd7061,17'd7728,17'd7225,17'd6437,17'd6598,17'd5379,17'd4894,17'd2605,17'd38865,17'd37171,17'd35772,17'd1560,17'd3436,17'd3437,17'd38866,17'd2950,17'd38867,17'd38868,17'd27717,17'd21336,17'd25796,17'd38869,17'd38870,17'd38871,17'd38872,17'd34520,17'd14893,17'd16168,17'd16034,17'd20425,17'd19891,17'd17941,17'd27217,17'd34675,17'd38873,17'd38874,17'd38875,17'd18537,17'd38876,17'd38877,17'd38878,17'd38595,17'd38596,17'd38879,17'd38880,17'd38881,17'd38882,17'd38883,17'd36466,17'd38473,17'd38884,17'd38885,17'd38886,17'd32423,17'd15399,17'd14230,17'd12822,17'd9164,17'd8851,17'd38218,17'd38887,17'd38888,17'd38889,17'd38739,17'd38890,17'd38890,17'd6645,17'd6645,17'd38891,17'd38349,17'd38604,17'd37320,17'd38892,17'd38893,17'd38894,17'd38895,17'd38896,17'd38897,17'd38898,17'd38899,17'd38900,17'd38901,17'd38902,17'd38903,17'd10179,17'd17483,17'd8249,17'd9196,17'd12865,17'd13003,17'd17126,17'd8413,17'd8726,17'd9194,17'd24361,17'd10175,17'd38904,17'd38905,17'd15945,17'd8409,17'd9191,17'd24709,17'd11669,17'd14259,17'd38906,17'd37733,17'd37065,17'd31941,17'd34835,17'd34835,17'd31941,17'd31439,17'd30370,17'd26872,17'd21505,17'd11396,17'd28352,17'd10328,17'd17719,17'd9883,17'd10024,17'd9885,17'd10743,17'd10857,17'd10743,17'd9346,17'd9043,17'd16067,17'd8569,17'd9482,17'd8725,17'd8886,17'd9194,17'd9045,17'd9043,17'd15180,17'd24037,17'd12116,17'd11671,17'd19280,17'd38499,17'd24995,17'd25925,17'd30077,17'd38907,17'd30979,17'd38108,17'd38908,17'd38108,17'd38909,17'd38910,17'd38911,17'd30234,17'd37071,17'd31603,17'd38912,17'd30841,17'd37741,17'd37860,17'd38913,17'd10161,17'd32778,17'd38914,17'd38915,17'd38916,17'd38917,17'd38918,17'd38919,17'd36225,17'd38920,17'd38921,17'd38922,17'd38923,17'd38924,17'd38925,17'd38926,17'd38927,17'd38928,17'd38929,17'd38930,17'd38931,17'd38932,17'd38933,17'd38934,17'd38935,17'd38936,17'd38937,17'd38938,17'd38939,17'd38940,17'd38941,17'd38942,17'd38943,17'd38944,17'd38945,17'd38946,17'd38947,17'd38947,17'd38948,17'd38949,17'd38950,17'd38951,17'd38952,17'd38953,17'd38954,17'd34425,17'd36387,17'd36515,17'd36962,17'd38955,17'd38956,17'd36962,17'd37228,17'd36661,17'd37366,17'd36670,17'd36670,17'd37367,17'd36813,17'd36669,17'd37366,17'd37368,17'd37097,17'd36964,17'd38957,17'd38648,17'd36105,17'd35683,17'd35684,17'd38958,17'd38959,17'd38960,17'd38961,17'd38962,17'd38963,17'd38964,17'd38655,17'd38965,17'd38966,17'd38967,17'd38968,17'd38659,17'd38969,17'd38400,17'd37899,17'd38660,17'd38965,17'd38970,17'd38971,17'd38972,17'd38973,17'd37905,17'd37508,17'd38974,17'd38975,17'd32185,17'd26902,17'd28725,17'd27767,17'd27765,17'd25320,17'd32659,17'd38976,17'd36986,17'd22330,17'd22678,17'd22329,17'd29973,17'd23923,17'd29376,17'd23736,17'd38806,17'd32008,17'd23216,17'd23566,17'd29100,17'd33484,17'd26062,17'd27146,17'd34637,17'd30586,17'd28486,17'd27642,17'd35707,17'd38807,17'd38977,17'd29537,17'd29690,17'd29106,17'd29380,17'd32355,17'd32505,17'd29248,17'd32017,17'd29246,17'd25565,17'd38978,17'd38979,17'd29830,17'd38980,17'd24094,17'd35455,17'd23921,17'd38811,17'd25029,17'd29101,17'd30432,17'd24745,17'd28718,17'd24896,17'd27511,17'd28484,17'd28597,17'd33000,17'd31520,17'd31055,17'd27514,17'd28486,17'd31503,17'd27885,17'd37514,17'd38813,17'd38981,17'd38982,17'd38983,17'd38409,17'd38984,17'd38985,17'd38986,17'd38987,17'd37265,17'd37405,17'd38676,17'd35300,17'd38988,17'd31358,17'd25439,17'd24090,17'd28851,17'd29548,17'd38989,17'd31364,17'd28375,17'd38822,17'd38990,17'd38991,17'd38992,17'd38993,17'd29701,17'd38994,17'd38995,17'd24747,17'd38552,17'd38996,17'd38997,17'd38998,17'd34319,17'd38999,17'd39000,17'd39001,17'd39002,17'd39003,17'd23612,17'd22728,17'd21124,17'd39004,17'd39005,17'd39006,17'd39007,17'd39008,17'd39009,17'd39010,17'd38437,17'd38313,17'd22089,17'd39011,17'd39012,17'd38056,17'd39013,17'd39014,17'd35340,17'd31551,17'd31888,17'd29593,17'd27815,17'd10515,17'd31243,17'd29593,17'd6220,17'd27935,17'd5160,17'd25627,17'd30637,17'd25627,17'd5762,17'd5160,17'd5163,17'd4847,17'd33533,17'd33534,17'd4688,17'd5335,17'd9091,17'd29740,17'd37289,17'd39015,17'd39016,17'd39017,17'd39018,17'd39019,17'd4201,17'd39020,17'd39021,17'd3537,17'd39022,17'd39023,17'd39024,17'd39025,17'd38067,17'd39026,17'd2364,17'd39027,17'd39028,17'd39029,17'd23642,17'd39030,17'd39031,17'd4710,17'd4553,17'd4865,17'd39032,17'd11048,17'd39033,17'd38334,17'd37958,17'd38459,17'd6418,17'd7537,17'd9124,17'd9124,17'd9124,17'd38460,17'd33051,17'd33051,17'd31562,17'd28066,17'd33050,17'd6721,17'd1946,17'd5371,17'd1261,17'd1261,17'd446,17'd623,17'd234,17'd955,17'd39034,17'd39035,17'd39036,17'd39037
},
'{
17'd25384,17'd6420,17'd4245,17'd6420,17'd4245,17'd4733,17'd4245,17'd25384,17'd6420,17'd6420,17'd3251,17'd38864,17'd27714,17'd4247,17'd17,17'd17,17'd3905,17'd3905,17'd1278,17'd980,17'd7385,17'd7385,17'd7225,17'd6437,17'd6598,17'd5379,17'd4894,17'd2606,17'd38865,17'd1841,17'd35772,17'd1708,17'd3436,17'd3437,17'd1288,17'd39038,17'd38867,17'd29899,17'd2959,17'd39039,17'd5071,17'd38869,17'd39040,17'd39041,17'd38872,17'd39042,17'd17691,17'd16411,17'd17445,17'd17572,17'd19891,17'd18412,17'd11628,17'd37581,17'd37453,17'd39043,17'd35778,17'd39044,17'd38877,17'd39045,17'd39046,17'd39047,17'd38346,17'd39048,17'd39049,17'd38882,17'd38882,17'd39050,17'd39051,17'd38473,17'd38884,17'd39052,17'd39053,17'd36616,17'd35784,17'd14230,17'd14109,17'd9015,17'd8852,17'd8547,17'd39054,17'd39055,17'd39056,17'd38739,17'd38890,17'd38890,17'd39057,17'd6645,17'd39058,17'd38891,17'd38604,17'd37320,17'd38892,17'd39059,17'd39060,17'd39061,17'd39062,17'd39063,17'd39064,17'd39065,17'd6801,17'd39066,17'd39067,17'd38903,17'd10179,17'd17352,17'd10028,17'd9196,17'd12865,17'd8100,17'd9349,17'd8572,17'd10027,17'd9194,17'd24361,17'd10175,17'd38904,17'd24547,17'd9196,17'd12723,17'd9191,17'd10168,17'd28463,17'd24363,17'd39068,17'd37733,17'd32919,17'd31941,17'd34381,17'd34835,17'd31941,17'd31439,17'd30370,17'd29065,17'd24363,17'd24029,17'd24996,17'd10328,17'd17719,17'd9883,17'd10024,17'd10169,17'd10992,17'd9341,17'd9885,17'd9620,17'd9189,17'd9038,17'd9348,17'd9482,17'd8879,17'd17607,17'd10336,17'd9043,17'd9192,17'd9345,17'd9619,17'd12116,17'd9883,17'd13647,17'd39069,17'd24995,17'd26036,17'd27485,17'd29649,17'd30836,17'd39070,17'd39071,17'd38364,17'd38501,17'd17844,17'd39072,17'd39073,17'd31778,17'd37342,17'd33419,17'd38752,17'd29655,17'd34050,17'd39074,17'd29470,17'd29210,17'd39075,17'd34714,17'd39076,17'd39077,17'd36224,17'd35662,17'd39078,17'd39079,17'd35531,17'd39080,17'd39081,17'd39082,17'd39083,17'd39084,17'd39085,17'd39086,17'd39087,17'd39088,17'd39089,17'd39090,17'd39091,17'd39092,17'd39093,17'd39094,17'd39095,17'd39096,17'd39097,17'd39098,17'd39099,17'd39100,17'd39101,17'd39102,17'd39103,17'd39104,17'd39105,17'd39106,17'd39107,17'd39108,17'd39109,17'd33281,17'd39110,17'd39111,17'd39112,17'd39113,17'd39114,17'd39115,17'd34859,17'd35405,17'd36961,17'd38129,17'd37094,17'd37366,17'd37366,17'd37634,17'd36384,17'd36244,17'd39116,17'd38391,17'd38006,17'd38006,17'd36819,17'd36964,17'd38788,17'd38647,17'd36105,17'd36105,17'd36246,17'd38958,17'd39117,17'd39118,17'd39119,17'd39120,17'd39121,17'd39122,17'd39123,17'd38796,17'd39124,17'd39125,17'd39126,17'd38659,17'd38969,17'd38400,17'd37899,17'd38660,17'd38796,17'd39127,17'd39128,17'd39129,17'd37904,17'd39130,17'd37508,17'd38974,17'd38975,17'd32185,17'd26902,17'd26782,17'd27767,17'd25567,17'd25320,17'd30431,17'd29973,17'd22331,17'd22330,17'd39131,17'd23218,17'd29973,17'd23387,17'd29099,17'd23736,17'd23567,17'd32351,17'd37117,17'd29242,17'd28601,17'd33000,17'd27514,17'd27372,17'd33163,17'd26902,17'd26901,17'd31353,17'd35707,17'd38807,17'd38977,17'd29537,17'd30884,17'd29106,17'd29380,17'd32355,17'd32505,17'd32018,17'd32017,17'd28980,17'd27766,17'd33652,17'd39132,17'd37386,17'd39133,17'd34759,17'd30729,17'd39134,17'd33339,17'd28974,17'd29101,17'd32353,17'd24895,17'd24417,17'd24896,17'd27511,17'd25317,17'd28597,17'd33000,17'd33484,17'd32669,17'd27514,17'd28486,17'd31503,17'd27885,17'd37514,17'd38813,17'd38981,17'd38982,17'd38983,17'd39135,17'd35167,17'd34633,17'd39136,17'd38987,17'd37265,17'd38546,17'd35433,17'd35300,17'd39137,17'd33180,17'd24088,17'd29100,17'd24416,17'd24895,17'd39138,17'd39139,17'd30902,17'd38991,17'd38990,17'd39140,17'd27517,17'd35876,17'd39141,17'd39142,17'd39143,17'd39144,17'd39145,17'd39146,17'd39147,17'd39148,17'd39149,17'd39150,17'd39151,17'd36723,17'd38835,17'd39003,17'd21598,17'd39152,17'd39153,17'd39154,17'd39155,17'd39156,17'd39157,17'd39158,17'd39159,17'd39160,17'd22417,17'd38566,17'd22089,17'd39011,17'd39161,17'd39162,17'd39013,17'd39163,17'd34922,17'd31551,17'd39164,17'd29593,17'd10515,17'd10642,17'd30933,17'd31243,17'd9091,17'd27935,17'd25627,17'd5004,17'd4842,17'd5002,17'd5336,17'd30638,17'd5165,17'd37153,17'd33533,17'd39165,17'd39166,17'd5330,17'd9091,17'd29740,17'd5763,17'd28778,17'd39167,17'd4194,17'd39168,17'd39169,17'd38571,17'd39170,17'd39171,17'd3537,17'd39172,17'd39173,17'd39174,17'd39175,17'd37039,17'd39026,17'd2368,17'd39027,17'd39028,17'd39029,17'd39176,17'd39177,17'd39178,17'd4227,17'd39179,17'd39180,17'd10906,17'd39181,17'd38859,17'd39182,17'd39183,17'd38861,17'd15484,17'd7364,17'd9124,17'd7538,17'd7538,17'd38460,17'd33051,17'd33051,17'd31562,17'd28066,17'd33050,17'd5631,17'd5940,17'd5371,17'd1261,17'd1261,17'd446,17'd623,17'd1122,17'd792,17'd1238,17'd435,17'd39184,17'd32252
},
'{
17'd6420,17'd6420,17'd4245,17'd6420,17'd4245,17'd4245,17'd4245,17'd25384,17'd6420,17'd4245,17'd3251,17'd38864,17'd27714,17'd1127,17'd17,17'd3905,17'd3905,17'd3905,17'd1278,17'd980,17'd7385,17'd7385,17'd7225,17'd6437,17'd5804,17'd5210,17'd4894,17'd2431,17'd38865,17'd37171,17'd3598,17'd24830,17'd3600,17'd3437,17'd1288,17'd836,17'd2619,17'd29899,17'd2959,17'd39039,17'd5071,17'd36326,17'd39040,17'd39185,17'd38872,17'd39042,17'd17691,17'd16411,17'd17320,17'd18656,17'd19511,17'd11362,17'd12680,17'd39043,17'd37176,17'd39186,17'd18780,17'd39187,17'd39188,17'd39189,17'd39190,17'd39191,17'd39191,17'd39192,17'd39049,17'd38882,17'd38882,17'd39193,17'd38089,17'd36467,17'd39194,17'd39195,17'd39196,17'd15535,17'd35920,17'd13104,17'd14109,17'd9014,17'd39197,17'd8547,17'd39198,17'd39199,17'd38889,17'd38739,17'd38349,17'd38890,17'd39057,17'd39057,17'd39200,17'd38891,17'd38604,17'd39201,17'd38604,17'd39059,17'd39060,17'd39202,17'd39203,17'd39063,17'd39204,17'd39205,17'd39206,17'd39207,17'd39208,17'd7456,17'd10179,17'd17483,17'd8249,17'd9196,17'd8578,17'd12867,17'd17481,17'd10607,17'd12118,17'd9194,17'd14811,17'd26498,17'd38904,17'd24547,17'd8578,17'd8409,17'd9339,17'd10167,17'd11668,17'd29488,17'd39209,17'd39210,17'd32919,17'd31941,17'd34381,17'd34381,17'd30834,17'd39211,17'd30071,17'd24856,17'd21361,17'd19533,17'd24996,17'd10328,17'd10329,17'd10330,17'd9884,17'd10169,17'd9885,17'd11136,17'd9741,17'd10742,17'd12117,17'd9188,17'd8567,17'd30522,17'd8878,17'd24212,17'd17480,17'd9189,17'd9347,17'd25525,17'd24037,17'd12116,17'd9883,17'd19532,17'd19533,17'd24995,17'd18084,17'd28234,17'd30679,17'd28349,17'd39212,17'd39071,17'd38364,17'd39213,17'd39214,17'd39215,17'd33579,17'd32773,17'd31778,17'd30088,17'd39216,17'd33420,17'd32612,17'd39074,17'd33422,17'd39217,17'd39218,17'd39219,17'd39220,17'd39221,17'd39222,17'd37478,17'd31627,17'd39223,17'd39224,17'd34062,17'd33121,17'd37870,17'd39225,17'd39226,17'd39227,17'd39228,17'd39229,17'd39230,17'd39231,17'd39232,17'd39233,17'd39234,17'd39235,17'd39236,17'd39237,17'd39238,17'd39239,17'd39240,17'd39241,17'd39242,17'd39243,17'd39244,17'd39245,17'd39246,17'd39247,17'd39248,17'd39249,17'd39250,17'd39251,17'd39252,17'd39253,17'd39254,17'd39255,17'd39256,17'd39257,17'd39258,17'd39259,17'd33451,17'd35544,17'd35684,17'd37366,17'd37231,17'd39260,17'd38260,17'd39261,17'd36820,17'd36814,17'd36515,17'd37634,17'd37367,17'd36815,17'd36515,17'd36820,17'd38957,17'd36385,17'd36385,17'd35971,17'd39262,17'd39117,17'd39263,17'd39264,17'd39265,17'd39266,17'd39267,17'd39268,17'd39269,17'd39124,17'd39125,17'd39270,17'd38658,17'd39271,17'd37244,17'd37899,17'd38660,17'd39272,17'd39273,17'd39128,17'd39129,17'd39274,17'd37905,17'd37904,17'd39275,17'd39276,17'd39277,17'd26902,17'd28853,17'd26064,17'd28369,17'd30432,17'd30431,17'd39278,17'd23038,17'd22330,17'd22680,17'd22329,17'd39278,17'd29376,17'd31502,17'd23736,17'd30579,17'd32351,17'd37117,17'd29242,17'd23561,17'd25567,17'd27515,17'd27372,17'd30586,17'd26782,17'd26781,17'd31353,17'd36541,17'd38666,17'd38405,17'd28728,17'd28857,17'd29248,17'd32017,17'd33485,17'd33165,17'd28982,17'd32017,17'd38537,17'd26064,17'd31033,17'd39279,17'd38976,17'd39280,17'd39281,17'd39282,17'd24592,17'd24089,17'd34284,17'd29101,17'd33318,17'd25180,17'd24744,17'd24897,17'd25438,17'd25317,17'd28597,17'd33000,17'd33484,17'd39283,17'd26530,17'd28486,17'd31503,17'd27885,17'd37514,17'd39284,17'd39285,17'd38982,17'd38983,17'd39286,17'd35167,17'd34633,17'd39136,17'd38986,17'd37265,17'd38546,17'd28013,17'd26905,17'd39287,17'd31046,17'd25439,17'd30879,17'd24590,17'd24744,17'd30903,17'd32848,17'd38992,17'd27517,17'd39288,17'd39289,17'd39290,17'd39291,17'd33671,17'd39292,17'd39293,17'd39294,17'd39295,17'd39296,17'd39147,17'd39297,17'd33352,17'd39298,17'd39299,17'd36294,17'd39300,17'd39301,17'd19695,17'd39302,17'd39153,17'd39303,17'd37686,17'd39304,17'd39305,17'd39306,17'd39159,17'd39307,17'd38700,17'd39308,17'd39309,17'd39310,17'd39311,17'd22250,17'd38439,17'd39312,17'd34922,17'd31551,17'd29593,17'd29593,17'd10515,17'd10642,17'd30933,17'd29592,17'd6219,17'd27935,17'd25627,17'd5004,17'd28536,17'd4842,17'd5336,17'd30638,17'd5163,17'd4847,17'd33533,17'd39313,17'd5756,17'd27570,17'd6554,17'd9091,17'd34334,17'd39314,17'd4196,17'd39315,17'd39316,17'd39317,17'd38706,17'd39318,17'd39021,17'd39319,17'd39172,17'd39320,17'd39321,17'd39322,17'd39323,17'd39026,17'd2368,17'd2546,17'd39324,17'd39325,17'd39176,17'd39177,17'd7026,17'd39326,17'd39179,17'd39180,17'd10906,17'd39032,17'd11867,17'd38202,17'd39327,17'd39328,17'd6418,17'd7364,17'd9124,17'd7538,17'd7538,17'd9124,17'd33051,17'd33051,17'd31562,17'd28066,17'd33050,17'd6721,17'd1946,17'd5371,17'd1261,17'd1261,17'd446,17'd623,17'd447,17'd800,17'd38863,17'd29753,17'd39329,17'd39330
},
'{
17'd6420,17'd4245,17'd4245,17'd6420,17'd6420,17'd4245,17'd6420,17'd25384,17'd6420,17'd4245,17'd3101,17'd14188,17'd27714,17'd1127,17'd17,17'd3905,17'd3905,17'd3905,17'd1278,17'd980,17'd7385,17'd7385,17'd7225,17'd6437,17'd5804,17'd4250,17'd4580,17'd2431,17'd1704,17'd1841,17'd35772,17'd1425,17'd1561,17'd3266,17'd1709,17'd1290,17'd2619,17'd14875,17'd39331,17'd5068,17'd20017,17'd36326,17'd39040,17'd39185,17'd38872,17'd39042,17'd17811,17'd16033,17'd16519,17'd17206,17'd18655,17'd17204,17'd39332,17'd38591,17'd38591,17'd36611,17'd39333,17'd39334,17'd39335,17'd39336,17'd39191,17'd39337,17'd39338,17'd39339,17'd39340,17'd39341,17'd38881,17'd39342,17'd39343,17'd38473,17'd39344,17'd39195,17'd39345,17'd17213,17'd14782,17'd13104,17'd14109,17'd29182,17'd38477,17'd39346,17'd39347,17'd39348,17'd39349,17'd38739,17'd38349,17'd38890,17'd39057,17'd6645,17'd39058,17'd38891,17'd37971,17'd37837,17'd37838,17'd6949,17'd39350,17'd39351,17'd39062,17'd39352,17'd39353,17'd39354,17'd39355,17'd39356,17'd39357,17'd7456,17'd10860,17'd17352,17'd10028,17'd8578,17'd19923,17'd12867,17'd17481,17'd8571,17'd8725,17'd9041,17'd14811,17'd26498,17'd38904,17'd31760,17'd9887,17'd8409,17'd23679,17'd27487,17'd24029,17'd27985,17'd39358,17'd39210,17'd32919,17'd31941,17'd34381,17'd34381,17'd30834,17'd31587,17'd28344,17'd26371,17'd24858,17'd22816,17'd19281,17'd10328,17'd10329,17'd11670,17'd11671,17'd10024,17'd9885,17'd10992,17'd9741,17'd11809,17'd10174,17'd9039,17'd15297,17'd21507,17'd8885,17'd17480,17'd24361,17'd10174,17'd13887,17'd15569,17'd15048,17'd11277,17'd10329,17'd28352,17'd22817,17'd21505,17'd26758,17'd27485,17'd30078,17'd39359,17'd39212,17'd38908,17'd38364,17'd38751,17'd17476,17'd39360,17'd32447,17'd31603,17'd33578,17'd33246,17'd33244,17'd39361,17'd39362,17'd9613,17'd39363,17'd39364,17'd39365,17'd39366,17'd39367,17'd39368,17'd31625,17'd31797,17'd39369,17'd39370,17'd39371,17'd39372,17'd39373,17'd39374,17'd39375,17'd39376,17'd39377,17'd39378,17'd39379,17'd39380,17'd39381,17'd39382,17'd39383,17'd39384,17'd39385,17'd39386,17'd39387,17'd39388,17'd39389,17'd39390,17'd39391,17'd39392,17'd39393,17'd39394,17'd39395,17'd39395,17'd39396,17'd39397,17'd39398,17'd39399,17'd39400,17'd39401,17'd39402,17'd39403,17'd39404,17'd39405,17'd39406,17'd39407,17'd39408,17'd39409,17'd39410,17'd39411,17'd33915,17'd38133,17'd39412,17'd39413,17'd39414,17'd36964,17'd37226,17'd36820,17'd39415,17'd39416,17'd36819,17'd37097,17'd39417,17'd38957,17'd36385,17'd36385,17'd36385,17'd38133,17'd39418,17'd39419,17'd39420,17'd39421,17'd39422,17'd39423,17'd39424,17'd39425,17'd39426,17'd39427,17'd39428,17'd38968,17'd39429,17'd39430,17'd37899,17'd38660,17'd39431,17'd39432,17'd39433,17'd39434,17'd39435,17'd37905,17'd37904,17'd39275,17'd39436,17'd32184,17'd26902,17'd26902,17'd26062,17'd25567,17'd29244,17'd30431,17'd39278,17'd22859,17'd22330,17'd32827,17'd30277,17'd39278,17'd29376,17'd23918,17'd29099,17'd30579,17'd32008,17'd29828,17'd34137,17'd24417,17'd27765,17'd27515,17'd27146,17'd30586,17'd26782,17'd26901,17'd39437,17'd39438,17'd39439,17'd38405,17'd28728,17'd28857,17'd29248,17'd32017,17'd28373,17'd32505,17'd36989,17'd28373,17'd28726,17'd28720,17'd23565,17'd31191,17'd39278,17'd39440,17'd39441,17'd39442,17'd34452,17'd25439,17'd27763,17'd28850,17'd39443,17'd29976,17'd24898,17'd24897,17'd25438,17'd28369,17'd28597,17'd28597,17'd33484,17'd39444,17'd26530,17'd28486,17'd27642,17'd27885,17'd37514,17'd38813,17'd38981,17'd39445,17'd38160,17'd39286,17'd35167,17'd34769,17'd34633,17'd38029,17'd37265,17'd38546,17'd36283,17'd38032,17'd39446,17'd37123,17'd25439,17'd29100,17'd26657,17'd24589,17'd25568,17'd33510,17'd39447,17'd39448,17'd39289,17'd39290,17'd39290,17'd37251,17'd39449,17'd38812,17'd39450,17'd33820,17'd39451,17'd39452,17'd39453,17'd39454,17'd39455,17'd39456,17'd39457,17'd38833,17'd39458,17'd39459,17'd19691,17'd39460,17'd20979,17'd38562,17'd39461,17'd39462,17'd39463,17'd39464,17'd39465,17'd39466,17'd38566,17'd39308,17'd39309,17'd39011,17'd22250,17'd22250,17'd38439,17'd39467,17'd35196,17'd31551,17'd29593,17'd29593,17'd10515,17'd10515,17'd31243,17'd29592,17'd6220,17'd5614,17'd25627,17'd5002,17'd5327,17'd5327,17'd5335,17'd30638,17'd5163,17'd4846,17'd39468,17'd39469,17'd4837,17'd4687,17'd31717,17'd9091,17'd34334,17'd39470,17'd4193,17'd39471,17'd39472,17'd39473,17'd38850,17'd39474,17'd39475,17'd39476,17'd39023,17'd39320,17'd39477,17'd39478,17'd39479,17'd39480,17'd2368,17'd2546,17'd39324,17'd39325,17'd39176,17'd39481,17'd7026,17'd39326,17'd39179,17'd39180,17'd10790,17'd39482,17'd39483,17'd38859,17'd39484,17'd38861,17'd15484,17'd7364,17'd7538,17'd7538,17'd7538,17'd9124,17'd33051,17'd33051,17'd31562,17'd28066,17'd33050,17'd5631,17'd5940,17'd5371,17'd1261,17'd1261,17'd446,17'd623,17'd447,17'd1540,17'd27948,17'd787,17'd16264,17'd16006
},
'{
17'd6420,17'd4245,17'd4245,17'd6420,17'd6420,17'd4245,17'd6420,17'd25384,17'd6420,17'd4245,17'd3101,17'd14188,17'd10535,17'd466,17'd18,17'd3905,17'd3905,17'd3905,17'd1278,17'd980,17'd7385,17'd7385,17'd6745,17'd5971,17'd5804,17'd4250,17'd2605,17'd2431,17'd1704,17'd1705,17'd1707,17'd3108,17'd3439,17'd3266,17'd1710,17'd1290,17'd39485,17'd14875,17'd14197,17'd5068,17'd20017,17'd39486,17'd39487,17'd39185,17'd39488,17'd17574,17'd16768,17'd16034,17'd17319,17'd17206,17'd18655,17'd17204,17'd33859,17'd39489,17'd39490,17'd38211,17'd38593,17'd39491,17'd39492,17'd39493,17'd39494,17'd39495,17'd39495,17'd39496,17'd39497,17'd39498,17'd38881,17'd39499,17'd37456,17'd36467,17'd39500,17'd39501,17'd35216,17'd17213,17'd14782,17'd13104,17'd9164,17'd29182,17'd38477,17'd39346,17'd39502,17'd6782,17'd39349,17'd39503,17'd38891,17'd38891,17'd39504,17'd39057,17'd39505,17'd38891,17'd37971,17'd38484,17'd38604,17'd6949,17'd39350,17'd39351,17'd39062,17'd39506,17'd39507,17'd39508,17'd39509,17'd39510,17'd39511,17'd18567,17'd15441,17'd17850,17'd8580,17'd23343,17'd21208,17'd12867,17'd25147,17'd8571,17'd8725,17'd9040,17'd17123,17'd17848,17'd38904,17'd26260,17'd9483,17'd10607,17'd9340,17'd19281,17'd18327,17'd24208,17'd34542,17'd30832,17'd31439,17'd34381,17'd34381,17'd34381,17'd30676,17'd31587,17'd28344,17'd24537,17'd14258,17'd29789,17'd19281,17'd10328,17'd10330,17'd11670,17'd10329,17'd17719,17'd9741,17'd9885,17'd9884,17'd9741,17'd9346,17'd9038,17'd15297,17'd21507,17'd9045,17'd14811,17'd17716,17'd10173,17'd9345,17'd24037,17'd9618,17'd9739,17'd10330,17'd11669,17'd18327,17'd19408,17'd26758,17'd27485,17'd30078,17'd38751,17'd37611,17'd39359,17'd38750,17'd39512,17'd39513,17'd30840,17'd32608,17'd31603,17'd30088,17'd39514,17'd38370,17'd39515,17'd39516,17'd10021,17'd39517,17'd39518,17'd39519,17'd39520,17'd39521,17'd39522,17'd31625,17'd39523,17'd39524,17'd39525,17'd39526,17'd33268,17'd39527,17'd39528,17'd39529,17'd39530,17'd39531,17'd39532,17'd39533,17'd39534,17'd39535,17'd39536,17'd39537,17'd39538,17'd39107,17'd39539,17'd39388,17'd39540,17'd39541,17'd39542,17'd39543,17'd39544,17'd39545,17'd39546,17'd39547,17'd39548,17'd39549,17'd39550,17'd39551,17'd39552,17'd39553,17'd39554,17'd39555,17'd39556,17'd39557,17'd39558,17'd39559,17'd39560,17'd39561,17'd39562,17'd39563,17'd39564,17'd39565,17'd39566,17'd35137,17'd39567,17'd38130,17'd36818,17'd36810,17'd36243,17'd39568,17'd36669,17'd39569,17'd39569,17'd36964,17'd38957,17'd36385,17'd36385,17'd36385,17'd38009,17'd39570,17'd39571,17'd39572,17'd39573,17'd39574,17'd39575,17'd38795,17'd39576,17'd39426,17'd39427,17'd39577,17'd39578,17'd39579,17'd38020,17'd37899,17'd38660,17'd39580,17'd39581,17'd39582,17'd39583,17'd39435,17'd38973,17'd37904,17'd39584,17'd39585,17'd32495,17'd26902,17'd27258,17'd28602,17'd25567,17'd29103,17'd23916,17'd29973,17'd35018,17'd22330,17'd22330,17'd22328,17'd29973,17'd29376,17'd29099,17'd23736,17'd30579,17'd23569,17'd30128,17'd34137,17'd24744,17'd27638,17'd26903,17'd27372,17'd30586,17'd26782,17'd26901,17'd39437,17'd39438,17'd39439,17'd39586,17'd28728,17'd28857,17'd29248,17'd32017,17'd28373,17'd33165,17'd37250,17'd28373,17'd26901,17'd28130,17'd23386,17'd39587,17'd29973,17'd39588,17'd31834,17'd39589,17'd39590,17'd30883,17'd27763,17'd25438,17'd39591,17'd25320,17'd25029,17'd28596,17'd25177,17'd28369,17'd28597,17'd28597,17'd33484,17'd31856,17'd26530,17'd26901,17'd27642,17'd30279,17'd37514,17'd39284,17'd39285,17'd38982,17'd38983,17'd39286,17'd38284,17'd34769,17'd34633,17'd39592,17'd39593,17'd38546,17'd39594,17'd39595,17'd26066,17'd39596,17'd36565,17'd29100,17'd26283,17'd23728,17'd28719,17'd39597,17'd27028,17'd35734,17'd34480,17'd34480,17'd36869,17'd29535,17'd38538,17'd39591,17'd34883,17'd31836,17'd39598,17'd39599,17'd39600,17'd39601,17'd39602,17'd39603,17'd39604,17'd38426,17'd39605,17'd39606,17'd39607,17'd20658,17'd22727,17'd39608,17'd39609,17'd35331,17'd39610,17'd38312,17'd38436,17'd39307,17'd38437,17'd39308,17'd20250,17'd39011,17'd22250,17'd22250,17'd38439,17'd39467,17'd35196,17'd31551,17'd39611,17'd29593,17'd10515,17'd27815,17'd29592,17'd29592,17'd6391,17'd5919,17'd25627,17'd5002,17'd5153,17'd4996,17'd5334,17'd5335,17'd5161,17'd4529,17'd4515,17'd39469,17'd4523,17'd32552,17'd30638,17'd6390,17'd34334,17'd39612,17'd39613,17'd39614,17'd39615,17'd39616,17'd39617,17'd39618,17'd39619,17'd39476,17'd39620,17'd39621,17'd39622,17'd39623,17'd39624,17'd39625,17'd2363,17'd2546,17'd36746,17'd39626,17'd39176,17'd39481,17'd7026,17'd5353,17'd3872,17'd39180,17'd10790,17'd39032,17'd38458,17'd38202,17'd37958,17'd38459,17'd6417,17'd7364,17'd7538,17'd7538,17'd7538,17'd9124,17'd38460,17'd33051,17'd31562,17'd28066,17'd11882,17'd4559,17'd6415,17'd4880,17'd1261,17'd1261,17'd446,17'd623,17'd447,17'd1540,17'd39627,17'd1116,17'd39628,17'd39629
},
'{
17'd6420,17'd4245,17'd6420,17'd6420,17'd6420,17'd4245,17'd6420,17'd25384,17'd4245,17'd4733,17'd3101,17'd14188,17'd10535,17'd1127,17'd16,17'd3905,17'd3905,17'd3905,17'd1278,17'd27,17'd7385,17'd7061,17'd6437,17'd5971,17'd5656,17'd4250,17'd2605,17'd1422,17'd39630,17'd1705,17'd3599,17'd1425,17'd1979,17'd1146,17'd1710,17'd1148,17'd39631,17'd39632,17'd15369,17'd5068,17'd29045,17'd39633,17'd39487,17'd39634,17'd34673,17'd17574,17'd16987,17'd17445,17'd19255,17'd17206,17'd18774,17'd19621,17'd39635,17'd19136,17'd36330,17'd18301,17'd38877,17'd39636,17'd39190,17'd39637,17'd39638,17'd39639,17'd39640,17'd39641,17'd39497,17'd39642,17'd39643,17'd39499,17'd37456,17'd36332,17'd39644,17'd38601,17'd34191,17'd39645,17'd17105,17'd14109,17'd9015,17'd29182,17'd38477,17'd25260,17'd39646,17'd39647,17'd6483,17'd39648,17'd38891,17'd38891,17'd39504,17'd6645,17'd39649,17'd39503,17'd37971,17'd37320,17'd37838,17'd39650,17'd39651,17'd39652,17'd39653,17'd39654,17'd39655,17'd39656,17'd39657,17'd39658,17'd39659,17'd18567,17'd15441,17'd15056,17'd11674,17'd8579,17'd8248,17'd18919,17'd25147,17'd8731,17'd8724,17'd9045,17'd14811,17'd39660,17'd26259,17'd24712,17'd9483,17'd8567,17'd10992,17'd28352,17'd23513,17'd26149,17'd34542,17'd30832,17'd31439,17'd34381,17'd34381,17'd34381,17'd30676,17'd30072,17'd28943,17'd24857,17'd25143,17'd29789,17'd19281,17'd10328,17'd10330,17'd12863,17'd10330,17'd26152,17'd9884,17'd9741,17'd9884,17'd9885,17'd9346,17'd8874,17'd9045,17'd16066,17'd9042,17'd14811,17'd14674,17'd15807,17'd15187,17'd9619,17'd17839,17'd11134,17'd11670,17'd28463,17'd23513,17'd19408,17'd26758,17'd29784,17'd39661,17'd38751,17'd37611,17'd28349,17'd38750,17'd38366,17'd17349,17'd39662,17'd37071,17'd31778,17'd39514,17'd37741,17'd39663,17'd39664,17'd39665,17'd39666,17'd39667,17'd39668,17'd39669,17'd39670,17'd39671,17'd36362,17'd31797,17'd39672,17'd39673,17'd39674,17'd39675,17'd39676,17'd39677,17'd39678,17'd39679,17'd39680,17'd39681,17'd39682,17'd39683,17'd39684,17'd39685,17'd39686,17'd39687,17'd39688,17'd39689,17'd39690,17'd39691,17'd39692,17'd39693,17'd39694,17'd39695,17'd39696,17'd39697,17'd39698,17'd39699,17'd39700,17'd39701,17'd39702,17'd39703,17'd39704,17'd39705,17'd39706,17'd39707,17'd39708,17'd39709,17'd39710,17'd39711,17'd39712,17'd39713,17'd39714,17'd39715,17'd39716,17'd39717,17'd39718,17'd39719,17'd33915,17'd35273,17'd37097,17'd36668,17'd36820,17'd39720,17'd38391,17'd36812,17'd36812,17'd36964,17'd38788,17'd36384,17'd36385,17'd35972,17'd38389,17'd39721,17'd39722,17'd39723,17'd39724,17'd39725,17'd39726,17'd39727,17'd39728,17'd39729,17'd39730,17'd39731,17'd39732,17'd39733,17'd39734,17'd38020,17'd38660,17'd39735,17'd39736,17'd39737,17'd39738,17'd39739,17'd38973,17'd37904,17'd39584,17'd39740,17'd39741,17'd26902,17'd27258,17'd27766,17'd25567,17'd29103,17'd23916,17'd23216,17'd39742,17'd22330,17'd36986,17'd22501,17'd23216,17'd29376,17'd23565,17'd31502,17'd29530,17'd23388,17'd23923,17'd23384,17'd24895,17'd28720,17'd28725,17'd34637,17'd30586,17'd26782,17'd26781,17'd31353,17'd39743,17'd38404,17'd39586,17'd28728,17'd28857,17'd29248,17'd32017,17'd28373,17'd33165,17'd32505,17'd33485,17'd28486,17'd25317,17'd36987,17'd39742,17'd23389,17'd39744,17'd39745,17'd39746,17'd39747,17'd39293,17'd24417,17'd25568,17'd39591,17'd25438,17'd28719,17'd27764,17'd28717,17'd25567,17'd28597,17'd28597,17'd25568,17'd31520,17'd28482,17'd26901,17'd27642,17'd30279,17'd38813,17'd38813,17'd38981,17'd39748,17'd38160,17'd38983,17'd38284,17'd39749,17'd36548,17'd39592,17'd38987,17'd30000,17'd39750,17'd39751,17'd39752,17'd36550,17'd36565,17'd24090,17'd26283,17'd23728,17'd27764,17'd25567,17'd39753,17'd34479,17'd39754,17'd34128,17'd27027,17'd28853,17'd25829,17'd26172,17'd28368,17'd36152,17'd39755,17'd39756,17'd39757,17'd39758,17'd39759,17'd39760,17'd39761,17'd39762,17'd39763,17'd39764,17'd39765,17'd39766,17'd27811,17'd21124,17'd39767,17'd5908,17'd36022,17'd39768,17'd39769,17'd39466,17'd38313,17'd39770,17'd19479,17'd22422,17'd22250,17'd22088,17'd38056,17'd39771,17'd39772,17'd31551,17'd39611,17'd29593,17'd10515,17'd27815,17'd29593,17'd29592,17'd6391,17'd6221,17'd25627,17'd5005,17'd38442,17'd33532,17'd5329,17'd5335,17'd5161,17'd34656,17'd4358,17'd39773,17'd5477,17'd4840,17'd31553,17'd6554,17'd34334,17'd39774,17'd39775,17'd39776,17'd39777,17'd39778,17'd39779,17'd39780,17'd39781,17'd39476,17'd39782,17'd39783,17'd39784,17'd39785,17'd39786,17'd39625,17'd39787,17'd2546,17'd36746,17'd36453,17'd35058,17'd39481,17'd6236,17'd39788,17'd3871,17'd39789,17'd10790,17'd10790,17'd39790,17'd38859,17'd38860,17'd38581,17'd39791,17'd7364,17'd7538,17'd7538,17'd7538,17'd9124,17'd38460,17'd38460,17'd38719,17'd28066,17'd11882,17'd5183,17'd5630,17'd4880,17'd1261,17'd1261,17'd446,17'd623,17'd447,17'd1540,17'd22264,17'd433,17'd29442,17'd16634
},
'{
17'd6420,17'd4245,17'd6420,17'd25384,17'd6420,17'd4245,17'd6420,17'd25384,17'd4245,17'd4246,17'd3252,17'd27714,17'd17917,17'd2,17'd18,17'd3905,17'd4089,17'd3905,17'd1278,17'd27,17'd7061,17'd7061,17'd6437,17'd5971,17'd5656,17'd4250,17'd2947,17'd1422,17'd39630,17'd1705,17'd3599,17'd3108,17'd3266,17'd1146,17'd835,17'd38867,17'd32256,17'd39792,17'd3767,17'd39793,17'd25508,17'd39794,17'd39795,17'd39634,17'd34673,17'd39796,17'd17810,17'd17320,17'd19255,17'd27461,17'd17689,17'd39797,17'd39798,17'd19016,17'd18780,17'd38593,17'd39799,17'd39492,17'd39800,17'd39801,17'd39802,17'd39803,17'd39804,17'd39805,17'd39806,17'd39642,17'd39643,17'd39807,17'd38089,17'd39808,17'd39644,17'd37459,17'd32268,17'd39809,17'd16779,17'd9707,17'd9164,17'd39810,17'd39811,17'd24978,17'd39812,17'd39647,17'd6483,17'd39813,17'd39503,17'd38891,17'd39814,17'd39815,17'd39816,17'd39503,17'd38351,17'd37839,17'd38892,17'd39650,17'd39651,17'd39817,17'd39818,17'd39819,17'd39820,17'd39656,17'd39821,17'd39822,17'd7134,17'd39823,17'd18920,17'd17016,17'd11674,17'd8579,17'd8248,17'd18919,17'd21987,17'd8731,17'd8724,17'd9348,17'd17123,17'd28353,17'd26259,17'd30217,17'd9483,17'd8877,17'd9741,17'd28463,17'd24706,17'd26371,17'd39824,17'd37065,17'd30834,17'd34381,17'd34381,17'd30221,17'd31440,17'd29645,17'd28816,17'd23512,17'd18681,17'd14381,17'd27623,17'd19281,17'd19280,17'd11400,17'd11526,17'd10329,17'd9883,17'd9740,17'd9884,17'd9885,17'd9346,17'd9039,17'd9040,17'd8882,17'd9194,17'd14811,17'd14674,17'd9479,17'd17011,17'd15048,17'd17839,17'd10479,17'd11133,17'd21206,17'd14264,17'd19408,17'd27486,17'd37856,17'd39825,17'd39826,17'd39826,17'd38366,17'd38366,17'd38910,17'd39827,17'd32446,17'd38109,17'd33250,17'd39514,17'd33244,17'd39828,17'd39829,17'd39830,17'd39831,17'd39832,17'd39833,17'd39834,17'd39835,17'd39836,17'd39837,17'd39838,17'd39839,17'd39840,17'd39841,17'd39842,17'd39843,17'd39844,17'd39845,17'd39846,17'd39847,17'd39848,17'd39849,17'd39850,17'd39851,17'd39852,17'd39853,17'd39854,17'd39855,17'd39856,17'd39857,17'd39858,17'd39859,17'd39860,17'd39861,17'd39862,17'd39863,17'd39864,17'd39865,17'd39866,17'd39867,17'd39868,17'd39869,17'd39870,17'd39871,17'd39872,17'd39873,17'd39874,17'd39875,17'd39876,17'd39877,17'd39709,17'd39878,17'd39879,17'd39880,17'd39881,17'd39882,17'd39883,17'd39884,17'd39091,17'd39885,17'd39886,17'd34858,17'd35839,17'd39261,17'd39720,17'd36244,17'd39116,17'd36812,17'd36660,17'd39417,17'd36244,17'd36384,17'd36385,17'd39887,17'd39888,17'd39889,17'd39890,17'd39891,17'd39892,17'd39893,17'd38964,17'd39894,17'd39895,17'd39896,17'd39897,17'd38660,17'd39898,17'd39126,17'd37900,17'd39899,17'd39900,17'd39901,17'd39902,17'd39903,17'd39904,17'd37904,17'd39905,17'd39906,17'd39907,17'd39741,17'd28853,17'd27146,17'd25708,17'd25567,17'd29103,17'd23916,17'd37386,17'd39908,17'd36986,17'd22329,17'd33158,17'd23217,17'd29099,17'd23918,17'd31502,17'd23387,17'd23388,17'd23387,17'd23564,17'd25030,17'd28720,17'd28725,17'd33163,17'd30586,17'd27371,17'd26902,17'd37908,17'd35854,17'd39909,17'd39586,17'd32018,17'd29249,17'd29248,17'd32017,17'd28373,17'd33485,17'd32505,17'd39910,17'd30586,17'd27511,17'd33651,17'd39911,17'd22329,17'd39912,17'd31658,17'd39913,17'd34638,17'd39914,17'd28851,17'd28719,17'd29970,17'd28369,17'd27512,17'd27764,17'd25709,17'd25567,17'd28597,17'd28597,17'd25568,17'd33484,17'd28482,17'd26901,17'd27642,17'd30279,17'd33319,17'd29977,17'd27643,17'd27769,17'd38982,17'd38160,17'd35725,17'd39749,17'd38984,17'd34633,17'd38986,17'd30000,17'd32849,17'd39915,17'd26532,17'd36409,17'd39916,17'd24415,17'd39917,17'd39918,17'd28596,17'd28597,17'd25833,17'd27146,17'd31035,17'd28486,17'd27027,17'd28853,17'd25829,17'd26060,17'd29533,17'd34895,17'd39919,17'd39920,17'd39921,17'd39922,17'd39923,17'd39924,17'd39925,17'd39926,17'd39927,17'd39928,17'd39929,17'd39930,17'd39931,17'd21441,17'd39932,17'd36729,17'd4829,17'd39933,17'd39769,17'd38437,17'd39934,17'd39935,17'd19479,17'd22422,17'd22088,17'd22088,17'd38056,17'd37286,17'd35051,17'd29158,17'd29593,17'd29592,17'd10515,17'd27815,17'd29593,17'd27815,17'd7668,17'd6221,17'd5004,17'd4686,17'd4188,17'd38441,17'd4845,17'd5160,17'd5162,17'd4529,17'd4833,17'd39936,17'd4186,17'd4682,17'd37029,17'd37030,17'd39937,17'd39938,17'd39939,17'd39777,17'd39940,17'd39941,17'd39942,17'd39943,17'd39781,17'd39476,17'd39782,17'd39944,17'd39945,17'd39946,17'd22775,17'd39625,17'd39787,17'd2546,17'd36746,17'd36453,17'd35058,17'd39481,17'd6236,17'd39788,17'd3871,17'd39947,17'd10790,17'd10906,17'd11048,17'd39948,17'd39327,17'd4867,17'd6258,17'd7364,17'd7538,17'd7538,17'd7538,17'd9124,17'd38460,17'd33051,17'd31899,17'd28066,17'd11882,17'd4559,17'd6415,17'd4880,17'd1261,17'd1680,17'd2249,17'd627,17'd3100,17'd39949,17'd431,17'd251,17'd649,17'd39950
},
'{
17'd6420,17'd6420,17'd6420,17'd25384,17'd6420,17'd4245,17'd4245,17'd6420,17'd4245,17'd4733,17'd2935,17'd14070,17'd10535,17'd14,17'd16,17'd3905,17'd4089,17'd4089,17'd1278,17'd27,17'd7061,17'd7061,17'd6437,17'd5971,17'd5656,17'd4251,17'd2947,17'd1422,17'd39630,17'd1285,17'd1560,17'd2949,17'd1428,17'd998,17'd1290,17'd38867,17'd32256,17'd15749,17'd3767,17'd39951,17'd25254,17'd39794,17'd39795,17'd39634,17'd34673,17'd39796,17'd17810,17'd19008,17'd25512,17'd27461,17'd17689,17'd20150,17'd20025,17'd18417,17'd39952,17'd39953,17'd39954,17'd39955,17'd39048,17'd39956,17'd39957,17'd39958,17'd39959,17'd39960,17'd39961,17'd39962,17'd39050,17'd37717,17'd39963,17'd39808,17'd39644,17'd37319,17'd39964,17'd14639,17'd13104,17'd9164,17'd29182,17'd38477,17'd39965,17'd25913,17'd39812,17'd6640,17'd39966,17'd39813,17'd39503,17'd38891,17'd39814,17'd39200,17'd39967,17'd39968,17'd38093,17'd6947,17'd38606,17'd6950,17'd39969,17'd39970,17'd39971,17'd39819,17'd39820,17'd39972,17'd39973,17'd39974,17'd39975,17'd25415,17'd18920,17'd17016,17'd17240,17'd8579,17'd8248,17'd10339,17'd35514,17'd8729,17'd8878,17'd9045,17'd16795,17'd17123,17'd8878,17'd39976,17'd12586,17'd24999,17'd12116,17'd11275,17'd21363,17'd29065,17'd37733,17'd37065,17'd30834,17'd34835,17'd30677,17'd30221,17'd31587,17'd35372,17'd29778,17'd24705,17'd24994,17'd14381,17'd28352,17'd19281,17'd19280,17'd11400,17'd11526,17'd10329,17'd9883,17'd9739,17'd9884,17'd9885,17'd9346,17'd10174,17'd9194,17'd8883,17'd10175,17'd39977,17'd10334,17'd9479,17'd17011,17'd15048,17'd17839,17'd10479,17'd11132,17'd11275,17'd16325,17'd21671,17'd27486,17'd37856,17'd38366,17'd39978,17'd39978,17'd38366,17'd38366,17'd38910,17'd39979,17'd39980,17'd38109,17'd30088,17'd16434,17'd18446,17'd39361,17'd39664,17'd39665,17'd39981,17'd39982,17'd39983,17'd39984,17'd39835,17'd39985,17'd39837,17'd39986,17'd39987,17'd39988,17'd39989,17'd39842,17'd33750,17'd39990,17'd39991,17'd39992,17'd39993,17'd39994,17'd39995,17'd39996,17'd39997,17'd39998,17'd39248,17'd39999,17'd39553,17'd40000,17'd40001,17'd40002,17'd40003,17'd40004,17'd40005,17'd39865,17'd40006,17'd40007,17'd40008,17'd40009,17'd40010,17'd40011,17'd40012,17'd40013,17'd40014,17'd40015,17'd40016,17'd40017,17'd40018,17'd40019,17'd40020,17'd40021,17'd40022,17'd40023,17'd40024,17'd40025,17'd40026,17'd40027,17'd40028,17'd40029,17'd40030,17'd40031,17'd40032,17'd40033,17'd40034,17'd38958,17'd36384,17'd36512,17'd36813,17'd37097,17'd40035,17'd38391,17'd36244,17'd36384,17'd39262,17'd40036,17'd40037,17'd40038,17'd40039,17'd40040,17'd40041,17'd40042,17'd40043,17'd39576,17'd40044,17'd40045,17'd39899,17'd39577,17'd39732,17'd37900,17'd39899,17'd40046,17'd40047,17'd40048,17'd39903,17'd39904,17'd37904,17'd39905,17'd39906,17'd39907,17'd33308,17'd28853,17'd27146,17'd25565,17'd25567,17'd29103,17'd32659,17'd29828,17'd40049,17'd36986,17'd22329,17'd33158,17'd29828,17'd23733,17'd23732,17'd23918,17'd23386,17'd29686,17'd23386,17'd28849,17'd25180,17'd28720,17'd27259,17'd30586,17'd27027,17'd27259,17'd26902,17'd38025,17'd35425,17'd39909,17'd40050,17'd33486,17'd29249,17'd29248,17'd32017,17'd28373,17'd33485,17'd32505,17'd40051,17'd27146,17'd25320,17'd32680,17'd40052,17'd22328,17'd40053,17'd31192,17'd40054,17'd40055,17'd40056,17'd29688,17'd27764,17'd25435,17'd27765,17'd33484,17'd33803,17'd28597,17'd25567,17'd28599,17'd33000,17'd25568,17'd33484,17'd28482,17'd26901,17'd27642,17'd30279,17'd33319,17'd33001,17'd40057,17'd27769,17'd38982,17'd38982,17'd36001,17'd40058,17'd40059,17'd29695,17'd38986,17'd40060,17'd27771,17'd40061,17'd40062,17'd40063,17'd40064,17'd24088,17'd34884,17'd28718,17'd28974,17'd25709,17'd25708,17'd27146,17'd31035,17'd28727,17'd28486,17'd26902,17'd25703,17'd23554,17'd29103,17'd23921,17'd35455,17'd40065,17'd39921,17'd40066,17'd40067,17'd40068,17'd30310,17'd40069,17'd40070,17'd40071,17'd40072,17'd40073,17'd21128,17'd28415,17'd39303,17'd40074,17'd4669,17'd40075,17'd40076,17'd38700,17'd39934,17'd40077,17'd19087,17'd18619,17'd18131,17'd18131,17'd38056,17'd40078,17'd37151,17'd29158,17'd29593,17'd29592,17'd10642,17'd27815,17'd29593,17'd27815,17'd7668,17'd6391,17'd31553,17'd4686,17'd5477,17'd40079,17'd4687,17'd5329,17'd5157,17'd4529,17'd4833,17'd40080,17'd40081,17'd6067,17'd4685,17'd5163,17'd40082,17'd40083,17'd40084,17'd40085,17'd40086,17'd40087,17'd40088,17'd40089,17'd3685,17'd40090,17'd40091,17'd40092,17'd40093,17'd40094,17'd40095,17'd39625,17'd39787,17'd40096,17'd40097,17'd36453,17'd2737,17'd40098,17'd6082,17'd3567,17'd40099,17'd40100,17'd39789,17'd10388,17'd39181,17'd40101,17'd39484,17'd38581,17'd39791,17'd7364,17'd7538,17'd7538,17'd7538,17'd38460,17'd38460,17'd38460,17'd34002,17'd28066,17'd11882,17'd5183,17'd5630,17'd4880,17'd1261,17'd1261,17'd625,17'd623,17'd233,17'd39949,17'd611,17'd40102,17'd1543,17'd648
},
'{
17'd4428,17'd4088,17'd6420,17'd6420,17'd6420,17'd4245,17'd6420,17'd25384,17'd4245,17'd4246,17'd3252,17'd27714,17'd17917,17'd466,17'd18,17'd3905,17'd3905,17'd3905,17'd27,17'd980,17'd7728,17'd7060,17'd6903,17'd5971,17'd5379,17'd4739,17'd2431,17'd38865,17'd37171,17'd1705,17'd3599,17'd1561,17'd1146,17'd998,17'd23659,17'd40103,17'd22970,17'd14753,17'd3929,17'd39951,17'd18766,17'd35912,17'd40104,17'd40105,17'd40106,17'd18175,17'd19257,17'd19255,17'd19007,17'd18655,17'd17941,17'd19622,17'd20295,17'd18537,17'd39333,17'd40107,17'd40108,17'd39190,17'd40109,17'd40110,17'd40111,17'd40112,17'd40113,17'd39960,17'd40114,17'd39642,17'd38087,17'd37718,17'd40115,17'd40116,17'd39195,17'd37721,17'd39645,17'd16665,17'd9707,17'd9581,17'd9014,17'd39197,17'd40117,17'd40118,17'd6939,17'd6640,17'd39966,17'd40119,17'd39816,17'd39813,17'd6485,17'd39505,17'd40120,17'd39967,17'd38093,17'd40121,17'd40122,17'd40123,17'd40124,17'd40125,17'd40126,17'd40127,17'd40128,17'd40129,17'd40130,17'd40131,17'd40132,17'd18086,17'd18920,17'd15435,17'd11674,17'd23343,17'd8248,17'd12867,17'd24862,17'd8731,17'd8725,17'd15684,17'd24361,17'd17480,17'd8878,17'd34958,17'd30969,17'd17123,17'd9884,17'd19533,17'd23170,17'd28343,17'd30370,17'd34827,17'd31765,17'd34835,17'd30677,17'd36937,17'd40133,17'd36629,17'd26370,17'd23170,17'd22817,17'd22647,17'd28352,17'd24996,17'd28352,17'd11669,17'd11400,17'd10330,17'd17719,17'd17719,17'd11671,17'd9885,17'd9345,17'd12117,17'd8720,17'd9045,17'd10336,17'd39977,17'd17232,17'd11809,17'd9619,17'd9618,17'd40134,17'd10606,17'd11132,17'd11275,17'd19920,17'd14807,17'd16558,17'd17725,17'd37857,17'd40135,17'd18562,17'd18448,17'd40136,17'd17844,17'd31776,17'd34392,17'd32448,17'd30380,17'd40137,17'd40138,17'd39515,17'd32942,17'd40139,17'd40140,17'd40141,17'd40142,17'd40143,17'd40144,17'd40145,17'd40146,17'd40147,17'd39987,17'd40148,17'd40149,17'd40150,17'd40151,17'd40152,17'd40153,17'd40154,17'd40155,17'd40156,17'd39099,17'd40157,17'd40158,17'd40159,17'd40160,17'd40161,17'd40162,17'd40163,17'd40164,17'd40165,17'd40166,17'd40167,17'd40168,17'd40169,17'd40170,17'd40171,17'd40172,17'd40173,17'd40174,17'd40175,17'd40176,17'd40177,17'd40178,17'd40179,17'd40180,17'd40181,17'd40182,17'd40183,17'd40184,17'd40185,17'd40186,17'd40187,17'd40188,17'd40189,17'd40190,17'd40191,17'd40192,17'd40193,17'd40194,17'd40195,17'd40196,17'd40197,17'd40198,17'd40199,17'd36245,17'd36512,17'd39116,17'd37097,17'd40035,17'd36670,17'd36670,17'd36385,17'd39262,17'd40200,17'd40201,17'd40202,17'd40203,17'd40204,17'd40205,17'd40206,17'd40207,17'd40208,17'd40209,17'd40044,17'd40210,17'd40211,17'd38801,17'd39734,17'd40212,17'd40213,17'd40214,17'd40215,17'd40216,17'd40217,17'd37904,17'd39905,17'd39906,17'd40218,17'd32495,17'd27372,17'd28853,17'd25708,17'd27765,17'd25320,17'd35159,17'd29828,17'd40049,17'd22679,17'd22328,17'd23218,17'd29829,17'd23733,17'd29241,17'd29099,17'd23923,17'd30579,17'd29827,17'd24902,17'd25180,17'd28723,17'd27259,17'd30586,17'd27027,17'd27259,17'd26902,17'd35426,17'd40219,17'd40220,17'd28982,17'd29249,17'd33486,17'd32355,17'd28373,17'd32017,17'd32505,17'd32355,17'd28258,17'd32826,17'd25029,17'd31191,17'd35429,17'd22331,17'd40221,17'd32997,17'd40222,17'd40223,17'd40224,17'd30431,17'd25320,17'd25435,17'd28594,17'd28717,17'd33484,17'd33000,17'd27765,17'd27638,17'd33000,17'd25568,17'd28717,17'd28481,17'd26902,17'd31352,17'd27885,17'd33001,17'd37513,17'd35579,17'd35579,17'd38982,17'd40225,17'd40226,17'd40227,17'd34769,17'd40228,17'd40229,17'd38545,17'd40230,17'd40061,17'd35860,17'd40231,17'd40232,17'd37532,17'd35722,17'd34622,17'd24896,17'd25568,17'd30606,17'd28853,17'd35426,17'd31352,17'd26901,17'd26782,17'd25830,17'd23553,17'd29101,17'd25439,17'd34277,17'd40233,17'd40234,17'd40235,17'd31867,17'd40236,17'd19794,17'd33827,17'd40237,17'd40238,17'd40239,17'd40240,17'd37793,17'd20677,17'd21744,17'd37547,17'd36020,17'd37689,17'd40241,17'd40242,17'd40243,17'd39309,17'd19087,17'd22422,17'd22250,17'd40244,17'd40245,17'd37428,17'd40246,17'd28183,17'd31888,17'd29592,17'd29592,17'd29593,17'd9933,17'd9933,17'd7499,17'd6219,17'd28185,17'd4841,17'd39468,17'd39165,17'd4689,17'd5162,17'd34921,17'd4529,17'd4359,17'd39936,17'd40247,17'd4681,17'd4684,17'd5162,17'd40082,17'd40248,17'd40249,17'd40250,17'd40251,17'd40252,17'd40253,17'd40254,17'd40255,17'd40256,17'd40091,17'd40092,17'd39945,17'd39785,17'd40095,17'd40257,17'd39787,17'd40258,17'd36746,17'd19490,17'd39029,17'd38070,17'd6082,17'd5494,17'd3871,17'd3709,17'd39789,17'd10790,17'd39482,17'd38333,17'd37957,17'd37709,17'd6258,17'd6417,17'd8507,17'd7537,17'd9124,17'd38460,17'd38460,17'd38460,17'd34002,17'd33051,17'd11882,17'd4714,17'd4713,17'd3895,17'd1261,17'd1680,17'd626,17'd627,17'd3100,17'd211,17'd2420,17'd639,17'd1826,17'd22106
},
'{
17'd4428,17'd4088,17'd6420,17'd6420,17'd6420,17'd4245,17'd6420,17'd25384,17'd4245,17'd4246,17'd3252,17'd27714,17'd17917,17'd2,17'd18,17'd3905,17'd3905,17'd3905,17'd27,17'd980,17'd7728,17'd7060,17'd6437,17'd5971,17'd5379,17'd4739,17'd2431,17'd1283,17'd1424,17'd1285,17'd1560,17'd2949,17'd1145,17'd836,17'd38867,17'd40259,17'd2273,17'd13442,17'd4591,17'd5397,17'd38585,17'd35912,17'd40104,17'd40105,17'd40106,17'd18175,17'd19257,17'd18656,17'd18774,17'd18655,17'd17941,17'd19388,17'd21040,17'd40260,17'd40261,17'd40262,17'd40263,17'd40264,17'd40265,17'd40111,17'd40112,17'd40112,17'd40113,17'd40266,17'd40114,17'd40267,17'd40268,17'd37718,17'd39963,17'd40116,17'd39052,17'd36054,17'd39645,17'd14358,17'd9848,17'd9014,17'd8851,17'd40269,17'd24978,17'd39502,17'd6780,17'd40270,17'd40271,17'd40119,17'd39816,17'd39813,17'd6485,17'd40272,17'd40273,17'd40274,17'd38093,17'd40275,17'd40276,17'd40277,17'd40278,17'd40279,17'd40280,17'd40127,17'd40128,17'd40281,17'd40282,17'd6809,17'd40283,17'd18086,17'd15692,17'd15435,17'd11674,17'd23343,17'd8248,17'd10339,17'd24545,17'd12425,17'd8879,17'd15684,17'd24361,17'd14811,17'd10027,17'd34958,17'd9482,17'd15430,17'd9883,17'd24029,17'd24209,17'd28343,17'd30370,17'd34827,17'd30676,17'd34381,17'd30677,17'd29785,17'd31286,17'd30218,17'd26371,17'd21363,17'd30532,17'd22647,17'd28352,17'd19532,17'd28352,17'd11669,17'd11525,17'd11526,17'd10329,17'd17719,17'd11671,17'd9741,17'd9345,17'd12117,17'd8873,17'd29334,17'd22813,17'd15807,17'd9479,17'd16549,17'd9619,17'd9739,17'd10164,17'd10991,17'd11132,17'd11808,17'd19920,17'd14807,17'd16558,17'd18685,17'd40135,17'd40135,17'd17724,17'd17724,17'd40136,17'd40284,17'd30839,17'd40285,17'd33418,17'd40286,17'd40137,17'd32934,17'd40287,17'd40288,17'd10325,17'd40289,17'd40290,17'd40291,17'd40292,17'd40293,17'd40294,17'd40295,17'd40147,17'd40296,17'd40297,17'd40149,17'd40298,17'd40299,17'd40300,17'd40301,17'd40302,17'd40303,17'd40304,17'd40305,17'd40306,17'd40307,17'd40308,17'd40309,17'd40310,17'd40311,17'd40312,17'd40313,17'd40314,17'd40315,17'd40316,17'd40317,17'd40318,17'd40319,17'd40320,17'd40321,17'd40322,17'd40323,17'd40324,17'd40325,17'd40326,17'd40327,17'd40328,17'd40329,17'd40330,17'd40331,17'd40332,17'd40333,17'd40334,17'd40335,17'd40336,17'd40337,17'd40338,17'd40339,17'd40340,17'd40341,17'd40342,17'd40343,17'd40344,17'd40345,17'd40346,17'd40347,17'd40348,17'd37101,17'd40349,17'd40350,17'd36820,17'd39261,17'd37367,17'd36244,17'd36384,17'd36385,17'd38262,17'd40351,17'd40352,17'd40353,17'd40354,17'd40355,17'd40356,17'd40357,17'd39268,17'd39894,17'd40358,17'd39124,17'd40359,17'd40360,17'd38968,17'd38533,17'd40361,17'd40362,17'd40363,17'd40364,17'd40217,17'd37904,17'd40365,17'd40366,17'd39907,17'd32495,17'd27372,17'd28853,17'd25708,17'd27765,17'd29244,17'd32659,17'd32191,17'd40049,17'd22679,17'd22501,17'd23217,17'd30579,17'd23733,17'd31033,17'd23565,17'd23386,17'd29530,17'd23566,17'd28722,17'd25178,17'd26064,17'd28725,17'd30586,17'd26902,17'd27640,17'd28853,17'd36690,17'd35425,17'd38154,17'd28982,17'd29249,17'd33486,17'd32355,17'd28373,17'd32017,17'd32505,17'd32355,17'd40367,17'd33309,17'd24897,17'd39587,17'd31496,17'd22330,17'd40368,17'd32997,17'd34757,17'd40369,17'd40370,17'd29375,17'd25179,17'd28600,17'd28594,17'd31366,17'd33484,17'd33000,17'd28130,17'd28594,17'd31055,17'd33484,17'd28717,17'd28481,17'd26902,17'd31352,17'd30279,17'd33001,17'd40371,17'd39284,17'd35579,17'd38982,17'd38982,17'd36001,17'd40226,17'd39749,17'd40228,17'd40229,17'd33502,17'd40372,17'd40373,17'd35995,17'd40374,17'd40375,17'd40376,17'd40377,17'd40378,17'd24417,17'd28254,17'd27638,17'd28978,17'd35426,17'd29379,17'd28726,17'd26902,17'd25702,17'd25708,17'd40379,17'd30446,17'd33971,17'd40380,17'd40381,17'd40382,17'd40383,17'd40384,17'd40385,17'd40386,17'd40387,17'd40388,17'd40389,17'd23609,17'd40390,17'd22555,17'd38051,17'd39461,17'd36164,17'd40391,17'd40392,17'd40242,17'd40393,17'd22251,17'd19087,17'd18619,17'd21772,17'd40244,17'd40245,17'd37428,17'd40394,17'd28057,17'd31888,17'd29592,17'd27933,17'd29592,17'd9933,17'd8780,17'd6220,17'd6219,17'd27935,17'd5328,17'd4356,17'd40395,17'd5156,17'd5162,17'd5157,17'd4529,17'd4190,17'd39773,17'd40396,17'd4681,17'd40397,17'd5157,17'd40398,17'd40399,17'd40400,17'd34916,17'd40401,17'd40402,17'd40403,17'd40404,17'd40405,17'd40256,17'd40406,17'd40092,17'd39945,17'd39785,17'd40095,17'd40257,17'd39787,17'd40407,17'd40097,17'd2236,17'd40408,17'd40409,17'd40410,17'd4394,17'd3870,17'd40411,17'd39789,17'd10790,17'd39482,17'd40101,17'd38860,17'd38861,17'd39791,17'd6417,17'd8507,17'd7537,17'd9124,17'd38460,17'd38460,17'd38460,17'd33051,17'd33051,17'd11061,17'd11335,17'd4869,17'd5193,17'd229,17'd1261,17'd446,17'd623,17'd233,17'd40412,17'd211,17'd1682,17'd186,17'd404
},
'{
17'd4428,17'd4088,17'd6420,17'd25384,17'd6420,17'd6420,17'd6420,17'd25384,17'd14743,17'd4246,17'd3252,17'd27714,17'd2594,17'd2,17'd18,17'd20404,17'd3905,17'd4089,17'd27,17'd980,17'd7728,17'd6745,17'd6437,17'd3910,17'd5379,17'd4739,17'd2431,17'd1704,17'd1705,17'd1285,17'd1560,17'd1427,17'd998,17'd1290,17'd38867,17'd40103,17'd22970,17'd27102,17'd4591,17'd40413,17'd18525,17'd40414,17'd40104,17'd40105,17'd40415,17'd17810,17'd19008,17'd17206,17'd18774,17'd19892,17'd17204,17'd20024,17'd18416,17'd36612,17'd38083,17'd40416,17'd40417,17'd38879,17'd40418,17'd40419,17'd40420,17'd40421,17'd40422,17'd40266,17'd39961,17'd39498,17'd38472,17'd37717,17'd40423,17'd40424,17'd39501,17'd34367,17'd16778,17'd14358,17'd19900,17'd9581,17'd9013,17'd8849,17'd24977,17'd7758,17'd6780,17'd40270,17'd40271,17'd40120,17'd39813,17'd39813,17'd40425,17'd40426,17'd40427,17'd40428,17'd38603,17'd38482,17'd6949,17'd40429,17'd40430,17'd40431,17'd40432,17'd40433,17'd40434,17'd6799,17'd40435,17'd40436,17'd40437,17'd21366,17'd15692,17'd15435,17'd17353,17'd23343,17'd8248,17'd14812,17'd8571,17'd8729,17'd8879,17'd9194,17'd17716,17'd14811,17'd8410,17'd40438,17'd8726,17'd24361,17'd11134,17'd11397,17'd24031,17'd28227,17'd30370,17'd29330,17'd36491,17'd31773,17'd31765,17'd31587,17'd40439,17'd40440,17'd24859,17'd21362,17'd30532,17'd14263,17'd19532,17'd19532,17'd11669,17'd21206,17'd11669,17'd24996,17'd10166,17'd17124,17'd9883,17'd9741,17'd9345,17'd12117,17'd8873,17'd8720,17'd8874,17'd15807,17'd9479,17'd12116,17'd9740,17'd9740,17'd10164,17'd11133,17'd10475,17'd11808,17'd13646,17'd12580,17'd14524,17'd17013,17'd40441,17'd40442,17'd17349,17'd17349,17'd40284,17'd40443,17'd40444,17'd36784,17'd34393,17'd40445,17'd18683,17'd32934,17'd32942,17'd40446,17'd40447,17'd40448,17'd40449,17'd40450,17'd39984,17'd40451,17'd39522,17'd39837,17'd40452,17'd40453,17'd40297,17'd40149,17'd40150,17'd40454,17'd40455,17'd40456,17'd40457,17'd40458,17'd40459,17'd40460,17'd40461,17'd40462,17'd40463,17'd40464,17'd40465,17'd40466,17'd40467,17'd40468,17'd40469,17'd40470,17'd40471,17'd40472,17'd40473,17'd40474,17'd40475,17'd40476,17'd40477,17'd40478,17'd40479,17'd40480,17'd40481,17'd40482,17'd40483,17'd40484,17'd40485,17'd40486,17'd40487,17'd40488,17'd40489,17'd40490,17'd40491,17'd40492,17'd40493,17'd40494,17'd40495,17'd39995,17'd40496,17'd40497,17'd40498,17'd39884,17'd40499,17'd40500,17'd40501,17'd40502,17'd37637,17'd40349,17'd36820,17'd36964,17'd37634,17'd38391,17'd36244,17'd36384,17'd38389,17'd37638,17'd40503,17'd40504,17'd40505,17'd40506,17'd40507,17'd40508,17'd40509,17'd40510,17'd40511,17'd40512,17'd40513,17'd40514,17'd38968,17'd38533,17'd40515,17'd40516,17'd40517,17'd40518,17'd40519,17'd40365,17'd39739,17'd40366,17'd39907,17'd40520,17'd32343,17'd28853,17'd25708,17'd27765,17'd29244,17'd32659,17'd23388,17'd40049,17'd39131,17'd22502,17'd23218,17'd23567,17'd23920,17'd29241,17'd29376,17'd23923,17'd30579,17'd23566,17'd30879,17'd25179,17'd28720,17'd28724,17'd27146,17'd26902,17'd27640,17'd28853,17'd33941,17'd35990,17'd38154,17'd32018,17'd29249,17'd33486,17'd32355,17'd28134,17'd32017,17'd32355,17'd32355,17'd40367,17'd33310,17'd24417,17'd39908,17'd32660,17'd22500,17'd40521,17'd21694,17'd40522,17'd32012,17'd40523,17'd33801,17'd30432,17'd28130,17'd30606,17'd33000,17'd28717,17'd28597,17'd28594,17'd30606,17'd28599,17'd28717,17'd33000,17'd28481,17'd26902,17'd29245,17'd31503,17'd29977,17'd37513,17'd31503,17'd31503,17'd40524,17'd28011,17'd38160,17'd39286,17'd35167,17'd40525,17'd40526,17'd36867,17'd40230,17'd40373,17'd33504,17'd40527,17'd38412,17'd38410,17'd37532,17'd40378,17'd24743,17'd24897,17'd28597,17'd28724,17'd35426,17'd31352,17'd26901,17'd26902,17'd28725,17'd25833,17'd33510,17'd40528,17'd29376,17'd40529,17'd40530,17'd25037,17'd40531,17'd40532,17'd40533,17'd40534,17'd40535,17'd40536,17'd40537,17'd40538,17'd40539,17'd40540,17'd40541,17'd40542,17'd9213,17'd40543,17'd40544,17'd40242,17'd40545,17'd39770,17'd40546,17'd18619,17'd21772,17'd40244,17'd40245,17'd37556,17'd40394,17'd28057,17'd29593,17'd27933,17'd28183,17'd29592,17'd27815,17'd8780,17'd6391,17'd6220,17'd5614,17'd5328,17'd4185,17'd40547,17'd4525,17'd5162,17'd5157,17'd4529,17'd4524,17'd40548,17'd39165,17'd4360,17'd4526,17'd4846,17'd40549,17'd40399,17'd40550,17'd40551,17'd40552,17'd40553,17'd40554,17'd40555,17'd40556,17'd40256,17'd40406,17'd40092,17'd39945,17'd40557,17'd22775,17'd40558,17'd40559,17'd40407,17'd40560,17'd2236,17'd40408,17'd40561,17'd40562,17'd4394,17'd3870,17'd40411,17'd39789,17'd39180,17'd10906,17'd11048,17'd38334,17'd4867,17'd6258,17'd6417,17'd35769,17'd7537,17'd7705,17'd9261,17'd9261,17'd9261,17'd11882,17'd11882,17'd11061,17'd4714,17'd4729,17'd3895,17'd1119,17'd624,17'd626,17'd627,17'd608,17'd40563,17'd2255,17'd2255,17'd2115,17'd40564
},
'{
17'd4428,17'd4088,17'd6420,17'd25384,17'd6420,17'd6420,17'd6420,17'd25384,17'd14743,17'd4246,17'd3252,17'd27714,17'd2594,17'd2,17'd18,17'd20404,17'd3905,17'd4089,17'd27,17'd980,17'd7061,17'd6438,17'd6598,17'd3910,17'd5379,17'd4739,17'd2431,17'd1283,17'd1424,17'd1285,17'd1425,17'd2949,17'd996,17'd1290,17'd2792,17'd2443,17'd39632,17'd2626,17'd39039,17'd40565,17'd17561,17'd40414,17'd40566,17'd40105,17'd40415,17'd17448,17'd19008,17'd27461,17'd19892,17'd19892,17'd19621,17'd20024,17'd18416,17'd40567,17'd40568,17'd40569,17'd39493,17'd40570,17'd40571,17'd40572,17'd40573,17'd40421,17'd40422,17'd40266,17'd39961,17'd40574,17'd38472,17'd37717,17'd40575,17'd40576,17'd38601,17'd40577,17'd14639,17'd18306,17'd19900,17'd40578,17'd39197,17'd8383,17'd40579,17'd7101,17'd7915,17'd40580,17'd40581,17'd40273,17'd39813,17'd40582,17'd40425,17'd40583,17'd40584,17'd40585,17'd40586,17'd6788,17'd39650,17'd40587,17'd40588,17'd40589,17'd40590,17'd40591,17'd40592,17'd40593,17'd40594,17'd6973,17'd40437,17'd21366,17'd15692,17'd15435,17'd17353,17'd23343,17'd8248,17'd24213,17'd12425,17'd8569,17'd15297,17'd9194,17'd25814,17'd24361,17'd40595,17'd40596,17'd8886,17'd24361,17'd11134,17'd11397,17'd24538,17'd28943,17'd30370,17'd31940,17'd39211,17'd36491,17'd30972,17'd29330,17'd29480,17'd40597,17'd24705,17'd14258,17'd22816,17'd14263,17'd19282,17'd28352,17'd13521,17'd28463,17'd21206,17'd19532,17'd10166,17'd17124,17'd9883,17'd9741,17'd9345,17'd12117,17'd9038,17'd9043,17'd9190,17'd10334,17'd18556,17'd12116,17'd9740,17'd9740,17'd10164,17'd11133,17'd10475,17'd11965,17'd13135,17'd12580,17'd14672,17'd16560,17'd17477,17'd40598,17'd17349,17'd17349,17'd40284,17'd40599,17'd40600,17'd40601,17'd30535,17'd40445,17'd16548,17'd32292,17'd40602,17'd40603,17'd40604,17'd40605,17'd40606,17'd40607,17'd40292,17'd35660,17'd40608,17'd40609,17'd40610,17'd40611,17'd40612,17'd40613,17'd40614,17'd40615,17'd40616,17'd35824,17'd40617,17'd40618,17'd40619,17'd40620,17'd40621,17'd40622,17'd40623,17'd40624,17'd40625,17'd40626,17'd40627,17'd40628,17'd40629,17'd40630,17'd40473,17'd40631,17'd40632,17'd40633,17'd40634,17'd40635,17'd40635,17'd40636,17'd40637,17'd40638,17'd40639,17'd40640,17'd40641,17'd40642,17'd40643,17'd40644,17'd40645,17'd40646,17'd40647,17'd40648,17'd40649,17'd40650,17'd40651,17'd40652,17'd40653,17'd40654,17'd40655,17'd40656,17'd40657,17'd40498,17'd40658,17'd40659,17'd40660,17'd40661,17'd34734,17'd35684,17'd36243,17'd37226,17'd36669,17'd36669,17'd36670,17'd36384,17'd38389,17'd40662,17'd40663,17'd40664,17'd40665,17'd40666,17'd40667,17'd40668,17'd40669,17'd40361,17'd40670,17'd40671,17'd40672,17'd39124,17'd38968,17'd38533,17'd40673,17'd40674,17'd40675,17'd40676,17'd40519,17'd37508,17'd40365,17'd40366,17'd39907,17'd39741,17'd32496,17'd27258,17'd25708,17'd27765,17'd29244,17'd32659,17'd23388,17'd40049,17'd39131,17'd33158,17'd23217,17'd38806,17'd23920,17'd24086,17'd23565,17'd29827,17'd29530,17'd23566,17'd23731,17'd25320,17'd26064,17'd28725,17'd30586,17'd28853,17'd27514,17'd28978,17'd33476,17'd40677,17'd28858,17'd32018,17'd29249,17'd33486,17'd32355,17'd28134,17'd33654,17'd32355,17'd32355,17'd40367,17'd33310,17'd24743,17'd40678,17'd22157,17'd33315,17'd36846,17'd21693,17'd34616,17'd33798,17'd40679,17'd40680,17'd38667,17'd28130,17'd28602,17'd33000,17'd28717,17'd28597,17'd28720,17'd26064,17'd38671,17'd31366,17'd31055,17'd28482,17'd26902,17'd29245,17'd29977,17'd40681,17'd40371,17'd30279,17'd31354,17'd40524,17'd40524,17'd38982,17'd36001,17'd39749,17'd40525,17'd40526,17'd36867,17'd40230,17'd40373,17'd37913,17'd40682,17'd38412,17'd40683,17'd40684,17'd40685,17'd24089,17'd24744,17'd25709,17'd28252,17'd35426,17'd31352,17'd26901,17'd26902,17'd28725,17'd25833,17'd26661,17'd25710,17'd23732,17'd38040,17'd40686,17'd40687,17'd40688,17'd40689,17'd40236,17'd40690,17'd40691,17'd40692,17'd40693,17'd40694,17'd40695,17'd40696,17'd40697,17'd37418,17'd35467,17'd36304,17'd40698,17'd40242,17'd40545,17'd39770,17'd18741,17'd18619,17'd18021,17'd40244,17'd40245,17'd38845,17'd40699,17'd27934,17'd29592,17'd27933,17'd28183,17'd29592,17'd9933,17'd8780,17'd6220,17'd6220,17'd5614,17'd5328,17'd5476,17'd40700,17'd4999,17'd5162,17'd4846,17'd4529,17'd4524,17'd40548,17'd39313,17'd4360,17'd4526,17'd4847,17'd40549,17'd40701,17'd40702,17'd34787,17'd40703,17'd40704,17'd40705,17'd40706,17'd40707,17'd40708,17'd40709,17'd40710,17'd39945,17'd40711,17'd3046,17'd40558,17'd40712,17'd40713,17'd40714,17'd36746,17'd19237,17'd40561,17'd40715,17'd4054,17'd4055,17'd40411,17'd39947,17'd18629,17'd40716,17'd40101,17'd38860,17'd38072,17'd16492,17'd6417,17'd35769,17'd8507,17'd7705,17'd9261,17'd9261,17'd7705,17'd11882,17'd11882,17'd11061,17'd11335,17'd5194,17'd40717,17'd40718,17'd228,17'd625,17'd626,17'd1539,17'd40563,17'd40563,17'd595,17'd265,17'd189
},
'{
17'd4088,17'd4088,17'd6420,17'd25384,17'd25384,17'd6420,17'd6420,17'd25384,17'd14743,17'd4246,17'd3252,17'd10535,17'd2594,17'd13,17'd1128,17'd20404,17'd3905,17'd4089,17'd27,17'd27444,17'd7225,17'd40719,17'd6437,17'd3910,17'd5210,17'd2946,17'd2431,17'd1704,17'd1705,17'd1285,17'd1425,17'd1427,17'd835,17'd2614,17'd2792,17'd2443,17'd29307,17'd14876,17'd5232,17'd40565,17'd17561,17'd40414,17'd40566,17'd35350,17'd40415,17'd17448,17'd18656,17'd18774,17'd20422,17'd20422,17'd39797,17'd19756,17'd18416,17'd40720,17'd15906,17'd39492,17'd40721,17'd40722,17'd40723,17'd40724,17'd40725,17'd40726,17'd39804,17'd39960,17'd39806,17'd40574,17'd38472,17'd37833,17'd40727,17'd40728,17'd38091,17'd39964,17'd16665,17'd18179,17'd9581,17'd40729,17'd9013,17'd8383,17'd40579,17'd7100,17'd7915,17'd40730,17'd40731,17'd40273,17'd40583,17'd40732,17'd40732,17'd40120,17'd40733,17'd40585,17'd40586,17'd40734,17'd40735,17'd40587,17'd40736,17'd40737,17'd40738,17'd40739,17'd40592,17'd40740,17'd40741,17'd40742,17'd40437,17'd22301,17'd15692,17'd15435,17'd8580,17'd19923,17'd9483,17'd9349,17'd8569,17'd8886,17'd9348,17'd8873,17'd18080,17'd15944,17'd15178,17'd32921,17'd9040,17'd14674,17'd11134,17'd11964,17'd24859,17'd28943,17'd30370,17'd29330,17'd30220,17'd37335,17'd31440,17'd29067,17'd29923,17'd25527,17'd25926,17'd18681,17'd22816,17'd14263,17'd19282,17'd19532,17'd11669,17'd28463,17'd21206,17'd19532,17'd10023,17'd20044,17'd17719,17'd9740,17'd27856,17'd12117,17'd9039,17'd8873,17'd9189,17'd15807,17'd11809,17'd12116,17'd9740,17'd20044,17'd10163,17'd10855,17'd10475,17'd11965,17'd11963,17'd13519,17'd13643,17'd31599,17'd40743,17'd39979,17'd17233,17'd40744,17'd17349,17'd31775,17'd32446,17'd31777,17'd40745,17'd40746,17'd18682,17'd29203,17'd40602,17'd40747,17'd40748,17'd40749,17'd40750,17'd40751,17'd40292,17'd35660,17'd40608,17'd40752,17'd40753,17'd40754,17'd40755,17'd40756,17'd40757,17'd40758,17'd40759,17'd40760,17'd40761,17'd40762,17'd40763,17'd40764,17'd40765,17'd40766,17'd40767,17'd40768,17'd40769,17'd40770,17'd40771,17'd40772,17'd40773,17'd40774,17'd40775,17'd40776,17'd40777,17'd40636,17'd40778,17'd40779,17'd40779,17'd40780,17'd40781,17'd40782,17'd40638,17'd40783,17'd40784,17'd40785,17'd40786,17'd40787,17'd40788,17'd40789,17'd40790,17'd40791,17'd40792,17'd40793,17'd40794,17'd40795,17'd40796,17'd40797,17'd40798,17'd40799,17'd40800,17'd40801,17'd40802,17'd40803,17'd40804,17'd40805,17'd35399,17'd40806,17'd35405,17'd36243,17'd36669,17'd38391,17'd38391,17'd36244,17'd38645,17'd40807,17'd40808,17'd40809,17'd40810,17'd40811,17'd39893,17'd40812,17'd40813,17'd40814,17'd40357,17'd40815,17'd40816,17'd40817,17'd39126,17'd40818,17'd40819,17'd40820,17'd40821,17'd40676,17'd40822,17'd38665,17'd40823,17'd40824,17'd40825,17'd40218,17'd32185,17'd27258,17'd25708,17'd27765,17'd25320,17'd32659,17'd23388,17'd40049,17'd36426,17'd22501,17'd23215,17'd24421,17'd23920,17'd23920,17'd29099,17'd29827,17'd29530,17'd29376,17'd23917,17'd25179,17'd28594,17'd28724,17'd27258,17'd28725,17'd26530,17'd29535,17'd37777,17'd40677,17'd33320,17'd32018,17'd29249,17'd33486,17'd33485,17'd28134,17'd33654,17'd32017,17'd32017,17'd40367,17'd40826,17'd24743,17'd40827,17'd22157,17'd33315,17'd37115,17'd32010,17'd34616,17'd22338,17'd40223,17'd23567,17'd33793,17'd28600,17'd27766,17'd28597,17'd25709,17'd25567,17'd28723,17'd26062,17'd40828,17'd31055,17'd28599,17'd26530,17'd27027,17'd29245,17'd27642,17'd26652,17'd25697,17'd31354,17'd31354,17'd36555,17'd40524,17'd28011,17'd40227,17'd35167,17'd40525,17'd40229,17'd38822,17'd40829,17'd30002,17'd40830,17'd40831,17'd40832,17'd38543,17'd38542,17'd37256,17'd30879,17'd24416,17'd25028,17'd26285,17'd27369,17'd26524,17'd26901,17'd26902,17'd28725,17'd26903,17'd32364,17'd27511,17'd23382,17'd40833,17'd40834,17'd40835,17'd40836,17'd40837,17'd40384,17'd40838,17'd33026,17'd40839,17'd40840,17'd36573,17'd38835,17'd21114,17'd40841,17'd40842,17'd40843,17'd39305,17'd40844,17'd40845,17'd39308,17'd22251,17'd18134,17'd18498,17'd18021,17'd40846,17'd40847,17'd38845,17'd36171,17'd30639,17'd28533,17'd28306,17'd30933,17'd29592,17'd9933,17'd8780,17'd6219,17'd6219,17'd6853,17'd4684,17'd40848,17'd40849,17'd4189,17'd34921,17'd4846,17'd4689,17'd4999,17'd40548,17'd39313,17'd4190,17'd5000,17'd4529,17'd4691,17'd40701,17'd40850,17'd34652,17'd40851,17'd40852,17'd40853,17'd40854,17'd40707,17'd40855,17'd40406,17'd40092,17'd40856,17'd40711,17'd3046,17'd40558,17'd40857,17'd40858,17'd40714,17'd40859,17'd19237,17'd40860,17'd40861,17'd4224,17'd4055,17'd4056,17'd39947,17'd39180,17'd18383,17'd11048,17'd38334,17'd4867,17'd6095,17'd6095,17'd35769,17'd8507,17'd7705,17'd7705,17'd9261,17'd7705,17'd11882,17'd11882,17'd11061,17'd9123,17'd4729,17'd229,17'd228,17'd625,17'd2249,17'd626,17'd1539,17'd408,17'd802,17'd802,17'd40862,17'd40863
},
'{
17'd4088,17'd4088,17'd6420,17'd25384,17'd25384,17'd6420,17'd6420,17'd25384,17'd14743,17'd4246,17'd2422,17'd10535,17'd2594,17'd2,17'd18,17'd20404,17'd3905,17'd3905,17'd27,17'd1278,17'd7061,17'd6438,17'd5971,17'd3910,17'd5210,17'd2946,17'd2431,17'd1283,17'd1424,17'd1285,17'd1425,17'd2949,17'd996,17'd2615,17'd2618,17'd2443,17'd29307,17'd2626,17'd39039,17'd25507,17'd15371,17'd36186,17'd36187,17'd35350,17'd32738,17'd17448,17'd18656,17'd18774,17'd20422,17'd19382,17'd19755,17'd40864,17'd20429,17'd17099,17'd40865,17'd40866,17'd40867,17'd39956,17'd40572,17'd40724,17'd40868,17'd40726,17'd39804,17'd40869,17'd40870,17'd40574,17'd38472,17'd34185,17'd40727,17'd40871,17'd37589,17'd39964,17'd16665,17'd18179,17'd9581,17'd9013,17'd9162,17'd27327,17'd7757,17'd40872,17'd40873,17'd40874,17'd40581,17'd40273,17'd40732,17'd40732,17'd40732,17'd40875,17'd40733,17'd40876,17'd40877,17'd40878,17'd40879,17'd40880,17'd6793,17'd40881,17'd40882,17'd40883,17'd40592,17'd6660,17'd40884,17'd40742,17'd40437,17'd19537,17'd18920,17'd17016,17'd10028,17'd19923,17'd9483,17'd11404,17'd8569,17'd8886,17'd9348,17'd9039,17'd18080,17'd10174,17'd15178,17'd30523,17'd16067,17'd22814,17'd11134,17'd11396,17'd26493,17'd28943,17'd30370,17'd31940,17'd31587,17'd36211,17'd29330,17'd31768,17'd30218,17'd29326,17'd26035,17'd19921,17'd11130,17'd14263,17'd19282,17'd28352,17'd13521,17'd28463,17'd21206,17'd19532,17'd10023,17'd20044,17'd17719,17'd12116,17'd9345,17'd12117,17'd15430,17'd8874,17'd9190,17'd10334,17'd18556,17'd11277,17'd9740,17'd26870,17'd10163,17'd10855,17'd10475,17'd11965,17'd13362,17'd14670,17'd14809,17'd31775,17'd40885,17'd40743,17'd40744,17'd30683,17'd40443,17'd40886,17'd32446,17'd34215,17'd40887,17'd40137,17'd19922,17'd29203,17'd40288,17'd10162,17'd40888,17'd40889,17'd40890,17'd40891,17'd40892,17'd35660,17'd40893,17'd40894,17'd40753,17'd40895,17'd40896,17'd40756,17'd40757,17'd40897,17'd40898,17'd40899,17'd40900,17'd40901,17'd40902,17'd40903,17'd40904,17'd40905,17'd40906,17'd40907,17'd40908,17'd40909,17'd40910,17'd40911,17'd40912,17'd40913,17'd40635,17'd40914,17'd40915,17'd40916,17'd40780,17'd40917,17'd40918,17'd40919,17'd40920,17'd40921,17'd40922,17'd40923,17'd40924,17'd40925,17'd40926,17'd40927,17'd40928,17'd40929,17'd40930,17'd40931,17'd40932,17'd40933,17'd40934,17'd40935,17'd40936,17'd40937,17'd40938,17'd40339,17'd40939,17'd40940,17'd40941,17'd40942,17'd40943,17'd33762,17'd40944,17'd40945,17'd36106,17'd36105,17'd36384,17'd37634,17'd38391,17'd36670,17'd35972,17'd40946,17'd40947,17'd37236,17'd40948,17'd40949,17'd40950,17'd40951,17'd40952,17'd39122,17'd40953,17'd40213,17'd40954,17'd40817,17'd39126,17'd40955,17'd40956,17'd40820,17'd40821,17'd40957,17'd40822,17'd36686,17'd38536,17'd40958,17'd40959,17'd40218,17'd32185,17'd27258,17'd25708,17'd27765,17'd25320,17'd29688,17'd23388,17'd39908,17'd36426,17'd23215,17'd30128,17'd40960,17'd29241,17'd24086,17'd23918,17'd23566,17'd29530,17'd34137,17'd24415,17'd25320,17'd30606,17'd28725,17'd26902,17'd28725,17'd27514,17'd31827,17'd40961,17'd40677,17'd33320,17'd29249,17'd33166,17'd33486,17'd28373,17'd28134,17'd33654,17'd32017,17'd32017,17'd32506,17'd40826,17'd24252,17'd40962,17'd30580,17'd22325,17'd33650,17'd22338,17'd33481,17'd22511,17'd40963,17'd23216,17'd40964,17'd25435,17'd25708,17'd28597,17'd25709,17'd25567,17'd28723,17'd26062,17'd40965,17'd28599,17'd28598,17'd26530,17'd27027,17'd28727,17'd33952,17'd27636,17'd40966,17'd27885,17'd31354,17'd36555,17'd40967,17'd28011,17'd39286,17'd35167,17'd40525,17'd40229,17'd40968,17'd40829,17'd40969,17'd38827,17'd36699,17'd40970,17'd38543,17'd38542,17'd37256,17'd23732,17'd23916,17'd27509,17'd24242,17'd25553,17'd26525,17'd28486,17'd26782,17'd28725,17'd26903,17'd33970,17'd28369,17'd24590,17'd32351,17'd40971,17'd40972,17'd25443,17'd40973,17'd40974,17'd40975,17'd40976,17'd19549,17'd40977,17'd40978,17'd40979,17'd22904,17'd40980,17'd40981,17'd36577,17'd40982,17'd40983,17'd40984,17'd39308,17'd22251,17'd18134,17'd18498,17'd19478,17'd40244,17'd40985,17'd39013,17'd38701,17'd30488,17'd28650,17'd28306,17'd31243,17'd29593,17'd9933,17'd8780,17'd6554,17'd6390,17'd6853,17'd4847,17'd4829,17'd40986,17'd33838,17'd5157,17'd4846,17'd4689,17'd4525,17'd40987,17'd40548,17'd4359,17'd5000,17'd4689,17'd40988,17'd40701,17'd40989,17'd40990,17'd40991,17'd40992,17'd40993,17'd40994,17'd40995,17'd40708,17'd40996,17'd39944,17'd40856,17'd40711,17'd3046,17'd40558,17'd40857,17'd40997,17'd2546,17'd40560,17'd40998,17'd40999,17'd41000,17'd41001,17'd4055,17'd5493,17'd41002,17'd41003,17'd41004,17'd40101,17'd38860,17'd38072,17'd37959,17'd6095,17'd35769,17'd8507,17'd7705,17'd7705,17'd7705,17'd7705,17'd11882,17'd11882,17'd11061,17'd5029,17'd5194,17'd40717,17'd40718,17'd228,17'd625,17'd626,17'd607,17'd17787,17'd802,17'd41005,17'd7539,17'd41006
},
'{
17'd4088,17'd4088,17'd6420,17'd25384,17'd25384,17'd6420,17'd6420,17'd25384,17'd4246,17'd4887,17'd2422,17'd10535,17'd4247,17'd13,17'd1128,17'd20404,17'd18,17'd3905,17'd27,17'd41007,17'd7225,17'd40719,17'd6438,17'd3910,17'd4250,17'd2946,17'd41008,17'd1704,17'd1705,17'd1285,17'd1425,17'd1427,17'd835,17'd2615,17'd2618,17'd2443,17'd29307,17'd3928,17'd41009,17'd25507,17'd38869,17'd41010,17'd41011,17'd35350,17'd32738,17'd27219,17'd25512,17'd19753,17'd20422,17'd19006,17'd7746,17'd20025,17'd19015,17'd16662,17'd38877,17'd40866,17'd40264,17'd41012,17'd41013,17'd40724,17'd40868,17'd40726,17'd41014,17'd41015,17'd40870,17'd40574,17'd38087,17'd41016,17'd40727,17'd39644,17'd41017,17'd41018,17'd17456,17'd18179,17'd9581,17'd9443,17'd8696,17'd27327,17'd7757,17'd41019,17'd7915,17'd40874,17'd40581,17'd41020,17'd40732,17'd40732,17'd41021,17'd41020,17'd41022,17'd41023,17'd40877,17'd41024,17'd6790,17'd41025,17'd6793,17'd41026,17'd41027,17'd40883,17'd41028,17'd6660,17'd40884,17'd41029,17'd41030,17'd21991,17'd41031,17'd16690,17'd19780,17'd8578,17'd9349,17'd8409,17'd9046,17'd9040,17'd8721,17'd15430,17'd15569,17'd8874,17'd40595,17'd15568,17'd24999,17'd16065,17'd10164,17'd13762,17'd24537,17'd30831,17'd34696,17'd29924,17'd29067,17'd36211,17'd28686,17'd28461,17'd30218,17'd28817,17'd20608,17'd19921,17'd11130,17'd16555,17'd19282,17'd19282,17'd11669,17'd28463,17'd11399,17'd19282,17'd10023,17'd20044,17'd17719,17'd9740,17'd27856,17'd12117,17'd16553,17'd8874,17'd9190,17'd9479,17'd12116,17'd9739,17'd26870,17'd26870,17'd10325,17'd10855,17'd27859,17'd11129,17'd13362,17'd14002,17'd29208,17'd40886,17'd41032,17'd41033,17'd39360,17'd31600,17'd30683,17'd41034,17'd39980,17'd30087,17'd40887,17'd37741,17'd41035,17'd29203,17'd41036,17'd39666,17'd39832,17'd41037,17'd41038,17'd40891,17'd41039,17'd40451,17'd41040,17'd41041,17'd41042,17'd40895,17'd40896,17'd40756,17'd41043,17'd41044,17'd41045,17'd37756,17'd41046,17'd41047,17'd41048,17'd41049,17'd41050,17'd41051,17'd41052,17'd41053,17'd41054,17'd41055,17'd41056,17'd41057,17'd41058,17'd41059,17'd41060,17'd41061,17'd41062,17'd41063,17'd41064,17'd41065,17'd41066,17'd41067,17'd41068,17'd41069,17'd41070,17'd41071,17'd41072,17'd40635,17'd41073,17'd41074,17'd41075,17'd41076,17'd41077,17'd41078,17'd41079,17'd41080,17'd41081,17'd41082,17'd41083,17'd41084,17'd41085,17'd41086,17'd41087,17'd41088,17'd41089,17'd41090,17'd41091,17'd39410,17'd41092,17'd34589,17'd36521,17'd35839,17'd35972,17'd37634,17'd38391,17'd36670,17'd36384,17'd40946,17'd41093,17'd41094,17'd41095,17'd41096,17'd38963,17'd41097,17'd41098,17'd39267,17'd41099,17'd40510,17'd41100,17'd41101,17'd41102,17'd41103,17'd40956,17'd41104,17'd41105,17'd41106,17'd40822,17'd38665,17'd41107,17'd41108,17'd40959,17'd40218,17'd32826,17'd27258,17'd25708,17'd27765,17'd25178,17'd34621,17'd29686,17'd31191,17'd30425,17'd23218,17'd29974,17'd40960,17'd29241,17'd23920,17'd31502,17'd29376,17'd29530,17'd29376,17'd23917,17'd29976,17'd28594,17'd28724,17'd28725,17'd27259,17'd27514,17'd32006,17'd41109,17'd41110,17'd33320,17'd29248,17'd33486,17'd33486,17'd28373,17'd27885,17'd32354,17'd33654,17'd33321,17'd32506,17'd41111,17'd24742,17'd40962,17'd32497,17'd22331,17'd22860,17'd22511,17'd41112,17'd35015,17'd41113,17'd41114,17'd34106,17'd25435,17'd27766,17'd28597,17'd25709,17'd25567,17'd28723,17'd28482,17'd41115,17'd38671,17'd30734,17'd27514,17'd27027,17'd28727,17'd29379,17'd26652,17'd25697,17'd31354,17'd31354,17'd35707,17'd41116,17'd28374,17'd41117,17'd41118,17'd40525,17'd37009,17'd41119,17'd41120,17'd38679,17'd40374,17'd41121,17'd41122,17'd32852,17'd41123,17'd23921,17'd23565,17'd24083,17'd23547,17'd24077,17'd26167,17'd26525,17'd33163,17'd28725,17'd27259,17'd26903,17'd41124,17'd25317,17'd41125,17'd41126,17'd41127,17'd39452,17'd41128,17'd41129,17'd41130,17'd41131,17'd41132,17'd41133,17'd41134,17'd36432,17'd41135,17'd41136,17'd41137,17'd34325,17'd41138,17'd41139,17'd39306,17'd40984,17'd38843,17'd22251,17'd18134,17'd18498,17'd19478,17'd40846,17'd41140,17'd38439,17'd41141,17'd41142,17'd28650,17'd28650,17'd31243,17'd29593,17'd8780,17'd28058,17'd6554,17'd6390,17'd6853,17'd4847,17'd36166,17'd41143,17'd34157,17'd4846,17'd4846,17'd4689,17'd5000,17'd41144,17'd40548,17'd4359,17'd4525,17'd4526,17'd40988,17'd40701,17'd41145,17'd41146,17'd40991,17'd41147,17'd41148,17'd41149,17'd41150,17'd41151,17'd41152,17'd41153,17'd40856,17'd40711,17'd41154,17'd40558,17'd40857,17'd40997,17'd41155,17'd41156,17'd41157,17'd19489,17'd41158,17'd41001,17'd4055,17'd4056,17'd41159,17'd41160,17'd18383,17'd11048,17'd38334,17'd4867,17'd6095,17'd6095,17'd35769,17'd8507,17'd7705,17'd7705,17'd7705,17'd7705,17'd11882,17'd11882,17'd11061,17'd9123,17'd4729,17'd229,17'd228,17'd625,17'd626,17'd626,17'd607,17'd41161,17'd41005,17'd261,17'd269,17'd18985
},
'{
17'd4088,17'd4088,17'd6420,17'd25384,17'd25384,17'd6420,17'd6420,17'd25384,17'd4246,17'd7545,17'd2422,17'd10535,17'd2595,17'd13,17'd18,17'd20404,17'd18,17'd3905,17'd27,17'd1278,17'd7061,17'd6438,17'd5971,17'd3910,17'd4250,17'd2946,17'd1422,17'd1283,17'd1424,17'd1285,17'd1425,17'd2612,17'd669,17'd41162,17'd2618,17'd30351,17'd41163,17'd41164,17'd41009,17'd5071,17'd38869,17'd41165,17'd41011,17'd33699,17'd32738,17'd19257,17'd25512,17'd19753,17'd20422,17'd19006,17'd19388,17'd20295,17'd18300,17'd41166,17'd41167,17'd38735,17'd41168,17'd41169,17'd41170,17'd40573,17'd41171,17'd41172,17'd41173,17'd41015,17'd39961,17'd39498,17'd41174,17'd41016,17'd40727,17'd39052,17'd36615,17'd41018,17'd17456,17'd18666,17'd9581,17'd9013,17'd8849,17'd8382,17'd7757,17'd41019,17'd7915,17'd40874,17'd40581,17'd41021,17'd40732,17'd40732,17'd41021,17'd41020,17'd41022,17'd41175,17'd6647,17'd41176,17'd41177,17'd41178,17'd41179,17'd41180,17'd41181,17'd41182,17'd41183,17'd41184,17'd41185,17'd41029,17'd41186,17'd21991,17'd15814,17'd16690,17'd19780,17'd25147,17'd17481,17'd8409,17'd25677,17'd9040,17'd8875,17'd16553,17'd15569,17'd9189,17'd40595,17'd30522,17'd15684,17'd16065,17'd11670,17'd14264,17'd26371,17'd30830,17'd30071,17'd29924,17'd29067,17'd29645,17'd28571,17'd29328,17'd29778,17'd41187,17'd20450,17'd18444,17'd11130,17'd16555,17'd19282,17'd28352,17'd13521,17'd28463,17'd11399,17'd19282,17'd10023,17'd9740,17'd17719,17'd12116,17'd9345,17'd12117,17'd24361,17'd8874,17'd9190,17'd17232,17'd16549,17'd11277,17'd9739,17'd10741,17'd17720,17'd10855,17'd16555,17'd25144,17'd13362,17'd14002,17'd29792,17'd41188,17'd40600,17'd41189,17'd31776,17'd40444,17'd30232,17'd41190,17'd41191,17'd30087,17'd41192,17'd37741,17'd41035,17'd41193,17'd41194,17'd41195,17'd41196,17'd41197,17'd41198,17'd41199,17'd41200,17'd41201,17'd41202,17'd41203,17'd41204,17'd40754,17'd41205,17'd41206,17'd41207,17'd41208,17'd41209,17'd41210,17'd41211,17'd41212,17'd41213,17'd41214,17'd41215,17'd41216,17'd41217,17'd41218,17'd41219,17'd41220,17'd41221,17'd41222,17'd41223,17'd41224,17'd41225,17'd41226,17'd41227,17'd41228,17'd41065,17'd41229,17'd41230,17'd41231,17'd41232,17'd41232,17'd41233,17'd41234,17'd41235,17'd41236,17'd41071,17'd41237,17'd41238,17'd41239,17'd41240,17'd41241,17'd41242,17'd41243,17'd41244,17'd41245,17'd41246,17'd41247,17'd41248,17'd41249,17'd41250,17'd41251,17'd41252,17'd41253,17'd41254,17'd40804,17'd41255,17'd37493,17'd35274,17'd36385,17'd36384,17'd36670,17'd38391,17'd36670,17'd39567,17'd39570,17'd41256,17'd41257,17'd41258,17'd41259,17'd41260,17'd41261,17'd41262,17'd39423,17'd41263,17'd41264,17'd41265,17'd41101,17'd41266,17'd41103,17'd41267,17'd41268,17'd41269,17'd40676,17'd40822,17'd38665,17'd38665,17'd41108,17'd41270,17'd41271,17'd32826,17'd27258,17'd25949,17'd27765,17'd25178,17'd34106,17'd29686,17'd41272,17'd41273,17'd23216,17'd30579,17'd23734,17'd29241,17'd24086,17'd23733,17'd29099,17'd35865,17'd34137,17'd24415,17'd25178,17'd30606,17'd28724,17'd28725,17'd27259,17'd27514,17'd33154,17'd41274,17'd41110,17'd37250,17'd33486,17'd33486,17'd29248,17'd28373,17'd32354,17'd32354,17'd33654,17'd33654,17'd32356,17'd41111,17'd24416,17'd40827,17'd32345,17'd30276,17'd22682,17'd22511,17'd41112,17'd41275,17'd41276,17'd41277,17'd38978,17'd29970,17'd28602,17'd28597,17'd33000,17'd25567,17'd28602,17'd26530,17'd41115,17'd38671,17'd30734,17'd27514,17'd27027,17'd28727,17'd29379,17'd26652,17'd26652,17'd31354,17'd32356,17'd35707,17'd36541,17'd41116,17'd41117,17'd40227,17'd28730,17'd33965,17'd41119,17'd41120,17'd30447,17'd41278,17'd41279,17'd41280,17'd41281,17'd41282,17'd23921,17'd29689,17'd24590,17'd24245,17'd41283,17'd25311,17'd30577,17'd34637,17'd27259,17'd27259,17'd26903,17'd27766,17'd28484,17'd24246,17'd29827,17'd41284,17'd41285,17'd41286,17'd41287,17'd40689,17'd33351,17'd41288,17'd41289,17'd41290,17'd39000,17'd41291,17'd41292,17'd41293,17'd38183,17'd41294,17'd6066,17'd41295,17'd38055,17'd41296,17'd18620,17'd40546,17'd22422,17'd22250,17'd40846,17'd41297,17'd38439,17'd36444,17'd36735,17'd28650,17'd28650,17'd31243,17'd29593,17'd8780,17'd28058,17'd27935,17'd5614,17'd5337,17'd4846,17'd4829,17'd41298,17'd4515,17'd5156,17'd4846,17'd4847,17'd5001,17'd41299,17'd39313,17'd4362,17'd4999,17'd5155,17'd40988,17'd40399,17'd41300,17'd41301,17'd41302,17'd41303,17'd40552,17'd41304,17'd41305,17'd41306,17'd41307,17'd41308,17'd40856,17'd40711,17'd41309,17'd41310,17'd41311,17'd40997,17'd41312,17'd41313,17'd3066,17'd41314,17'd41158,17'd8786,17'd7849,17'd5493,17'd41315,17'd41003,17'd41004,17'd11048,17'd38334,17'd38072,17'd37959,17'd6095,17'd6417,17'd8507,17'd7705,17'd7705,17'd7705,17'd7705,17'd11882,17'd11882,17'd11061,17'd9123,17'd4729,17'd229,17'd228,17'd624,17'd626,17'd626,17'd1679,17'd41316,17'd261,17'd2779,17'd206,17'd2577
},
'{
17'd4245,17'd4245,17'd4892,17'd4243,17'd4892,17'd4892,17'd25384,17'd6420,17'd2935,17'd3252,17'd1831,17'd2594,17'd1416,17'd18,17'd18,17'd3905,17'd3905,17'd18,17'd980,17'd26,17'd7060,17'd4430,17'd3910,17'd3756,17'd4739,17'd2265,17'd1976,17'd38865,17'd1705,17'd18150,17'd2949,17'd832,17'd486,17'd15631,17'd2618,17'd30351,17'd13442,17'd15249,17'd39951,17'd18160,17'd39486,17'd41165,17'd41317,17'd41318,17'd41319,17'd41320,17'd19007,17'd17689,17'd19382,17'd18884,17'd19388,17'd18416,17'd36612,17'd14898,17'd38469,17'd41321,17'd40570,17'd40572,17'd41322,17'd41323,17'd41323,17'd41172,17'd41324,17'd41015,17'd39961,17'd39498,17'd41174,17'd41325,17'd41326,17'd41327,17'd39345,17'd17816,17'd17456,17'd19267,17'd9443,17'd41328,17'd8849,17'd8381,17'd9011,17'd8691,17'd7914,17'd6632,17'd41329,17'd40732,17'd41330,17'd41021,17'd41020,17'd40584,17'd41331,17'd41332,17'd6647,17'd41176,17'd41333,17'd41334,17'd41335,17'd40432,17'd41336,17'd41337,17'd41338,17'd41339,17'd41340,17'd41341,17'd41342,17'd19288,17'd15693,17'd13258,17'd23343,17'd11967,17'd11404,17'd12425,17'd25677,17'd15684,17'd9038,17'd12117,17'd25814,17'd10174,17'd15428,17'd8883,17'd15944,17'd16549,17'd19280,17'd23513,17'd26493,17'd28943,17'd29329,17'd29645,17'd28686,17'd28571,17'd29480,17'd28343,17'd27004,17'd23170,17'd20609,17'd41343,17'd22647,17'd14263,17'd14263,17'd22647,17'd11130,17'd11130,17'd11399,17'd19282,17'd9883,17'd16796,17'd10856,17'd12116,17'd9480,17'd9344,17'd13887,17'd9192,17'd9043,17'd15807,17'd16549,17'd11277,17'd12116,17'd9883,17'd10326,17'd16555,17'd10475,17'd10737,17'd11963,17'd18081,17'd14521,17'd35520,17'd31449,17'd31139,17'd32936,17'd41344,17'd41345,17'd31601,17'd35520,17'd29653,17'd29793,17'd37741,17'd41346,17'd32135,17'd41194,17'd41347,17'd41348,17'd41038,17'd41349,17'd41350,17'd41200,17'd40293,17'd41351,17'd41352,17'd41353,17'd41354,17'd41355,17'd41356,17'd41357,17'd41358,17'd41359,17'd41360,17'd41361,17'd41362,17'd41363,17'd41364,17'd41365,17'd40004,17'd41366,17'd41367,17'd40773,17'd41368,17'd41369,17'd41370,17'd41371,17'd41372,17'd41373,17'd41374,17'd40919,17'd41375,17'd41375,17'd41376,17'd41377,17'd41378,17'd41379,17'd41371,17'd41070,17'd41380,17'd41381,17'd41382,17'd41383,17'd41384,17'd41385,17'd40924,17'd41386,17'd41387,17'd41388,17'd41389,17'd41390,17'd41391,17'd41392,17'd41393,17'd41394,17'd41395,17'd41396,17'd41397,17'd41398,17'd41089,17'd41399,17'd41400,17'd41401,17'd41402,17'd40945,17'd35972,17'd36385,17'd36244,17'd36670,17'd39568,17'd41403,17'd41404,17'd36115,17'd41405,17'd41406,17'd38962,17'd41407,17'd41408,17'd41262,17'd41409,17'd41410,17'd40951,17'd40515,17'd41411,17'd41412,17'd41413,17'd41414,17'd40516,17'd40517,17'd41415,17'd41416,17'd38536,17'd38665,17'd41417,17'd41418,17'd41418,17'd32184,17'd27258,17'd26530,17'd27638,17'd27512,17'd34106,17'd23388,17'd41419,17'd33316,17'd23215,17'd29099,17'd23733,17'd31033,17'd31033,17'd23732,17'd23565,17'd29376,17'd23565,17'd34467,17'd29244,17'd28602,17'd28724,17'd27515,17'd26530,17'd25833,17'd39277,17'd41274,17'd35425,17'd29248,17'd36847,17'd32018,17'd32505,17'd28133,17'd28854,17'd28854,17'd28370,17'd32354,17'd32356,17'd32185,17'd25180,17'd41420,17'd23040,17'd31834,17'd33312,17'd32828,17'd35293,17'd41421,17'd41422,17'd41423,17'd31190,17'd29825,17'd28602,17'd28598,17'd28597,17'd27638,17'd25708,17'd41424,17'd41425,17'd41426,17'd41427,17'd28009,17'd26901,17'd31035,17'd31352,17'd28980,17'd27642,17'd27642,17'd35570,17'd41428,17'd41429,17'd41116,17'd28011,17'd40226,17'd34769,17'd28490,17'd27887,17'd41430,17'd30447,17'd41431,17'd38418,17'd41432,17'd41433,17'd41434,17'd38542,17'd23732,17'd26398,17'd24740,17'd23724,17'd24582,17'd36286,17'd34637,17'd26782,17'd41435,17'd34135,17'd41436,17'd23557,17'd27637,17'd37256,17'd41437,17'd25035,17'd41438,17'd41439,17'd41440,17'd41441,17'd41442,17'd41443,17'd41444,17'd41445,17'd36432,17'd41446,17'd20507,17'd41447,17'd30633,17'd6540,17'd41448,17'd41449,17'd41450,17'd18374,17'd22595,17'd41451,17'd39012,17'd40846,17'd41452,17'd39161,17'd41453,17'd41454,17'd28533,17'd28305,17'd29592,17'd31888,17'd10515,17'd6391,17'd5335,17'd5329,17'd34334,17'd4846,17'd41455,17'd41456,17'd4356,17'd41457,17'd4846,17'd4847,17'd4525,17'd41458,17'd5476,17'd4832,17'd33838,17'd41459,17'd41460,17'd41461,17'd41462,17'd41463,17'd41464,17'd41465,17'd41466,17'd41467,17'd41468,17'd41469,17'd41470,17'd41471,17'd41472,17'd41473,17'd41309,17'd37816,17'd41474,17'd2221,17'd41475,17'd41476,17'd41477,17'd41478,17'd41479,17'd3562,17'd41480,17'd7849,17'd41315,17'd39947,17'd10388,17'd38458,17'd41481,17'd12636,17'd13933,17'd4730,17'd6258,17'd6094,17'd7364,17'd7878,17'd9124,17'd7537,17'd9261,17'd9414,17'd9544,17'd8186,17'd4729,17'd229,17'd228,17'd625,17'd626,17'd627,17'd2924,17'd41316,17'd17661,17'd2779,17'd972,17'd41482
},
'{
17'd4245,17'd4245,17'd4892,17'd4243,17'd4892,17'd4892,17'd25384,17'd6420,17'd2935,17'd3252,17'd1831,17'd2594,17'd1416,17'd18,17'd18,17'd3905,17'd3905,17'd3905,17'd980,17'd26,17'd7060,17'd4430,17'd3910,17'd12335,17'd4739,17'd2265,17'd1976,17'd1423,17'd1424,17'd18150,17'd2437,17'd832,17'd487,17'd2440,17'd2618,17'd30351,17'd13442,17'd4751,17'd41483,17'd18766,17'd41484,17'd41165,17'd41317,17'd41485,17'd27459,17'd41320,17'd19007,17'd17689,17'd19382,17'd20886,17'd19756,17'd18660,17'd41486,17'd38468,17'd40866,17'd41487,17'd41488,17'd40725,17'd41489,17'd41490,17'd41323,17'd41491,17'd41172,17'd41492,17'd39961,17'd41493,17'd41494,17'd41325,17'd41495,17'd41327,17'd41496,17'd17816,17'd17701,17'd41497,17'd9443,17'd8695,17'd8694,17'd24841,17'd9011,17'd8540,17'd7914,17'd6632,17'd41329,17'd41498,17'd41330,17'd41021,17'd41020,17'd40584,17'd41331,17'd41499,17'd6647,17'd41500,17'd41501,17'd41334,17'd41502,17'd41503,17'd41504,17'd41505,17'd39656,17'd39509,17'd41340,17'd41506,17'd11281,17'd19288,17'd15693,17'd13258,17'd24713,17'd11967,17'd9886,17'd8570,17'd16317,17'd15684,17'd8874,17'd12117,17'd25814,17'd10174,17'd15428,17'd41507,17'd10173,17'd12116,17'd11525,17'd23513,17'd26493,17'd28943,17'd31286,17'd36777,17'd29645,17'd28571,17'd28943,17'd28343,17'd26371,17'd23170,17'd23169,17'd22816,17'd22647,17'd14263,17'd22647,17'd22647,17'd11130,17'd11130,17'd21206,17'd19282,17'd10329,17'd16796,17'd9741,17'd12116,17'd9480,17'd9620,17'd9344,17'd9192,17'd9043,17'd15807,17'd16549,17'd19531,17'd9884,17'd10329,17'd19532,17'd19282,17'd10475,17'd10737,17'd11963,17'd18081,17'd29491,17'd41508,17'd30087,17'd33414,17'd32936,17'd32936,17'd39662,17'd41509,17'd29652,17'd29491,17'd41510,17'd18446,17'd41511,17'd32135,17'd25811,17'd41512,17'd41513,17'd41514,17'd41515,17'd41516,17'd41200,17'd41517,17'd41203,17'd41352,17'd41518,17'd41519,17'd40895,17'd35665,17'd41520,17'd41521,17'd41522,17'd41523,17'd41524,17'd41525,17'd41526,17'd41527,17'd41528,17'd41529,17'd41530,17'd41531,17'd41532,17'd40632,17'd41533,17'd41072,17'd41236,17'd41534,17'd41535,17'd41536,17'd41537,17'd41538,17'd41539,17'd41540,17'd41541,17'd41542,17'd41543,17'd41544,17'd41545,17'd41546,17'd41072,17'd41547,17'd41548,17'd41061,17'd40915,17'd40637,17'd41549,17'd41550,17'd41551,17'd41552,17'd41553,17'd41554,17'd41555,17'd41556,17'd41557,17'd41558,17'd41559,17'd41560,17'd41561,17'd41562,17'd41563,17'd41564,17'd39094,17'd41565,17'd41566,17'd41567,17'd36384,17'd36244,17'd36669,17'd39568,17'd41568,17'd41569,17'd36115,17'd41570,17'd41571,17'd41572,17'd41573,17'd41574,17'd41575,17'd40667,17'd41576,17'd41577,17'd41264,17'd41411,17'd41578,17'd41413,17'd41579,17'd41580,17'd39432,17'd41581,17'd41416,17'd41107,17'd38665,17'd41582,17'd41583,17'd41583,17'd32184,17'd27146,17'd27514,17'd27513,17'd27512,17'd34621,17'd23388,17'd41419,17'd23740,17'd32351,17'd29099,17'd23732,17'd23731,17'd23917,17'd24086,17'd23565,17'd29376,17'd23918,17'd34467,17'd25320,17'd26064,17'd28724,17'd27515,17'd28482,17'd25833,17'd32184,17'd41274,17'd40219,17'd29248,17'd36847,17'd29248,17'd32505,17'd28133,17'd28854,17'd28854,17'd28370,17'd33319,17'd31354,17'd36542,17'd25320,17'd41277,17'd36691,17'd32502,17'd32665,17'd32828,17'd41584,17'd21690,17'd41585,17'd41586,17'd41587,17'd39443,17'd28602,17'd27638,17'd28599,17'd27513,17'd25708,17'd41424,17'd41588,17'd41589,17'd41425,17'd35578,17'd26901,17'd31035,17'd31352,17'd28980,17'd27642,17'd27642,17'd35707,17'd41590,17'd41429,17'd41116,17'd41591,17'd40226,17'd34769,17'd28490,17'd27887,17'd41430,17'd28867,17'd41592,17'd41593,17'd41594,17'd41595,17'd41596,17'd41123,17'd23922,17'd28852,17'd23914,17'd24079,17'd23908,17'd29525,17'd34637,17'd33963,17'd41435,17'd34135,17'd38027,17'd23376,17'd25437,17'd41597,17'd41598,17'd33675,17'd41438,17'd41599,17'd41600,17'd40384,17'd32701,17'd41601,17'd41602,17'd41603,17'd40070,17'd41604,17'd41605,17'd41606,17'd41607,17'd41608,17'd41609,17'd41449,17'd41450,17'd18374,17'd22595,17'd41610,17'd39012,17'd40846,17'd18131,17'd18132,17'd37694,17'd41454,17'd28533,17'd28306,17'd29592,17'd31888,17'd27815,17'd7668,17'd25627,17'd5002,17'd34334,17'd5157,17'd41458,17'd41611,17'd41612,17'd41613,17'd4689,17'd4847,17'd4525,17'd41458,17'd5476,17'd4672,17'd33991,17'd41459,17'd41460,17'd41461,17'd41614,17'd4179,17'd33688,17'd41615,17'd33988,17'd41616,17'd41617,17'd41469,17'd41618,17'd41619,17'd39945,17'd41473,17'd41309,17'd37816,17'd41474,17'd41620,17'd41621,17'd41476,17'd41622,17'd3379,17'd41623,17'd41624,17'd41480,17'd7849,17'd41625,17'd41626,17'd41004,17'd38458,17'd38334,17'd12636,17'd13933,17'd13933,17'd6258,17'd6094,17'd7364,17'd7878,17'd9124,17'd7538,17'd9261,17'd9414,17'd8187,17'd8186,17'd4729,17'd229,17'd228,17'd625,17'd626,17'd627,17'd2924,17'd41316,17'd3899,17'd1538,17'd204,17'd41627
},
'{
17'd4245,17'd4245,17'd4892,17'd4243,17'd4892,17'd4892,17'd25384,17'd15746,17'd3252,17'd10535,17'd2594,17'd2595,17'd4089,17'd18,17'd18,17'd3905,17'd3905,17'd20404,17'd3906,17'd26,17'd27444,17'd4430,17'd3910,17'd3435,17'd4739,17'd2265,17'd1976,17'd1704,17'd1705,17'd18150,17'd41628,17'd484,17'd487,17'd2440,17'd2618,17'd2273,17'd14876,17'd4751,17'd41483,17'd18160,17'd39486,17'd41165,17'd41317,17'd41629,17'd41630,17'd25512,17'd18774,17'd17689,17'd19006,17'd28925,17'd39798,17'd18537,17'd17099,17'd15266,17'd41631,17'd41632,17'd40265,17'd41633,17'd41634,17'd41635,17'd41636,17'd41637,17'd40726,17'd41638,17'd39961,17'd39498,17'd41639,17'd41325,17'd41495,17'd38737,17'd41496,17'd41640,17'd16890,17'd41497,17'd9308,17'd41641,17'd41642,17'd24976,17'd41643,17'd8540,17'd7914,17'd6632,17'd41329,17'd41498,17'd41021,17'd41644,17'd41020,17'd40427,17'd41645,17'd41499,17'd41646,17'd41647,17'd41648,17'd41649,17'd41502,17'd41650,17'd41651,17'd41652,17'd39656,17'd39509,17'd41653,17'd41654,17'd7623,17'd15303,17'd10179,17'd24044,17'd24713,17'd11967,17'd9886,17'd12425,17'd25677,17'd15684,17'd8874,17'd13887,17'd25814,17'd10174,17'd41655,17'd9044,17'd15180,17'd12116,17'd11525,17'd23167,17'd26493,17'd29923,17'd31286,17'd29645,17'd28571,17'd28571,17'd28943,17'd28816,17'd26493,17'd23170,17'd23169,17'd22816,17'd22647,17'd11131,17'd22647,17'd22647,17'd11130,17'd11131,17'd11132,17'd10326,17'd9883,17'd21503,17'd9741,17'd12116,17'd9480,17'd9344,17'd15180,17'd9347,17'd9192,17'd15180,17'd16065,17'd19279,17'd11277,17'd11134,17'd11133,17'd19282,17'd10475,17'd10737,17'd13362,17'd41656,17'd29491,17'd34215,17'd41657,17'd39073,17'd41658,17'd41658,17'd32446,17'd32446,17'd35520,17'd29491,17'd41659,17'd18446,17'd41511,17'd32942,17'd10600,17'd41660,17'd41661,17'd41516,17'd41515,17'd41662,17'd41663,17'd40293,17'd41664,17'd41352,17'd41518,17'd41354,17'd41665,17'd41666,17'd41667,17'd41668,17'd41669,17'd41670,17'd41671,17'd41672,17'd41673,17'd41674,17'd41675,17'd41676,17'd41677,17'd41678,17'd41679,17'd41680,17'd41681,17'd40914,17'd41682,17'd41237,17'd41073,17'd41683,17'd41684,17'd41685,17'd41686,17'd41687,17'd41688,17'd41689,17'd41690,17'd41691,17'd41692,17'd41693,17'd41694,17'd41540,17'd41695,17'd41696,17'd41697,17'd41698,17'd41699,17'd41386,17'd41700,17'd41701,17'd41702,17'd41703,17'd41704,17'd41705,17'd41706,17'd41707,17'd41708,17'd41709,17'd41710,17'd41711,17'd41712,17'd41713,17'd41714,17'd41715,17'd33915,17'd41716,17'd36245,17'd38391,17'd37227,17'd37367,17'd38788,17'd41404,17'd41717,17'd41718,17'd41719,17'd41572,17'd41720,17'd41721,17'd41722,17'd41723,17'd41724,17'd41410,17'd41264,17'd41725,17'd41578,17'd41413,17'd41579,17'd41580,17'd39432,17'd41581,17'd41416,17'd41107,17'd38665,17'd41582,17'd41583,17'd41583,17'd32184,17'd27146,17'd27515,17'd27638,17'd28719,17'd34621,17'd23387,17'd32830,17'd23740,17'd23569,17'd29099,17'd30275,17'd23731,17'd23917,17'd24086,17'd23565,17'd29099,17'd23733,17'd23916,17'd25320,17'd26064,17'd26903,17'd27515,17'd27639,17'd25833,17'd40520,17'd41109,17'd35854,17'd29248,17'd33486,17'd29248,17'd32505,17'd28133,17'd28854,17'd28854,17'd28370,17'd33001,17'd31503,17'd32185,17'd32353,17'd40827,17'd22164,17'd31658,17'd41726,17'd33646,17'd41727,17'd21530,17'd41728,17'd41729,17'd23217,17'd41730,17'd28602,17'd27638,17'd28597,17'd27638,17'd27766,17'd26174,17'd27767,17'd41589,17'd41588,17'd35578,17'd26901,17'd28486,17'd30735,17'd28727,17'd29379,17'd27642,17'd36403,17'd41731,17'd41429,17'd41116,17'd40524,17'd41732,17'd41733,17'd41734,17'd27887,17'd41430,17'd41735,17'd41736,17'd41737,17'd41738,17'd41739,17'd41740,17'd41741,17'd35021,17'd29102,17'd24412,17'd23725,17'd24584,17'd28365,17'd33163,17'd33963,17'd34301,17'd27515,17'd41436,17'd26284,17'd31367,17'd41742,17'd35020,17'd24747,17'd41743,17'd41744,17'd41600,17'd41745,17'd41746,17'd41747,17'd41748,17'd41603,17'd38426,17'd41604,17'd36296,17'd22907,17'd33983,17'd41749,17'd41750,17'd41751,17'd41752,17'd18374,17'd20697,17'd41753,17'd41754,17'd40846,17'd40244,17'd39162,17'd39467,17'd37430,17'd28650,17'd28306,17'd29592,17'd31888,17'd27815,17'd6391,17'd5005,17'd4686,17'd29429,17'd5157,17'd39468,17'd41755,17'd41612,17'd41756,17'd4689,17'd5156,17'd4525,17'd41612,17'd4829,17'd4672,17'd4358,17'd33841,17'd4531,17'd41757,17'd41614,17'd41758,17'd33688,17'd41759,17'd41760,17'd41761,17'd41762,17'd41763,17'd41618,17'd41764,17'd41765,17'd41766,17'd41767,17'd37952,17'd41474,17'd41620,17'd41768,17'd41769,17'd41770,17'd3379,17'd41623,17'd41624,17'd41480,17'd6081,17'd5493,17'd41159,17'd10388,17'd38458,17'd38334,17'd38072,17'd13933,17'd14060,17'd6258,17'd6094,17'd7364,17'd7878,17'd9124,17'd7705,17'd9414,17'd9414,17'd8187,17'd4882,17'd3391,17'd1261,17'd625,17'd625,17'd626,17'd623,17'd2924,17'd261,17'd2779,17'd1966,17'd2256,17'd41627
},
'{
17'd4245,17'd4245,17'd4892,17'd4243,17'd4892,17'd4892,17'd25384,17'd6420,17'd2935,17'd2422,17'd1831,17'd4247,17'd1416,17'd18,17'd18,17'd3905,17'd3905,17'd3905,17'd980,17'd3906,17'd27444,17'd4430,17'd3910,17'd3435,17'd2946,17'd19874,17'd1422,17'd1283,17'd1424,17'd18150,17'd41628,17'd484,17'd307,17'd2269,17'd2618,17'd34169,17'd27102,17'd4591,17'd41483,17'd18766,17'd38339,17'd41165,17'd41317,17'd41485,17'd41771,17'd27461,17'd18774,17'd17689,17'd19006,17'd19513,17'd36189,17'd20431,17'd16990,17'd41772,17'd39955,17'd41773,17'd40418,17'd40725,17'd41774,17'd41490,17'd41774,17'd41637,17'd41172,17'd41775,17'd39961,17'd41493,17'd41776,17'd41325,17'd41495,17'd38737,17'd41777,17'd41778,17'd41779,17'd41497,17'd9308,17'd9161,17'd8694,17'd24841,17'd8845,17'd8540,17'd6638,17'd41780,17'd41329,17'd41781,17'd41644,17'd41644,17'd41020,17'd40733,17'd41782,17'd41783,17'd41646,17'd41784,17'd41785,17'd41786,17'd41787,17'd41788,17'd40591,17'd41789,17'd41790,17'd39355,17'd39822,17'd41791,17'd7459,17'd15303,17'd10179,17'd8250,17'd25147,17'd11531,17'd8412,17'd8878,17'd9194,17'd15684,17'd8874,17'd13887,17'd25814,17'd8874,17'd41792,17'd9042,17'd15807,17'd11277,17'd12423,17'd23167,17'd26493,17'd29923,17'd40439,17'd31286,17'd35372,17'd35372,17'd29923,17'd28816,17'd24857,17'd25926,17'd23169,17'd22816,17'd22647,17'd11131,17'd22647,17'd11130,17'd11130,17'd11130,17'd21206,17'd19532,17'd26152,17'd21503,17'd9741,17'd12116,17'd9480,17'd9620,17'd9345,17'd9347,17'd9192,17'd9345,17'd16549,17'd19531,17'd11671,17'd10330,17'd19282,17'd19282,17'd10475,17'd10737,17'd13362,17'd41656,17'd41793,17'd41508,17'd41794,17'd41657,17'd41795,17'd33100,17'd32446,17'd41509,17'd29490,17'd29491,17'd41659,17'd18446,17'd41511,17'd23510,17'd41796,17'd40289,17'd41797,17'd41350,17'd41515,17'd41516,17'd40607,17'd40293,17'd41798,17'd41353,17'd41518,17'd41799,17'd41800,17'd35115,17'd41801,17'd41802,17'd41803,17'd41804,17'd41805,17'd41806,17'd41807,17'd41808,17'd41809,17'd41810,17'd41811,17'd41812,17'd41813,17'd41814,17'd41815,17'd41816,17'd41817,17'd41058,17'd41818,17'd41819,17'd41820,17'd41821,17'd41822,17'd41823,17'd41824,17'd41825,17'd41826,17'd41827,17'd41828,17'd41829,17'd41830,17'd41831,17'd41832,17'd41833,17'd41834,17'd41835,17'd40637,17'd40323,17'd41836,17'd41837,17'd41838,17'd41839,17'd41840,17'd41841,17'd41842,17'd41843,17'd41844,17'd41845,17'd41846,17'd41847,17'd41848,17'd41849,17'd41850,17'd41851,17'd41852,17'd35834,17'd35972,17'd35972,17'd37227,17'd37495,17'd40035,17'd41853,17'd41854,17'd41718,17'd41855,17'd41856,17'd41857,17'd41721,17'd41722,17'd41858,17'd41859,17'd41410,17'd41264,17'd41725,17'd41578,17'd41413,17'd41579,17'd41860,17'd41861,17'd41862,17'd41863,17'd41107,17'd38665,17'd41582,17'd41583,17'd41864,17'd32495,17'd27372,17'd26903,17'd27638,17'd28719,17'd34621,17'd23387,17'd32830,17'd23740,17'd29974,17'd31502,17'd23732,17'd23731,17'd23917,17'd24086,17'd30275,17'd23918,17'd24086,17'd24416,17'd25320,17'd30606,17'd26903,17'd27515,17'd27639,17'd25707,17'd33308,17'd41109,17'd36541,17'd29248,17'd33486,17'd29248,17'd32505,17'd29247,17'd28854,17'd26522,17'd28854,17'd33001,17'd31503,17'd32496,17'd33483,17'd40827,17'd41865,17'd31192,17'd34457,17'd34616,17'd41866,17'd21531,17'd35855,17'd41867,17'd32514,17'd29103,17'd25566,17'd28130,17'd28598,17'd27513,17'd27766,17'd26174,17'd27767,17'd41427,17'd34300,17'd33499,17'd26901,17'd28486,17'd29245,17'd38537,17'd29379,17'd27642,17'd36541,17'd41731,17'd34877,17'd41868,17'd28011,17'd36001,17'd34896,17'd41869,17'd41870,17'd41430,17'd36270,17'd41736,17'd41737,17'd41871,17'd41595,17'd41872,17'd41873,17'd41874,17'd28849,17'd24589,17'd23726,17'd24892,17'd25702,17'd30586,17'd26781,17'd34301,17'd27515,17'd41436,17'd26284,17'd34127,17'd29994,17'd33331,17'd24747,17'd38686,17'd41875,17'd41876,17'd41877,17'd41878,17'd41879,17'd41880,17'd41881,17'd41882,17'd41883,17'd41884,17'd22555,17'd33983,17'd41885,17'd41886,17'd41887,17'd41752,17'd18620,17'd20697,17'd41888,17'd37555,17'd41452,17'd40244,17'd18021,17'd37803,17'd37558,17'd28306,17'd28650,17'd29593,17'd31888,17'd9933,17'd6220,17'd5005,17'd4686,17'd41889,17'd4846,17'd39468,17'd41755,17'd41455,17'd33837,17'd5156,17'd5156,17'd4525,17'd33533,17'd5476,17'd41890,17'd4515,17'd41891,17'd34501,17'd41892,17'd41893,17'd5473,17'd41894,17'd41895,17'd4509,17'd41896,17'd41897,17'd41763,17'd41618,17'd41764,17'd41898,17'd41899,17'd41900,17'd37952,17'd41901,17'd41620,17'd41902,17'd2726,17'd3059,17'd41903,17'd41904,17'd4052,17'd41905,17'd41906,17'd41907,17'd41626,17'd41004,17'd39483,17'd38580,17'd38203,17'd13933,17'd14060,17'd6094,17'd6890,17'd7364,17'd7878,17'd9124,17'd9124,17'd9261,17'd9544,17'd6416,17'd7365,17'd3744,17'd229,17'd228,17'd625,17'd626,17'd443,17'd1678,17'd17661,17'd1538,17'd205,17'd1244,17'd41908
},
'{
17'd6420,17'd6420,17'd4243,17'd4243,17'd4892,17'd4892,17'd25384,17'd15746,17'd3252,17'd1831,17'd4247,17'd2595,17'd3905,17'd18,17'd18,17'd3905,17'd17,17'd3905,17'd980,17'd980,17'd27444,17'd4248,17'd3756,17'd3435,17'd2946,17'd19874,17'd1423,17'd1704,17'd1285,17'd2787,17'd2438,17'd14451,17'd14873,17'd16145,17'd2618,17'd41909,17'd14876,17'd4591,17'd41910,17'd18998,17'd38339,17'd15633,17'd41911,17'd41912,17'd41913,17'd27461,17'd17689,17'd17689,17'd17204,17'd7746,17'd18660,17'd20431,17'd14631,17'd39799,17'd39955,17'd41914,17'd41915,17'd40725,17'd41916,17'd41635,17'd41489,17'd41637,17'd40726,17'd41775,17'd39961,17'd41917,17'd41918,17'd41919,17'd41495,17'd41920,17'd41921,17'd17455,17'd41922,17'd41497,17'd9308,17'd9308,17'd9161,17'd24976,17'd41643,17'd8540,17'd6638,17'd6632,17'd41923,17'd41781,17'd41644,17'd41644,17'd41020,17'd41924,17'd41782,17'd40877,17'd41176,17'd41925,17'd41785,17'd41926,17'd41927,17'd41928,17'd40739,17'd41929,17'd41930,17'd6801,17'd39510,17'd41931,17'd41932,17'd24548,17'd10179,17'd8250,17'd25147,17'd11404,17'd8410,17'd8724,17'd16067,17'd9038,17'd9347,17'd13887,17'd17716,17'd10336,17'd16681,17'd8873,17'd15180,17'd11277,17'd21206,17'd14259,17'd26371,17'd29923,17'd29480,17'd31286,17'd35372,17'd28460,17'd28343,17'd26370,17'd24031,17'd21363,17'd23169,17'd22816,17'd22647,17'd11131,17'd22647,17'd11130,17'd11130,17'd10854,17'd11132,17'd10326,17'd17719,17'd21503,17'd9885,17'd12116,17'd9479,17'd9344,17'd15180,17'd12117,17'd9191,17'd9345,17'd16549,17'd15048,17'd9739,17'd11134,17'd11133,17'd19282,17'd10475,17'd10737,17'd13362,17'd18081,17'd33734,17'd30087,17'd41657,17'd41933,17'd33735,17'd33885,17'd33248,17'd35520,17'd29651,17'd34048,17'd41659,17'd18446,17'd41346,17'd41934,17'd41935,17'd41936,17'd41937,17'd41938,17'd41349,17'd41514,17'd40143,17'd40144,17'd41939,17'd41940,17'd41940,17'd41799,17'd41800,17'd35115,17'd41941,17'd41942,17'd41943,17'd41944,17'd41945,17'd41946,17'd41947,17'd41948,17'd41949,17'd41950,17'd41951,17'd41952,17'd41953,17'd41954,17'd41382,17'd41548,17'd41817,17'd41683,17'd41955,17'd41956,17'd41957,17'd41958,17'd41959,17'd41960,17'd41961,17'd41962,17'd41963,17'd41964,17'd41965,17'd41966,17'd41967,17'd41968,17'd41969,17'd41693,17'd41834,17'd41970,17'd41537,17'd41971,17'd41972,17'd41973,17'd41974,17'd41975,17'd41976,17'd41977,17'd41978,17'd41979,17'd41980,17'd41981,17'd41982,17'd41983,17'd41984,17'd41985,17'd41986,17'd41987,17'd40501,17'd33916,17'd41988,17'd35406,17'd38521,17'd36818,17'd41989,17'd41990,17'd41991,17'd41718,17'd41855,17'd41992,17'd41720,17'd41410,17'd41575,17'd41858,17'd41993,17'd41721,17'd41264,17'd41725,17'd41578,17'd41994,17'd41995,17'd41996,17'd41861,17'd41581,17'd41997,17'd41107,17'd41998,17'd41582,17'd41864,17'd41864,17'd32495,17'd32343,17'd25707,17'd27765,17'd27637,17'd30733,17'd29530,17'd32514,17'd32514,17'd30579,17'd31502,17'd23920,17'd31033,17'd23917,17'd23731,17'd23732,17'd24086,17'd23917,17'd28851,17'd25438,17'd28720,17'd25833,17'd27514,17'd41999,17'd31351,17'd39740,17'd34450,17'd40367,17'd32505,17'd33486,17'd29248,17'd32505,17'd29247,17'd28981,17'd26522,17'd28854,17'd33319,17'd31503,17'd32496,17'd38406,17'd42000,17'd42001,17'd32997,17'd22864,17'd42002,17'd42003,17'd21530,17'd33946,17'd31347,17'd42004,17'd25179,17'd32658,17'd28600,17'd27638,17'd30606,17'd26174,17'd26174,17'd27767,17'd27513,17'd26062,17'd33499,17'd26901,17'd26901,17'd30735,17'd28979,17'd29379,17'd39437,17'd35291,17'd34451,17'd34877,17'd41868,17'd42005,17'd40225,17'd41118,17'd41734,17'd32515,17'd42006,17'd36270,17'd32200,17'd42007,17'd42008,17'd42009,17'd42010,17'd42011,17'd35166,17'd29243,17'd42012,17'd24245,17'd24078,17'd25703,17'd27146,17'd27027,17'd34301,17'd27514,17'd24409,17'd42013,17'd28369,17'd42014,17'd42015,17'd42016,17'd42017,17'd42018,17'd42019,17'd42020,17'd42021,17'd42022,17'd41748,17'd42023,17'd41882,17'd42024,17'd23432,17'd22906,17'd42025,17'd36437,17'd42026,17'd42027,17'd39160,17'd18620,17'd42028,17'd42029,17'd37555,17'd41452,17'd40244,17'd22088,17'd37286,17'd42030,17'd28306,17'd28650,17'd9933,17'd29740,17'd8780,17'd6219,17'd5005,17'd4686,17'd42031,17'd4689,17'd4017,17'd41755,17'd39165,17'd4360,17'd5156,17'd5156,17'd4525,17'd4356,17'd4829,17'd4671,17'd39468,17'd34157,17'd42032,17'd42033,17'd41893,17'd12131,17'd41894,17'd41895,17'd33689,17'd42034,17'd42035,17'd42036,17'd42037,17'd41764,17'd42038,17'd42039,17'd42040,17'd37816,17'd41901,17'd42041,17'd2530,17'd42042,17'd3210,17'd41903,17'd41904,17'd4052,17'd3702,17'd42043,17'd5493,17'd41159,17'd10388,17'd38458,17'd41481,17'd38203,17'd13933,17'd14060,17'd6094,17'd6890,17'd7364,17'd7878,17'd9124,17'd7705,17'd9414,17'd9544,17'd6416,17'd4713,17'd3391,17'd1261,17'd1262,17'd1262,17'd2249,17'd623,17'd1380,17'd17661,17'd1538,17'd972,17'd1381,17'd41908
},
'{
17'd6420,17'd6420,17'd4243,17'd27713,17'd4892,17'd4892,17'd25384,17'd4245,17'd2935,17'd1831,17'd4247,17'd2595,17'd3905,17'd18,17'd18,17'd3905,17'd17,17'd16,17'd652,17'd980,17'd27444,17'd4248,17'd3434,17'd3258,17'd2946,17'd19874,17'd1423,17'd1559,17'd1138,17'd2787,17'd2438,17'd22269,17'd22449,17'd16145,17'd2793,17'd41909,17'd14876,17'd4591,17'd41910,17'd18998,17'd38339,17'd15633,17'd41911,17'd42044,17'd19131,17'd19007,17'd17689,17'd17689,17'd17204,17'd19388,17'd19015,17'd39952,17'd42045,17'd42046,17'd42047,17'd42048,17'd42049,17'd42050,17'd42051,17'd42052,17'd41489,17'd41637,17'd40112,17'd42053,17'd42054,17'd42055,17'd42056,17'd41919,17'd42057,17'd42058,17'd34190,17'd42059,17'd41922,17'd41497,17'd9308,17'd9161,17'd25259,17'd25659,17'd8845,17'd8540,17'd6638,17'd42060,17'd42061,17'd41781,17'd41644,17'd42062,17'd40584,17'd41924,17'd42063,17'd40877,17'd42064,17'd41925,17'd42065,17'd42066,17'd42067,17'd41928,17'd42068,17'd42069,17'd42070,17'd42071,17'd42072,17'd42073,17'd42074,17'd24548,17'd10179,17'd8250,17'd25147,17'd11404,17'd8726,17'd8886,17'd15684,17'd9039,17'd9347,17'd24361,17'd37605,17'd10336,17'd16066,17'd10175,17'd15807,17'd11277,17'd21206,17'd14259,17'd26371,17'd28943,17'd29480,17'd29480,17'd28460,17'd30222,17'd28343,17'd27004,17'd24031,17'd21363,17'd23169,17'd22816,17'd22647,17'd10854,17'd22647,17'd11130,17'd11275,17'd11668,17'd21206,17'd11526,17'd26152,17'd21503,17'd9885,17'd12116,17'd9479,17'd9620,17'd9345,17'd12117,17'd9339,17'd9345,17'd16549,17'd11277,17'd9883,17'd10330,17'd19282,17'd19282,17'd10475,17'd10737,17'd11963,17'd18081,17'd33734,17'd29653,17'd41794,17'd33582,17'd33735,17'd33885,17'd33248,17'd32294,17'd29651,17'd12998,17'd12114,17'd42075,17'd41346,17'd33082,17'd42076,17'd42077,17'd41038,17'd41938,17'd41349,17'd41514,17'd42078,17'd40144,17'd42079,17'd42080,17'd41940,17'd42081,17'd42082,17'd42083,17'd42084,17'd42085,17'd42086,17'd42087,17'd42088,17'd42089,17'd42090,17'd42091,17'd42092,17'd42093,17'd42094,17'd42095,17'd41385,17'd41383,17'd42096,17'd42097,17'd42098,17'd42099,17'd42100,17'd42101,17'd42102,17'd42103,17'd42104,17'd42105,17'd42106,17'd42107,17'd42108,17'd42109,17'd42110,17'd42111,17'd42112,17'd42113,17'd42114,17'd42115,17'd42116,17'd42117,17'd41224,17'd42118,17'd42119,17'd42120,17'd42121,17'd42122,17'd42123,17'd42124,17'd42125,17'd42126,17'd42127,17'd42128,17'd42129,17'd42130,17'd42131,17'd42132,17'd39715,17'd42133,17'd42134,17'd42135,17'd37637,17'd35551,17'd37885,17'd42136,17'd37097,17'd42137,17'd42138,17'd42139,17'd42140,17'd42141,17'd42142,17'd41721,17'd41722,17'd41724,17'd42143,17'd41858,17'd42144,17'd41725,17'd41578,17'd41994,17'd41995,17'd42145,17'd41861,17'd42146,17'd41863,17'd41998,17'd41107,17'd41417,17'd41864,17'd41864,17'd32495,17'd32496,17'd25707,17'd25567,17'd28254,17'd30733,17'd29530,17'd32514,17'd39132,17'd38806,17'd31502,17'd24086,17'd23731,17'd23917,17'd23731,17'd28722,17'd23731,17'd23916,17'd25032,17'd25438,17'd28720,17'd26174,17'd26530,17'd28481,17'd42147,17'd39436,17'd36983,17'd40367,17'd32505,17'd33486,17'd29248,17'd29248,17'd28257,17'd28981,17'd26522,17'd26522,17'd32354,17'd31503,17'd32496,17'd42148,17'd42149,17'd36130,17'd34457,17'd42150,17'd42151,17'd42152,17'd42153,17'd22337,17'd32829,17'd42154,17'd25180,17'd32658,17'd25435,17'd28594,17'd28481,17'd26174,17'd26174,17'd27767,17'd27513,17'd28481,17'd33499,17'd26781,17'd26901,17'd29245,17'd38537,17'd29379,17'd31353,17'd41731,17'd34877,17'd40961,17'd42155,17'd42005,17'd40225,17'd40227,17'd41869,17'd42156,17'd41430,17'd31215,17'd32200,17'd42007,17'd42157,17'd42158,17'd42159,17'd42160,17'd42161,17'd25033,17'd24252,17'd23727,17'd26658,17'd25431,17'd27258,17'd27027,17'd42162,17'd27514,17'd24409,17'd42013,17'd25317,17'd36287,17'd42163,17'd42164,17'd42165,17'd42166,17'd42167,17'd42168,17'd42169,17'd40068,17'd42170,17'd42171,17'd42172,17'd42173,17'd42174,17'd35046,17'd42175,17'd42176,17'd42177,17'd42178,17'd39160,17'd18620,17'd42028,17'd42029,17'd37940,17'd41452,17'd40244,17'd22088,17'd37286,17'd37287,17'd28305,17'd28650,17'd9933,17'd29740,17'd7668,17'd6219,17'd5005,17'd4686,17'd5162,17'd5156,17'd4017,17'd41755,17'd39313,17'd4359,17'd4526,17'd4526,17'd4525,17'd39468,17'd5476,17'd42179,17'd4356,17'd42180,17'd42181,17'd42182,17'd42183,17'd42184,17'd41894,17'd42185,17'd42186,17'd42187,17'd42188,17'd41763,17'd42037,17'd42189,17'd42190,17'd42191,17'd42192,17'd39323,17'd41901,17'd42041,17'd2369,17'd42193,17'd42194,17'd3378,17'd42195,17'd41623,17'd3702,17'd41906,17'd42196,17'd41626,17'd41004,17'd38859,17'd38580,17'd38072,17'd13933,17'd14060,17'd6094,17'd6890,17'd7364,17'd7364,17'd9124,17'd9124,17'd9261,17'd8187,17'd6416,17'd4869,17'd3744,17'd229,17'd1401,17'd1262,17'd2249,17'd954,17'd190,17'd3899,17'd1538,17'd204,17'd1381,17'd42197
},
'{
17'd4428,17'd4428,17'd4243,17'd27713,17'd4892,17'd4892,17'd25384,17'd14743,17'd2422,17'd1831,17'd4247,17'd466,17'd3905,17'd18,17'd18,17'd3905,17'd17,17'd18,17'd980,17'd27,17'd4430,17'd4091,17'd3434,17'd3105,17'd2946,17'd19608,17'd1423,17'd1424,17'd1285,17'd2787,17'd994,17'd22269,17'd22449,17'd16145,17'd2793,17'd41909,17'd14876,17'd5232,17'd42198,17'd19745,17'd42199,17'd35774,17'd41911,17'd42200,17'd42201,17'd18774,17'd19128,17'd19128,17'd17317,17'd20024,17'd19015,17'd39952,17'd15015,17'd42202,17'd42203,17'd42204,17'd42049,17'd40725,17'd42205,17'd42206,17'd42207,17'd41637,17'd40112,17'd42053,17'd42054,17'd41917,17'd42208,17'd41919,17'd42057,17'd42209,17'd17816,17'd42210,17'd18785,17'd9706,17'd9308,17'd9306,17'd9305,17'd9160,17'd8689,17'd8375,17'd7914,17'd6480,17'd41923,17'd42211,17'd42212,17'd42062,17'd42213,17'd42214,17'd42063,17'd41023,17'd42215,17'd42216,17'd42217,17'd42218,17'd42219,17'd42220,17'd42221,17'd42222,17'd42223,17'd42224,17'd42225,17'd42226,17'd42227,17'd42228,17'd14136,17'd8250,17'd25147,17'd15429,17'd8726,17'd8569,17'd24999,17'd9039,17'd9347,17'd15180,17'd17716,17'd10336,17'd42229,17'd8874,17'd9345,17'd11671,17'd21206,17'd16325,17'd24856,17'd28943,17'd35372,17'd29480,17'd29923,17'd28343,17'd28343,17'd25672,17'd24705,17'd21363,17'd18327,17'd22816,17'd22647,17'd10854,17'd22647,17'd11130,17'd11668,17'd11399,17'd11132,17'd19280,17'd26152,17'd10024,17'd10992,17'd12116,17'd9479,17'd9620,17'd9345,17'd9344,17'd9339,17'd9345,17'd9619,17'd15048,17'd17839,17'd10479,17'd10991,17'd19282,17'd10475,17'd10853,17'd12114,17'd14002,17'd30685,17'd41794,17'd41657,17'd33736,17'd41795,17'd33885,17'd33248,17'd32294,17'd18192,17'd29491,17'd33410,17'd33097,17'd41346,17'd42230,17'd42231,17'd42232,17'd42233,17'd41938,17'd41516,17'd41197,17'd42234,17'd40144,17'd42235,17'd42236,17'd41940,17'd42081,17'd39525,17'd41043,17'd42237,17'd42238,17'd42239,17'd42240,17'd42241,17'd42242,17'd42243,17'd42244,17'd42245,17'd42246,17'd42247,17'd42248,17'd41681,17'd42249,17'd42250,17'd42251,17'd42252,17'd42253,17'd42254,17'd26161,17'd42255,17'd42256,17'd42257,17'd42258,17'd42259,17'd42260,17'd42261,17'd42262,17'd42263,17'd42264,17'd42265,17'd42266,17'd41825,17'd42267,17'd42268,17'd41373,17'd41071,17'd41546,17'd42269,17'd40642,17'd42270,17'd42271,17'd42272,17'd42273,17'd42274,17'd42275,17'd42276,17'd42277,17'd42278,17'd42279,17'd42280,17'd42281,17'd42282,17'd42283,17'd42284,17'd34994,17'd35684,17'd41988,17'd42285,17'd37884,17'd36964,17'd42137,17'd42286,17'd42287,17'd42288,17'd42289,17'd42290,17'd41576,17'd42291,17'd41993,17'd42292,17'd41724,17'd42293,17'd42294,17'd41578,17'd41994,17'd42295,17'd42145,17'd42296,17'd42146,17'd41863,17'd38665,17'd42297,17'd42298,17'd42299,17'd42300,17'd42301,17'd33477,17'd38538,17'd28597,17'd25029,17'd29688,17'd29376,17'd33800,17'd33651,17'd24421,17'd31502,17'd23732,17'd30879,17'd24415,17'd23917,17'd30879,17'd24415,17'd28851,17'd25031,17'd27511,17'd28723,17'd25949,17'd26530,17'd28481,17'd33155,17'd39436,17'd34877,17'd40367,17'd32505,17'd29248,17'd29248,17'd29248,17'd32507,17'd32192,17'd33319,17'd33319,17'd30279,17'd31353,17'd32496,17'd42302,17'd42303,17'd42304,17'd21693,17'd34280,17'd42151,17'd42305,17'd21701,17'd22510,17'd32666,17'd42004,17'd24897,17'd28721,17'd25566,17'd28594,17'd26062,17'd27515,17'd25833,17'd28481,17'd27513,17'd28481,17'd33815,17'd26782,17'd26781,17'd30735,17'd28727,17'd29379,17'd31353,17'd41731,17'd40961,17'd40961,17'd34275,17'd42005,17'd40225,17'd40227,17'd41869,17'd30148,17'd41430,17'd31215,17'd42306,17'd42307,17'd25712,17'd42009,17'd42010,17'd42308,17'd37922,17'd29242,17'd24901,17'd24740,17'd27370,17'd23908,17'd28978,17'd27258,17'd27371,17'd26530,17'd23554,17'd24410,17'd25317,17'd25319,17'd42161,17'd42309,17'd42310,17'd42311,17'd42312,17'd42313,17'd42314,17'd42315,17'd42170,17'd42171,17'd42316,17'd42317,17'd42318,17'd42319,17'd42175,17'd42320,17'd42177,17'd42321,17'd39307,17'd18260,17'd42028,17'd42029,17'd37940,17'd21772,17'd40846,17'd22250,17'd39771,17'd37287,17'd28305,17'd28650,17'd27815,17'd29740,17'd7499,17'd6390,17'd4842,17'd4841,17'd4848,17'd4526,17'd4357,17'd42322,17'd40395,17'd4833,17'd5000,17'd4526,17'd4525,17'd39468,17'd5476,17'd4670,17'd41455,17'd33839,17'd4360,17'd36022,17'd42183,17'd42184,17'd42323,17'd42185,17'd41465,17'd42324,17'd42325,17'd42326,17'd41152,17'd42189,17'd42190,17'd42327,17'd42328,17'd42329,17'd42330,17'd42331,17'd42332,17'd42333,17'd42194,17'd42334,17'd2723,17'd41904,17'd3702,17'd42043,17'd4055,17'd41159,17'd10790,17'd11867,17'd41481,17'd38072,17'd37959,17'd16492,17'd6094,17'd6890,17'd7364,17'd7364,17'd9124,17'd7705,17'd9544,17'd8187,17'd8186,17'd4713,17'd3391,17'd229,17'd1401,17'd1263,17'd953,17'd953,17'd8812,17'd2779,17'd936,17'd204,17'd1381,17'd42335
},
'{
17'd4428,17'd4428,17'd4243,17'd27713,17'd4892,17'd4892,17'd25384,17'd14743,17'd2422,17'd1688,17'd4247,17'd466,17'd3905,17'd18,17'd18,17'd3905,17'd16,17'd16,17'd28,17'd27,17'd4430,17'd4091,17'd3434,17'd3105,17'd1975,17'd1839,17'd1559,17'd1135,17'd1138,17'd2787,17'd994,17'd42336,17'd22449,17'd16145,17'd2793,17'd41909,17'd14876,17'd5232,17'd42198,17'd17926,17'd42337,17'd15753,17'd42338,17'd42339,17'd41320,17'd18774,17'd19128,17'd19128,17'd17317,17'd42340,17'd14224,17'd17211,17'd15144,17'd42341,17'd42342,17'd42343,17'd41915,17'd42344,17'd42345,17'd42345,17'd42344,17'd42346,17'd40726,17'd39805,17'd42054,17'd42347,17'd42208,17'd41919,17'd42057,17'd42209,17'd17700,17'd42210,17'd42348,17'd9580,17'd42349,17'd9577,17'd9304,17'd8693,17'd5087,17'd8375,17'd6639,17'd42350,17'd6320,17'd42211,17'd42212,17'd42213,17'd42351,17'd42352,17'd42063,17'd41175,17'd42353,17'd42216,17'd42354,17'd42355,17'd42356,17'd42357,17'd42358,17'd42222,17'd42359,17'd42360,17'd42361,17'd42362,17'd42363,17'd42228,17'd14136,17'd8250,17'd25147,17'd15429,17'd8726,17'd8886,17'd15684,17'd9039,17'd9347,17'd24361,17'd37605,17'd10336,17'd42229,17'd9743,17'd9480,17'd11671,17'd21206,17'd16442,17'd24856,17'd28943,17'd35372,17'd29480,17'd29923,17'd28816,17'd28343,17'd25672,17'd24705,17'd21362,17'd18327,17'd22816,17'd22647,17'd10854,17'd22647,17'd11130,17'd11668,17'd11668,17'd12423,17'd19280,17'd19278,17'd13522,17'd16912,17'd12116,17'd9479,17'd9620,17'd9345,17'd9344,17'd9339,17'd9345,17'd9619,17'd11277,17'd11134,17'd11670,17'd11132,17'd19282,17'd10475,17'd10853,17'd11957,17'd14002,17'd30685,17'd42364,17'd41794,17'd33736,17'd41795,17'd33885,17'd42365,17'd35520,17'd18192,17'd12105,17'd16548,17'd33097,17'd41346,17'd28827,17'd42366,17'd42367,17'd41516,17'd42368,17'd41514,17'd40750,17'd42078,17'd40144,17'd42369,17'd42370,17'd41940,17'd41799,17'd32312,17'd42371,17'd42372,17'd42373,17'd42374,17'd42375,17'd42376,17'd42377,17'd42378,17'd42379,17'd42380,17'd42381,17'd42382,17'd42383,17'd41681,17'd42249,17'd42384,17'd42385,17'd42386,17'd42387,17'd42388,17'd42389,17'd42390,17'd42391,17'd42392,17'd42393,17'd42394,17'd42395,17'd42396,17'd42397,17'd42398,17'd42399,17'd42400,17'd42401,17'd42402,17'd42403,17'd42404,17'd42405,17'd41236,17'd42406,17'd42407,17'd42408,17'd42409,17'd42410,17'd42411,17'd42412,17'd42413,17'd42414,17'd42415,17'd42416,17'd42417,17'd42418,17'd42419,17'd42420,17'd42421,17'd42422,17'd42423,17'd42424,17'd35273,17'd35406,17'd42425,17'd37885,17'd37226,17'd41568,17'd42426,17'd42427,17'd42428,17'd42429,17'd42430,17'd42431,17'd42432,17'd42143,17'd42433,17'd41993,17'd42293,17'd42434,17'd41994,17'd41994,17'd42295,17'd42435,17'd42296,17'd42146,17'd41863,17'd38665,17'd42297,17'd42436,17'd42299,17'd42300,17'd42301,17'd33477,17'd38538,17'd25709,17'd24896,17'd35159,17'd29099,17'd33651,17'd32504,17'd40960,17'd31502,17'd30275,17'd30879,17'd24415,17'd23917,17'd24090,17'd24252,17'd24895,17'd25179,17'd28850,17'd25566,17'd27766,17'd26062,17'd26062,17'd42437,17'd39276,17'd34451,17'd39743,17'd32505,17'd29248,17'd29248,17'd29248,17'd32507,17'd32192,17'd33319,17'd33001,17'd30279,17'd31352,17'd32496,17'd42438,17'd42303,17'd35856,17'd42150,17'd34109,17'd42439,17'd42440,17'd42441,17'd32010,17'd33480,17'd42442,17'd24744,17'd25435,17'd25566,17'd26064,17'd26062,17'd26903,17'd25833,17'd28481,17'd27513,17'd28481,17'd33815,17'd26782,17'd26781,17'd29245,17'd28980,17'd29379,17'd31353,17'd41731,17'd40961,17'd38975,17'd37658,17'd42443,17'd41117,17'd35306,17'd42444,17'd30148,17'd41430,17'd36410,17'd42445,17'd32695,17'd42446,17'd42447,17'd41738,17'd42448,17'd42163,17'd42449,17'd23731,17'd23914,17'd24738,17'd24584,17'd28724,17'd27258,17'd26782,17'd33815,17'd24242,17'd24410,17'd25317,17'd30432,17'd39134,17'd42450,17'd24256,17'd42451,17'd42452,17'd42453,17'd42314,17'd42454,17'd42455,17'd42456,17'd42457,17'd42458,17'd39458,17'd19961,17'd42459,17'd42320,17'd42177,17'd42460,17'd39307,17'd18260,17'd19088,17'd22943,17'd37940,17'd21772,17'd41452,17'd22250,17'd39771,17'd42461,17'd28305,17'd28650,17'd27815,17'd29740,17'd7499,17'd27935,17'd4841,17'd4683,17'd5157,17'd4526,17'd42462,17'd42463,17'd42464,17'd4358,17'd5000,17'd4526,17'd4525,17'd39468,17'd5476,17'd4829,17'd4185,17'd4017,17'd4361,17'd42179,17'd42183,17'd42465,17'd42323,17'd42466,17'd42467,17'd42468,17'd42469,17'd41763,17'd42470,17'd42471,17'd42190,17'd42327,17'd42472,17'd42473,17'd42330,17'd42474,17'd42475,17'd42476,17'd42477,17'd42478,17'd42479,17'd41904,17'd3702,17'd41906,17'd42196,17'd41626,17'd40716,17'd38859,17'd38580,17'd38072,17'd38459,17'd37959,17'd6094,17'd6890,17'd7364,17'd7364,17'd9124,17'd9124,17'd7705,17'd8187,17'd8186,17'd4869,17'd3744,17'd3895,17'd1401,17'd230,17'd1263,17'd953,17'd8812,17'd42480,17'd42481,17'd1537,17'd202,17'd42482
},
'{
17'd4428,17'd4428,17'd3902,17'd4891,17'd4892,17'd4892,17'd6420,17'd14743,17'd3252,17'd1831,17'd4247,17'd466,17'd3905,17'd18,17'd18,17'd3905,17'd16,17'd18,17'd980,17'd980,17'd4430,17'd4091,17'd3104,17'd2601,17'd1974,17'd1839,17'd1559,17'd1424,17'd17079,17'd2788,17'd995,17'd14451,17'd22449,17'd14604,17'd40259,17'd41909,17'd42483,17'd5232,17'd25507,17'd18047,17'd15503,17'd15753,17'd42338,17'd42484,17'd42485,17'd17689,17'd19382,17'd19006,17'd19621,17'd19261,17'd18537,17'd41486,17'd42486,17'd42202,17'd38470,17'd42487,17'd42488,17'd42489,17'd42490,17'd42491,17'd42207,17'd42492,17'd39958,17'd39804,17'd42493,17'd42347,17'd42494,17'd42495,17'd42496,17'd41017,17'd17700,17'd42497,17'd20436,17'd10121,17'd42498,17'd9577,17'd9576,17'd42499,17'd42500,17'd8375,17'd6639,17'd6480,17'd42501,17'd6323,17'd42212,17'd42502,17'd42503,17'd42504,17'd42505,17'd42506,17'd42507,17'd42508,17'd42509,17'd42510,17'd42511,17'd42512,17'd42513,17'd42514,17'd42515,17'd42516,17'd42517,17'd42518,17'd42519,17'd42520,17'd7785,17'd9484,17'd8413,17'd15429,17'd8725,17'd9040,17'd8873,17'd10174,17'd8874,17'd10174,17'd16795,17'd10175,17'd17600,17'd8874,17'd15187,17'd9883,17'd11668,17'd22992,17'd24856,17'd28104,17'd28818,17'd28460,17'd28343,17'd28343,17'd26872,17'd24856,17'd24992,17'd22472,17'd21985,17'd22816,17'd11130,17'd11130,17'd11130,17'd11130,17'd11668,17'd11668,17'd12423,17'd19280,17'd17847,17'd10024,17'd11136,17'd12116,17'd9479,17'd9620,17'd15187,17'd9344,17'd9339,17'd9345,17'd15048,17'd14928,17'd11134,17'd12863,17'd19532,17'd10476,17'd10474,17'd10737,17'd12114,17'd41793,17'd42364,17'd30236,17'd41933,17'd41933,17'd33735,17'd33885,17'd33248,17'd30086,17'd18192,17'd34391,17'd38752,17'd33097,17'd41511,17'd28827,17'd42521,17'd41661,17'd41350,17'd42522,17'd41516,17'd42523,17'd40143,17'd42524,17'd42525,17'd42526,17'd42527,17'd42528,17'd42529,17'd42530,17'd42531,17'd42532,17'd42533,17'd42534,17'd42535,17'd42536,17'd42537,17'd42538,17'd42539,17'd42540,17'd42541,17'd42542,17'd42543,17'd42544,17'd42545,17'd40633,17'd42546,17'd42547,17'd42548,17'd42549,17'd42550,17'd42551,17'd42552,17'd42553,17'd42554,17'd42555,17'd42556,17'd42557,17'd42558,17'd42559,17'd42560,17'd42561,17'd42562,17'd42563,17'd41972,17'd41698,17'd42098,17'd42564,17'd42565,17'd42566,17'd42567,17'd42568,17'd42569,17'd42570,17'd42571,17'd42572,17'd42573,17'd42574,17'd42575,17'd42576,17'd42577,17'd42578,17'd40026,17'd42579,17'd42580,17'd42581,17'd35684,17'd38392,17'd42582,17'd40350,17'd36820,17'd42583,17'd42584,17'd42585,17'd42586,17'd42587,17'd42588,17'd38963,17'd42589,17'd42292,17'd42590,17'd42143,17'd42591,17'd42592,17'd42593,17'd42594,17'd42595,17'd42596,17'd41861,17'd42146,17'd40822,17'd38536,17'd42297,17'd42436,17'd42597,17'd42300,17'd42598,17'd33309,17'd28483,17'd27512,17'd24896,17'd23916,17'd29099,17'd38979,17'd29374,17'd34112,17'd30127,17'd34137,17'd28722,17'd24415,17'd23917,17'd24090,17'd24417,17'd25030,17'd25179,17'd29101,17'd28720,17'd25708,17'd27767,17'd25708,17'd42599,17'd42600,17'd35291,17'd32831,17'd33165,17'd29248,17'd29248,17'd33486,17'd29248,17'd32192,17'd40681,17'd29977,17'd32356,17'd28979,17'd32343,17'd42438,17'd42601,17'd34757,17'd22337,17'd35155,17'd21530,17'd42602,17'd42603,17'd34457,17'd33480,17'd42604,17'd23561,17'd28721,17'd32658,17'd27766,17'd28482,17'd26903,17'd25833,17'd28481,17'd26064,17'd28481,17'd28009,17'd26782,17'd26901,17'd28486,17'd29245,17'd29246,17'd39437,17'd34451,17'd38975,17'd38805,17'd34274,17'd34104,17'd42605,17'd42606,17'd27644,17'd37406,17'd31361,17'd31215,17'd42445,17'd42157,17'd42607,17'd42608,17'd42609,17'd42448,17'd42610,17'd42611,17'd23564,17'd24416,17'd23726,17'd24078,17'd28252,17'd27258,17'd25311,17'd24735,17'd27766,17'd28130,17'd23725,17'd30432,17'd30883,17'd42612,17'd42613,17'd42614,17'd32698,17'd42615,17'd42616,17'd42617,17'd42618,17'd42456,17'd42619,17'd42620,17'd42621,17'd20966,17'd42622,17'd42623,17'd16464,17'd42624,17'd42625,17'd20384,17'd42028,17'd36029,17'd37940,17'd21772,17'd42626,17'd39162,17'd39771,17'd37429,17'd28534,17'd10897,17'd27815,17'd29740,17'd9091,17'd28185,17'd5328,17'd42627,17'd4847,17'd5154,17'd42462,17'd42628,17'd42629,17'd33839,17'd4525,17'd4526,17'd4525,17'd4358,17'd42630,17'd4828,17'd42631,17'd4016,17'd4365,17'd4987,17'd42632,17'd42465,17'd42633,17'd42634,17'd42635,17'd42636,17'd41469,17'd42637,17'd42638,17'd42639,17'd42640,17'd42641,17'd42642,17'd42643,17'd42644,17'd2715,17'd42645,17'd42476,17'd42477,17'd42646,17'd2535,17'd42647,17'd41624,17'd9530,17'd4055,17'd41003,17'd11188,17'd39033,17'd38580,17'd38072,17'd16492,17'd37959,17'd6258,17'd6890,17'd7878,17'd7364,17'd7538,17'd9261,17'd9544,17'd8187,17'd8186,17'd4869,17'd3744,17'd3895,17'd1261,17'd1262,17'd1962,17'd1962,17'd1667,17'd606,17'd1537,17'd42648,17'd1527,17'd195
},
'{
17'd4428,17'd4428,17'd3902,17'd4891,17'd4892,17'd4892,17'd25384,17'd14743,17'd3252,17'd1831,17'd4247,17'd466,17'd3905,17'd18,17'd18,17'd3905,17'd16,17'd18,17'd980,17'd980,17'd4430,17'd4091,17'd3104,17'd2264,17'd1974,17'd1839,17'd1559,17'd1135,17'd992,17'd18275,17'd995,17'd14451,17'd22449,17'd14604,17'd40259,17'd29307,17'd22274,17'd42649,17'd42650,17'd18999,17'd36049,17'd35349,17'd42651,17'd42652,17'd19007,17'd17689,17'd19382,17'd19006,17'd19621,17'd21346,17'd20588,17'd41486,17'd42486,17'd42202,17'd38470,17'd42487,17'd42653,17'd41489,17'd42206,17'd42654,17'd42344,17'd42655,17'd41172,17'd39803,17'd39639,17'd42347,17'd42494,17'd42656,17'd42657,17'd42658,17'd42659,17'd42660,17'd9845,17'd10121,17'd42661,17'd9577,17'd9576,17'd5252,17'd5087,17'd8376,17'd6639,17'd42350,17'd42662,17'd42663,17'd42664,17'd42502,17'd42503,17'd42665,17'd42507,17'd42666,17'd42667,17'd42668,17'd42669,17'd41179,17'd42670,17'd42671,17'd39353,17'd42514,17'd42515,17'd42672,17'd42517,17'd42518,17'd42673,17'd42520,17'd7785,17'd9484,17'd17481,17'd15429,17'd8725,17'd9040,17'd8873,17'd10174,17'd8874,17'd10174,17'd16795,17'd10175,17'd17600,17'd9743,17'd9479,17'd9883,17'd11668,17'd22992,17'd24856,17'd30222,17'd35372,17'd28460,17'd28816,17'd28816,17'd26872,17'd24856,17'd24209,17'd22472,17'd21985,17'd22816,17'd11130,17'd11130,17'd11130,17'd11130,17'd11668,17'd11668,17'd12423,17'd13647,17'd42674,17'd13522,17'd20607,17'd9741,17'd9479,17'd9480,17'd15187,17'd9344,17'd9339,17'd9480,17'd12116,17'd11671,17'd10330,17'd11670,17'd19532,17'd11132,17'd10473,17'd10853,17'd12114,17'd14002,17'd42675,17'd42676,17'd30236,17'd41933,17'd33735,17'd33885,17'd31449,17'd30086,17'd18192,17'd41659,17'd16548,17'd42677,17'd24708,17'd25278,17'd42678,17'd41661,17'd41350,17'd42522,17'd41516,17'd42523,17'd42078,17'd42679,17'd42680,17'd42526,17'd42527,17'd42681,17'd42682,17'd42530,17'd42683,17'd42684,17'd42685,17'd42686,17'd42687,17'd42688,17'd42378,17'd42689,17'd42690,17'd42691,17'd42692,17'd42693,17'd42694,17'd42695,17'd42696,17'd41368,17'd42697,17'd42698,17'd25935,17'd42699,17'd42700,17'd42701,17'd42702,17'd42703,17'd42703,17'd42704,17'd42705,17'd42706,17'd42707,17'd42708,17'd42709,17'd42710,17'd42711,17'd42712,17'd42713,17'd40639,17'd41680,17'd42714,17'd42715,17'd42716,17'd42717,17'd42718,17'd42719,17'd42720,17'd42721,17'd42722,17'd42723,17'd42724,17'd42725,17'd41395,17'd42726,17'd38930,17'd42727,17'd42728,17'd42729,17'd40348,17'd34076,17'd35406,17'd42730,17'd40350,17'd37226,17'd42583,17'd41569,17'd42731,17'd42732,17'd42733,17'd42734,17'd41260,17'd42292,17'd42433,17'd42735,17'd42736,17'd42591,17'd42592,17'd42593,17'd42594,17'd42595,17'd42737,17'd42738,17'd41862,17'd42739,17'd41107,17'd42740,17'd42741,17'd42742,17'd42743,17'd42598,17'd33310,17'd32996,17'd27512,17'd24417,17'd34467,17'd34137,17'd42744,17'd23923,17'd31190,17'd29099,17'd28976,17'd28722,17'd34467,17'd24249,17'd24415,17'd24417,17'd28254,17'd25320,17'd28850,17'd28720,17'd25708,17'd27767,17'd25708,17'd41270,17'd42600,17'd35291,17'd32831,17'd33165,17'd29248,17'd33486,17'd33486,17'd29248,17'd32192,17'd29977,17'd27642,17'd29379,17'd26901,17'd32185,17'd42438,17'd42745,17'd42746,17'd22511,17'd35155,17'd42440,17'd42747,17'd34616,17'd32997,17'd31834,17'd42748,17'd29240,17'd42749,17'd32658,17'd27766,17'd28482,17'd27259,17'd27515,17'd28481,17'd26064,17'd28481,17'd28009,17'd26782,17'd26901,17'd28979,17'd29246,17'd29245,17'd37908,17'd34877,17'd38975,17'd41108,17'd33475,17'd42750,17'd27886,17'd42606,17'd27644,17'd37406,17'd30149,17'd36410,17'd42751,17'd42157,17'd42752,17'd42753,17'd42754,17'd42755,17'd42756,17'd25181,17'd25033,17'd24252,17'd23726,17'd24078,17'd25833,17'd28978,17'd25702,17'd24735,17'd27766,17'd28594,17'd24585,17'd25320,17'd25439,17'd34123,17'd42757,17'd42758,17'd42759,17'd42760,17'd42761,17'd42762,17'd42763,17'd42764,17'd41290,17'd39151,17'd42765,17'd42766,17'd38693,17'd42767,17'd42768,17'd42769,17'd42770,17'd20384,17'd19222,17'd36734,17'd17654,17'd21772,17'd42626,17'd22250,17'd37286,17'd37557,17'd30488,17'd27932,17'd10515,17'd7499,17'd6390,17'd30638,17'd5327,17'd42771,17'd4847,17'd34657,17'd42462,17'd40395,17'd39773,17'd33839,17'd4525,17'd4526,17'd4525,17'd34157,17'd42772,17'd4828,17'd42628,17'd4185,17'd4363,17'd42773,17'd42632,17'd42774,17'd42633,17'd42634,17'd42634,17'd42775,17'd42776,17'd42777,17'd3529,17'd42639,17'd42778,17'd42779,17'd42642,17'd42643,17'd42644,17'd39625,17'd42780,17'd42781,17'd42782,17'd42783,17'd42784,17'd2889,17'd3702,17'd41001,17'd42196,17'd41003,17'd11188,17'd39033,17'd38580,17'd38072,17'd16492,17'd16492,17'd6258,17'd6890,17'd7364,17'd7364,17'd7538,17'd9124,17'd7705,17'd6416,17'd8186,17'd4869,17'd3744,17'd5193,17'd229,17'd1401,17'd1262,17'd1962,17'd1667,17'd1112,17'd775,17'd42785,17'd421,17'd42786
},
'{
17'd3903,17'd3903,17'd3902,17'd4891,17'd4243,17'd4892,17'd25384,17'd14743,17'd3252,17'd2594,17'd2595,17'd466,17'd3905,17'd18,17'd18,17'd3905,17'd18,17'd18,17'd980,17'd980,17'd4430,17'd4091,17'd3104,17'd2264,17'd1974,17'd1839,17'd1559,17'd1138,17'd17079,17'd18275,17'd995,17'd14451,17'd22449,17'd14604,17'd40259,17'd29307,17'd3928,17'd5531,17'd42650,17'd18047,17'd42787,17'd35349,17'd42651,17'd42652,17'd19007,17'd17941,17'd19382,17'd19006,17'd39797,17'd19894,17'd18537,17'd16990,17'd42788,17'd42202,17'd42494,17'd42789,17'd40112,17'd41489,17'd42345,17'd42654,17'd42207,17'd42492,17'd39958,17'd39803,17'd39639,17'd39340,17'd42790,17'd42656,17'd42657,17'd42791,17'd42792,17'd19266,17'd9988,17'd42793,17'd42661,17'd42794,17'd9576,17'd5252,17'd5251,17'd42795,17'd42796,17'd42350,17'd42662,17'd42797,17'd42798,17'd42799,17'd42800,17'd42665,17'd42507,17'd42666,17'd42667,17'd42668,17'd42801,17'd41335,17'd42802,17'd42671,17'd39353,17'd42803,17'd42804,17'd42805,17'd42806,17'd42807,17'd38234,17'd42808,17'd42809,17'd13888,17'd12865,17'd15429,17'd8724,17'd9040,17'd9038,17'd12117,17'd8874,17'd8874,17'd16795,17'd10175,17'd17600,17'd9347,17'd16554,17'd9883,17'd11668,17'd22992,17'd24856,17'd27857,17'd28345,17'd28818,17'd28816,17'd26370,17'd26370,17'd24537,17'd24209,17'd22472,17'd21985,17'd19533,17'd11130,17'd11130,17'd11130,17'd11130,17'd11668,17'd11668,17'd12423,17'd19280,17'd17847,17'd10024,17'd11136,17'd9741,17'd9479,17'd9480,17'd15187,17'd9345,17'd9346,17'd9345,17'd9619,17'd11277,17'd11134,17'd11670,17'd24996,17'd11132,17'd10473,17'd10853,17'd12114,17'd41793,17'd42364,17'd30236,17'd33582,17'd33582,17'd33735,17'd33885,17'd31449,17'd30086,17'd18192,17'd41659,17'd16548,17'd42810,17'd28827,17'd10734,17'd42811,17'd42812,17'd41938,17'd40891,17'd40891,17'd42813,17'd42234,17'd42814,17'd42815,17'd42236,17'd42527,17'd42816,17'd42682,17'd42817,17'd42818,17'd38121,17'd42819,17'd42820,17'd42821,17'd42822,17'd42823,17'd42824,17'd42825,17'd42826,17'd42827,17'd41238,17'd41370,17'd42543,17'd42828,17'd42829,17'd42830,17'd42831,17'd42832,17'd42833,17'd42834,17'd42397,17'd42835,17'd42835,17'd42836,17'd42837,17'd42838,17'd42839,17'd42840,17'd42841,17'd42842,17'd42843,17'd42844,17'd42845,17'd42846,17'd42847,17'd42848,17'd41541,17'd42849,17'd42850,17'd42851,17'd42852,17'd42853,17'd42854,17'd42855,17'd42856,17'd42857,17'd42858,17'd42859,17'd42860,17'd42726,17'd42861,17'd42862,17'd42863,17'd42864,17'd42865,17'd42866,17'd42867,17'd35551,17'd40350,17'd36385,17'd42868,17'd42869,17'd42870,17'd41570,17'd42871,17'd42872,17'd42873,17'd42874,17'd42875,17'd42876,17'd42874,17'd40812,17'd42877,17'd42594,17'd42878,17'd42879,17'd42880,17'd42881,17'd41862,17'd42739,17'd42882,17'd42600,17'd42883,17'd42884,17'd42885,17'd40959,17'd33310,17'd33643,17'd28254,17'd24744,17'd34467,17'd23564,17'd29830,17'd29099,17'd33794,17'd29376,17'd23385,17'd24086,17'd30431,17'd30431,17'd24415,17'd24896,17'd27512,17'd25438,17'd28369,17'd28600,17'd27766,17'd27767,17'd25833,17'd42886,17'd40824,17'd36541,17'd33485,17'd32355,17'd32505,17'd29248,17'd33486,17'd29248,17'd33654,17'd29977,17'd39437,17'd28727,17'd26781,17'd32496,17'd42438,17'd39282,17'd42887,17'd22511,17'd35710,17'd42888,17'd42747,17'd40522,17'd31192,17'd22860,17'd33651,17'd34622,17'd42749,17'd32658,17'd26174,17'd33815,17'd27371,17'd27515,17'd28481,17'd28481,17'd27639,17'd28009,17'd26782,17'd26901,17'd28486,17'd29245,17'd29245,17'd37908,17'd34274,17'd42889,17'd40958,17'd33475,17'd42890,17'd42891,17'd42606,17'd27644,17'd37406,17'd30149,17'd42892,17'd42893,17'd42752,17'd42894,17'd42895,17'd42896,17'd42897,17'd24746,17'd36414,17'd29242,17'd24090,17'd24893,17'd23724,17'd27766,17'd28252,17'd25702,17'd24582,17'd27766,17'd28130,17'd23725,17'd23558,17'd24088,17'd32841,17'd24747,17'd38686,17'd42898,17'd42899,17'd42900,17'd42901,17'd42902,17'd42903,17'd42023,17'd18585,17'd42904,17'd42905,17'd42906,17'd21589,17'd42907,17'd42908,17'd38699,17'd38566,17'd18970,17'd22943,17'd17534,17'd21772,17'd42909,17'd41140,17'd37428,17'd36030,17'd29161,17'd11181,17'd10514,17'd7499,17'd6554,17'd25627,17'd42910,17'd4688,17'd4684,17'd41891,17'd42462,17'd5476,17'd42629,17'd39468,17'd4525,17'd4526,17'd5155,17'd34157,17'd42772,17'd4828,17'd42628,17'd42630,17'd33204,17'd4985,17'd42911,17'd33527,17'd42633,17'd42634,17'd42634,17'd42912,17'd42913,17'd42777,17'd42914,17'd42915,17'd42916,17'd42917,17'd42918,17'd42919,17'd42644,17'd2715,17'd42920,17'd42781,17'd42921,17'd42783,17'd42784,17'd2723,17'd41624,17'd9530,17'd4055,17'd41003,17'd11188,17'd39033,17'd38580,17'd38072,17'd16492,17'd16492,17'd6417,17'd7364,17'd7364,17'd7364,17'd9124,17'd7705,17'd8187,17'd6416,17'd7365,17'd4869,17'd3744,17'd3895,17'd1261,17'd1401,17'd1262,17'd1680,17'd4084,17'd425,17'd204,17'd42922,17'd419,17'd42923
},
'{
17'd3903,17'd3903,17'd3902,17'd4891,17'd4243,17'd4892,17'd25384,17'd14743,17'd3252,17'd1831,17'd4247,17'd466,17'd3905,17'd18,17'd18,17'd3905,17'd19,17'd18,17'd980,17'd980,17'd4430,17'd4091,17'd3104,17'd2264,17'd1974,17'd1282,17'd1135,17'd1137,17'd992,17'd18275,17'd995,17'd14451,17'd14873,17'd14604,17'd40259,17'd29307,17'd3928,17'd5531,17'd42650,17'd18999,17'd42924,17'd42925,17'd42926,17'd42927,17'd19007,17'd17941,17'd19006,17'd19006,17'd39797,17'd21039,17'd40260,17'd16662,17'd42928,17'd42929,17'd42494,17'd42789,17'd40726,17'd41774,17'd42345,17'd42654,17'd42207,17'd42655,17'd41172,17'd42930,17'd42931,17'd39340,17'd42790,17'd42656,17'd42657,17'd42791,17'd42792,17'd31748,17'd9845,17'd9843,17'd9987,17'd9986,17'd9009,17'd5252,17'd5087,17'd42795,17'd42932,17'd42350,17'd6320,17'd42933,17'd42934,17'd42799,17'd42800,17'd42935,17'd42936,17'd42937,17'd42938,17'd42939,17'd42940,17'd42941,17'd42802,17'd42942,17'd39353,17'd42943,17'd42944,17'd42945,17'd38362,17'd42946,17'd38234,17'd42808,17'd42947,17'd13888,17'd12865,17'd15429,17'd8724,17'd16067,17'd9038,17'd13887,17'd8874,17'd8874,17'd16795,17'd10175,17'd17600,17'd9743,17'd9479,17'd9883,17'd11668,17'd22992,17'd25927,17'd28460,17'd28571,17'd28818,17'd28816,17'd26370,17'd26370,17'd24537,17'd24209,17'd22472,17'd21985,17'd19533,17'd11130,17'd11275,17'd11130,17'd11275,17'd11668,17'd11668,17'd12423,17'd13647,17'd42674,17'd13522,17'd20607,17'd9885,17'd9479,17'd9479,17'd15569,17'd9345,17'd9344,17'd9480,17'd12116,17'd11671,17'd10330,17'd11670,17'd19532,17'd11132,17'd27743,17'd20910,17'd12114,17'd14002,17'd42675,17'd30984,17'd31450,17'd33582,17'd33735,17'd33416,17'd29936,17'd29489,17'd42948,17'd41659,17'd21822,17'd32137,17'd10852,17'd24702,17'd42949,17'd42950,17'd41938,17'd40891,17'd40891,17'd42813,17'd42951,17'd42952,17'd42815,17'd42236,17'd41353,17'd42953,17'd42954,17'd42955,17'd42956,17'd42957,17'd42958,17'd42959,17'd42960,17'd42961,17'd42962,17'd42963,17'd42964,17'd42965,17'd42966,17'd42967,17'd41222,17'd42968,17'd42969,17'd42970,17'd42971,17'd42972,17'd42973,17'd42974,17'd42975,17'd42976,17'd42977,17'd42978,17'd42979,17'd42980,17'd42981,17'd42982,17'd42983,17'd42984,17'd42985,17'd42986,17'd42987,17'd42988,17'd42989,17'd42990,17'd42991,17'd41541,17'd41679,17'd42992,17'd42409,17'd42993,17'd42994,17'd40010,17'd42995,17'd42996,17'd42997,17'd42998,17'd42859,17'd42999,17'd43000,17'd42861,17'd43001,17'd43002,17'd43003,17'd33452,17'd35973,17'd43004,17'd35551,17'd36385,17'd39262,17'd43005,17'd43006,17'd43007,17'd43008,17'd43009,17'd43010,17'd41857,17'd43011,17'd43012,17'd43013,17'd42875,17'd40951,17'd43014,17'd42594,17'd42878,17'd42879,17'd43015,17'd42881,17'd41862,17'd42739,17'd42882,17'd41582,17'd43016,17'd43017,17'd43018,17'd43019,17'd43020,17'd42749,17'd25029,17'd24895,17'd34467,17'd30275,17'd28976,17'd23734,17'd33950,17'd29376,17'd23385,17'd24086,17'd30431,17'd30431,17'd34467,17'd28596,17'd25568,17'd27511,17'd28369,17'd28600,17'd28602,17'd27767,17'd25707,17'd43021,17'd40824,17'd36541,17'd33485,17'd32355,17'd29248,17'd33486,17'd33656,17'd29248,17'd33654,17'd27642,17'd31353,17'd29245,17'd33963,17'd27146,17'd38282,17'd31194,17'd32348,17'd22337,17'd42603,17'd21532,17'd42747,17'd40522,17'd21846,17'd33311,17'd38979,17'd34622,17'd43022,17'd28253,17'd26174,17'd35578,17'd27371,17'd26903,17'd28481,17'd28481,17'd27639,17'd33815,17'd26782,17'd26781,17'd28726,17'd29246,17'd29245,17'd38025,17'd40961,17'd41108,17'd41582,17'd39436,17'd42750,17'd27886,17'd42606,17'd27644,17'd37406,17'd43023,17'd36410,17'd42751,17'd42446,17'd34296,17'd43024,17'd43025,17'd43026,17'd35165,17'd43027,17'd42611,17'd28975,17'd24893,17'd23724,17'd28723,17'd25707,17'd25703,17'd27514,17'd32364,17'd27638,17'd24585,17'd23558,17'd30731,17'd32201,17'd42016,17'd43028,17'd43029,17'd43030,17'd43031,17'd43032,17'd43033,17'd43034,17'd43035,17'd34144,17'd43036,17'd43037,17'd43038,17'd43039,17'd43040,17'd43041,17'd43042,17'd38566,17'd19087,17'd22942,17'd17534,17'd21772,17'd42909,17'd43043,17'd38845,17'd39312,17'd43044,17'd11709,17'd30332,17'd7499,17'd31717,17'd5004,17'd42910,17'd43045,17'd5156,17'd41891,17'd4018,17'd42772,17'd39469,17'd39468,17'd4525,17'd4526,17'd4526,17'd33992,17'd4185,17'd4828,17'd43046,17'd42630,17'd39610,17'd36303,17'd43047,17'd43048,17'd43049,17'd43050,17'd3526,17'd43051,17'd43052,17'd42777,17'd42914,17'd42915,17'd43053,17'd43054,17'd43055,17'd42919,17'd42644,17'd39625,17'd38328,17'd43056,17'd43057,17'd43058,17'd42784,17'd3208,17'd4392,17'd41001,17'd41907,17'd18629,17'd11587,17'd39033,17'd38580,17'd38072,17'd16492,17'd16492,17'd6417,17'd6418,17'd7364,17'd7364,17'd9124,17'd9124,17'd7537,17'd6416,17'd7365,17'd5194,17'd3744,17'd5193,17'd229,17'd1401,17'd1680,17'd2417,17'd4084,17'd1394,17'd1100,17'd43059,17'd600,17'd42923
},
'{
17'd3903,17'd3903,17'd3902,17'd4891,17'd3902,17'd4243,17'd25384,17'd14743,17'd3252,17'd4247,17'd466,17'd466,17'd3905,17'd19,17'd18,17'd3905,17'd19,17'd18,17'd980,17'd980,17'd4430,17'd4091,17'd3104,17'd2264,17'd1974,17'd16966,17'd1559,17'd1138,17'd17079,17'd18275,17'd832,17'd22269,17'd14873,17'd2615,17'd43060,17'd29307,17'd3928,17'd5531,17'd14995,17'd31264,17'd32735,17'd42925,17'd42926,17'd43061,17'd17689,17'd17204,17'd19006,17'd19006,17'd43062,17'd43063,17'd43064,17'd14773,17'd43065,17'd38734,17'd42790,17'd42789,17'd40726,17'd41916,17'd42345,17'd42654,17'd41489,17'd42492,17'd43066,17'd42930,17'd42931,17'd41773,17'd41487,17'd42656,17'd43067,17'd42791,17'd42792,17'd19266,17'd9988,17'd42793,17'd42661,17'd6466,17'd6305,17'd43068,17'd5086,17'd43069,17'd43070,17'd43071,17'd6312,17'd42933,17'd42934,17'd43072,17'd43073,17'd42935,17'd42936,17'd43074,17'd42938,17'd43075,17'd40588,17'd43076,17'd43077,17'd42942,17'd39353,17'd7278,17'd43078,17'd43079,17'd38233,17'd43080,17'd43081,17'd43082,17'd42947,17'd13888,17'd9196,17'd8573,17'd8728,17'd16067,17'd8874,17'd13887,17'd8874,17'd9038,17'd14811,17'd9042,17'd17600,17'd9339,17'd10742,17'd26152,17'd11275,17'd22992,17'd25927,17'd27857,17'd28462,17'd28818,17'd28816,17'd27004,17'd25927,17'd24707,17'd24209,17'd22472,17'd21985,17'd19533,17'd11275,17'd11275,17'd11275,17'd11275,17'd37196,17'd11668,17'd12584,17'd11400,17'd17847,17'd10024,17'd11136,17'd9885,17'd9479,17'd9479,17'd15569,17'd9345,17'd9341,17'd10743,17'd12116,17'd14928,17'd10479,17'd12863,17'd19532,17'd11132,17'd10473,17'd20910,17'd18447,17'd41793,17'd42676,17'd31450,17'd33736,17'd33582,17'd33735,17'd41795,17'd30085,17'd33099,17'd43083,17'd41659,17'd21822,17'd23336,17'd24702,17'd16907,17'd43084,17'd43085,17'd41938,17'd40891,17'd40891,17'd43086,17'd43087,17'd43088,17'd43089,17'd42236,17'd41353,17'd42953,17'd43090,17'd42955,17'd43091,17'd36804,17'd43092,17'd43093,17'd43094,17'd43095,17'd43096,17'd42091,17'd43097,17'd43098,17'd43099,17'd41058,17'd41682,17'd43100,17'd43101,17'd43102,17'd43103,17'd43104,17'd43105,17'd43106,17'd43107,17'd43108,17'd43109,17'd43110,17'd43111,17'd43112,17'd43113,17'd43114,17'd43115,17'd43116,17'd43117,17'd43118,17'd43119,17'd43120,17'd43121,17'd43122,17'd43123,17'd42565,17'd43124,17'd40642,17'd40644,17'd43125,17'd43126,17'd40009,17'd43127,17'd43128,17'd43129,17'd42998,17'd43130,17'd43131,17'd43000,17'd43132,17'd43133,17'd43134,17'd43135,17'd43136,17'd35973,17'd41567,17'd35971,17'd35972,17'd39887,17'd43137,17'd42869,17'd43138,17'd43139,17'd43140,17'd43141,17'd43142,17'd43143,17'd43144,17'd43145,17'd43146,17'd43147,17'd43148,17'd43149,17'd43150,17'd43151,17'd43152,17'd43153,17'd41581,17'd42739,17'd42882,17'd41582,17'd43154,17'd43155,17'd43156,17'd43019,17'd43020,17'd42749,17'd25030,17'd30126,17'd23917,17'd23384,17'd29242,17'd29241,17'd31029,17'd23386,17'd23386,17'd23732,17'd24249,17'd29375,17'd34467,17'd28596,17'd28717,17'd28850,17'd28369,17'd28600,17'd26064,17'd26062,17'd31351,17'd42436,17'd40958,17'd40367,17'd32017,17'd32355,17'd37250,17'd29248,17'd33656,17'd32507,17'd33654,17'd27642,17'd35426,17'd32016,17'd27371,17'd28853,17'd43157,17'd34278,17'd43158,17'd35295,17'd42603,17'd21529,17'd42439,17'd43159,17'd22008,17'd22504,17'd42744,17'd29240,17'd43022,17'd28253,17'd26174,17'd35578,17'd26782,17'd26903,17'd28481,17'd28481,17'd27639,17'd33815,17'd27371,17'd26781,17'd26901,17'd29245,17'd29245,17'd38025,17'd37907,17'd41582,17'd42600,17'd39436,17'd39741,17'd42891,17'd42606,17'd27644,17'd43160,17'd43023,17'd40063,17'd43161,17'd42446,17'd43162,17'd43163,17'd43025,17'd43164,17'd43165,17'd43166,17'd38668,17'd24902,17'd33340,17'd25173,17'd28130,17'd25565,17'd26285,17'd24583,17'd28602,17'd27765,17'd23725,17'd23558,17'd24416,17'd43167,17'd24095,17'd43168,17'd43169,17'd43170,17'd43031,17'd43171,17'd43172,17'd43173,17'd43174,17'd43175,17'd43176,17'd43177,17'd43178,17'd43179,17'd43040,17'd43180,17'd43181,17'd38566,17'd22251,17'd18619,17'd18132,17'd21772,17'd43182,17'd43043,17'd38845,17'd36734,17'd12906,17'd29161,17'd12160,17'd7499,17'd31891,17'd30637,17'd42910,17'd43045,17'd5156,17'd41891,17'd43183,17'd4671,17'd40395,17'd39468,17'd6067,17'd4683,17'd5327,17'd38442,17'd4016,17'd43046,17'd43046,17'd5476,17'd5142,17'd7654,17'd43184,17'd43048,17'd43049,17'd43050,17'd43185,17'd43186,17'd43187,17'd42777,17'd42914,17'd3357,17'd43188,17'd3043,17'd43055,17'd43189,17'd43190,17'd43191,17'd38328,17'd42781,17'd42921,17'd43058,17'd42477,17'd2723,17'd41479,17'd9530,17'd5493,17'd18629,17'd11587,17'd39033,17'd38580,17'd38581,17'd16492,17'd16492,17'd6418,17'd6418,17'd7364,17'd7878,17'd9124,17'd7705,17'd8187,17'd6416,17'd7365,17'd5194,17'd3744,17'd3895,17'd1261,17'd1401,17'd1680,17'd2559,17'd2764,17'd605,17'd424,17'd203,17'd195,17'd946
},
'{
17'd3903,17'd3903,17'd3902,17'd4891,17'd3902,17'd3902,17'd4892,17'd14743,17'd3252,17'd1688,17'd1127,17'd466,17'd3905,17'd19,17'd18,17'd3905,17'd18,17'd18,17'd980,17'd980,17'd4430,17'd4091,17'd3104,17'd2264,17'd1974,17'd1282,17'd1135,17'd1137,17'd992,17'd18275,17'd995,17'd22269,17'd14873,17'd2615,17'd43060,17'd2445,17'd3928,17'd20876,17'd32734,17'd18767,17'd43192,17'd43193,17'd43194,17'd43061,17'd17689,17'd17204,17'd19006,17'd19006,17'd43062,17'd21039,17'd40260,17'd41166,17'd43065,17'd38734,17'd42790,17'd42789,17'd40112,17'd43195,17'd42345,17'd43196,17'd41489,17'd42655,17'd40112,17'd41014,17'd42931,17'd43197,17'd42790,17'd42656,17'd43067,17'd43198,17'd42792,17'd19266,17'd9988,17'd9843,17'd11090,17'd43199,17'd42499,17'd6306,17'd4924,17'd43069,17'd43200,17'd43071,17'd6312,17'd43201,17'd43202,17'd43203,17'd43204,17'd43205,17'd42936,17'd43074,17'd43206,17'd43207,17'd43208,17'd43209,17'd43210,17'd43211,17'd43212,17'd7278,17'd7279,17'd43213,17'd43214,17'd43215,17'd43216,17'd43217,17'd43218,17'd13888,17'd9196,17'd24545,17'd8729,17'd16067,17'd8874,17'd9344,17'd8874,17'd9038,17'd14811,17'd9042,17'd17600,17'd9743,17'd9479,17'd26152,17'd11808,17'd24995,17'd25927,17'd28460,17'd28461,17'd28818,17'd28816,17'd27004,17'd24856,17'd24707,17'd24209,17'd22472,17'd21985,17'd19533,17'd11275,17'd11275,17'd11275,17'd11275,17'd18326,17'd18326,17'd28821,17'd11525,17'd42674,17'd19278,17'd16912,17'd9885,17'd9479,17'd9479,17'd15187,17'd15187,17'd10743,17'd10743,17'd11277,17'd11276,17'd11670,17'd11527,17'd19282,17'd11132,17'd27743,17'd20910,17'd18447,17'd14002,17'd29793,17'd30984,17'd31140,17'd33582,17'd41795,17'd33579,17'd30086,17'd32603,17'd42948,17'd41659,17'd21670,17'd18445,17'd43219,17'd43220,17'd43221,17'd43222,17'd42368,17'd40891,17'd40891,17'd43086,17'd43087,17'd43088,17'd43089,17'd42236,17'd41353,17'd42953,17'd41666,17'd40615,17'd43223,17'd43224,17'd43225,17'd43226,17'd43227,17'd43228,17'd43229,17'd43230,17'd43231,17'd43232,17'd43233,17'd43234,17'd43235,17'd42544,17'd43236,17'd43237,17'd43238,17'd43239,17'd43240,17'd43241,17'd43242,17'd43243,17'd43244,17'd43245,17'd43246,17'd43247,17'd43248,17'd43249,17'd43250,17'd43251,17'd42395,17'd43252,17'd43253,17'd43254,17'd43255,17'd40927,17'd43256,17'd43257,17'd43258,17'd40642,17'd41973,17'd43259,17'd43260,17'd43261,17'd43262,17'd43263,17'd43264,17'd43265,17'd43266,17'd43267,17'd43268,17'd43269,17'd43270,17'd43271,17'd43135,17'd35137,17'd43272,17'd43273,17'd35971,17'd35972,17'd39887,17'd43274,17'd43275,17'd37102,17'd43276,17'd43277,17'd43278,17'd42430,17'd43279,17'd42876,17'd43280,17'd43144,17'd43281,17'd43282,17'd43149,17'd43283,17'd43284,17'd43152,17'd43153,17'd41581,17'd42739,17'd42882,17'd41417,17'd41418,17'd43285,17'd43286,17'd43287,17'd43288,17'd29970,17'd25030,17'd28977,17'd23731,17'd23564,17'd23918,17'd29527,17'd23920,17'd23386,17'd29827,17'd30275,17'd24249,17'd29375,17'd34467,17'd33951,17'd33000,17'd28369,17'd28369,17'd28600,17'd26064,17'd25949,17'd27260,17'd43289,17'd41108,17'd32506,17'd32355,17'd32355,17'd32018,17'd33486,17'd33656,17'd32507,17'd28134,17'd31353,17'd32016,17'd30735,17'd43290,17'd28853,17'd43291,17'd43292,17'd43293,17'd34110,17'd33797,17'd42305,17'd43294,17'd43295,17'd43296,17'd22326,17'd29374,17'd28718,17'd29970,17'd28253,17'd27514,17'd35578,17'd26782,17'd26903,17'd28481,17'd28481,17'd27639,17'd33815,17'd27371,17'd33963,17'd28726,17'd29246,17'd28727,17'd38025,17'd37907,17'd42600,17'd43297,17'd43298,17'd39741,17'd42891,17'd35306,17'd34303,17'd43160,17'd43023,17'd36410,17'd42751,17'd43299,17'd43300,17'd43301,17'd43302,17'd43164,17'd43303,17'd43304,17'd36152,17'd28849,17'd23559,17'd23725,17'd27765,17'd25708,17'd24583,17'd26174,17'd33009,17'd27765,17'd23725,17'd23558,17'd30126,17'd43305,17'd43306,17'd43307,17'd43308,17'd43309,17'd43310,17'd43311,17'd20196,17'd43173,17'd40534,17'd38425,17'd43312,17'd43313,17'd43314,17'd22922,17'd43040,17'd43315,17'd43316,17'd38313,17'd22251,17'd18619,17'd19478,17'd18131,17'd43182,17'd43317,17'd39013,17'd37286,17'd36031,17'd11710,17'd13678,17'd7499,17'd31891,17'd31245,17'd5153,17'd43045,17'd4526,17'd33992,17'd4362,17'd4831,17'd39313,17'd39468,17'd6067,17'd4683,17'd5328,17'd5144,17'd41612,17'd42628,17'd43046,17'd5476,17'd33531,17'd7490,17'd43184,17'd43318,17'd43319,17'd43320,17'd43321,17'd42323,17'd43187,17'd43322,17'd43323,17'd43324,17'd43188,17'd43325,17'd43326,17'd43189,17'd43190,17'd43191,17'd2716,17'd43327,17'd43328,17'd43329,17'd42477,17'd42478,17'd3560,17'd41001,17'd41907,17'd18629,17'd11587,17'd39182,17'd43330,17'd38581,17'd16492,17'd16492,17'd6418,17'd6418,17'd6418,17'd7878,17'd9124,17'd9124,17'd7537,17'd6416,17'd7365,17'd5194,17'd3744,17'd5193,17'd229,17'd1401,17'd2417,17'd2559,17'd2922,17'd1394,17'd1525,17'd43331,17'd417,17'd946
},
'{
17'd3903,17'd3903,17'd4244,17'd4891,17'd3902,17'd4243,17'd25384,17'd14743,17'd3252,17'd4247,17'd466,17'd466,17'd18,17'd19,17'd18,17'd3905,17'd18,17'd1128,17'd3906,17'd3906,17'd27444,17'd3908,17'd3104,17'd2264,17'd1974,17'd16966,17'd1559,17'd1138,17'd17079,17'd18275,17'd995,17'd14451,17'd43332,17'd2615,17'd43060,17'd2445,17'd21798,17'd43333,17'd32734,17'd31264,17'd43334,17'd34517,17'd43335,17'd43336,17'd17689,17'd19006,17'd20292,17'd20292,17'd43337,17'd43063,17'd43338,17'd40261,17'd43065,17'd38469,17'd41632,17'd43339,17'd40112,17'd43340,17'd42345,17'd43341,17'd42207,17'd40112,17'd43342,17'd39802,17'd43343,17'd41914,17'd41487,17'd42656,17'd43344,17'd34528,17'd43345,17'd43346,17'd10566,17'd42793,17'd43347,17'd6467,17'd11089,17'd43348,17'd5086,17'd43069,17'd43349,17'd42501,17'd43350,17'd42797,17'd42934,17'd43351,17'd6161,17'd43352,17'd42936,17'd42936,17'd43353,17'd43354,17'd43355,17'd43209,17'd43210,17'd43356,17'd43357,17'd43358,17'd43359,17'd43360,17'd43361,17'd43362,17'd37849,17'd43217,17'd43218,17'd13888,17'd9196,17'd8573,17'd22473,17'd16067,17'd8874,17'd13887,17'd8873,17'd8873,17'd14811,17'd9042,17'd17600,17'd9346,17'd10742,17'd26152,17'd24029,17'd19408,17'd28107,17'd28460,17'd28461,17'd28818,17'd28816,17'd27004,17'd24856,17'd24707,17'd24362,17'd16442,17'd21985,17'd19533,17'd11275,17'd11275,17'd11808,17'd11808,17'd18326,17'd11398,17'd12584,17'd11400,17'd10331,17'd9884,17'd9885,17'd9885,17'd9479,17'd9479,17'd15187,17'd9345,17'd10743,17'd10743,17'd12116,17'd14928,17'd10479,17'd11527,17'd19282,17'd11132,17'd27743,17'd25144,17'd18447,17'd41793,17'd42676,17'd31450,17'd33736,17'd33582,17'd41795,17'd33581,17'd30234,17'd33099,17'd43083,17'd41659,17'd21670,17'd43363,17'd43364,17'd43364,17'd43221,17'd43222,17'd42368,17'd40891,17'd40751,17'd43086,17'd43365,17'd43366,17'd43089,17'd42236,17'd42527,17'd42953,17'd43367,17'd43368,17'd37999,17'd43369,17'd42686,17'd43370,17'd43371,17'd43372,17'd43373,17'd43374,17'd43375,17'd43376,17'd42850,17'd43377,17'd41375,17'd42117,17'd41060,17'd41953,17'd43378,17'd43379,17'd43380,17'd43381,17'd43382,17'd43383,17'd43384,17'd43385,17'd39688,17'd43386,17'd43387,17'd43388,17'd43389,17'd43390,17'd43391,17'd43392,17'd43393,17'd43394,17'd43395,17'd40477,17'd43396,17'd43397,17'd41694,17'd42992,17'd43398,17'd43399,17'd43400,17'd40488,17'd43401,17'd43402,17'd43403,17'd43265,17'd43404,17'd43405,17'd40938,17'd43406,17'd43407,17'd33448,17'd43408,17'd35834,17'd43409,17'd43273,17'd43410,17'd43411,17'd43412,17'd43412,17'd38393,17'd43413,17'd43414,17'd43415,17'd43416,17'd43417,17'd42430,17'd43013,17'd43418,17'd42876,17'd43419,17'd43420,17'd43421,17'd43283,17'd43422,17'd43423,17'd39273,17'd41581,17'd42739,17'd42882,17'd41417,17'd43424,17'd43425,17'd33157,17'd43288,17'd43020,17'd28484,17'd25030,17'd28977,17'd23731,17'd23564,17'd24086,17'd30424,17'd23920,17'd29826,17'd23566,17'd30275,17'd24249,17'd29375,17'd34467,17'd33951,17'd33000,17'd27882,17'd27882,17'd28130,17'd30606,17'd25833,17'd33478,17'd43426,17'd42889,17'd32506,17'd32507,17'd32355,17'd37250,17'd32018,17'd33656,17'd32193,17'd32354,17'd31352,17'd34637,17'd27027,17'd33499,17'd28725,17'd43157,17'd43292,17'd43427,17'd23044,17'd33946,17'd43428,17'd43429,17'd43430,17'd43431,17'd22326,17'd29686,17'd24417,17'd29970,17'd25565,17'd27515,17'd33499,17'd33963,17'd26903,17'd28481,17'd34300,17'd43432,17'd33815,17'd27371,17'd33963,17'd26901,17'd34632,17'd35441,17'd38025,17'd41109,17'd43433,17'd43434,17'd43298,17'd33308,17'd42891,17'd42606,17'd27644,17'd43160,17'd43023,17'd29549,17'd43435,17'd43436,17'd43437,17'd43438,17'd43302,17'd43439,17'd43440,17'd43441,17'd33971,17'd23564,17'd24246,17'd23726,17'd27765,17'd27766,17'd24583,17'd26174,17'd33009,17'd25951,17'd23912,17'd23558,17'd30126,17'd43305,17'd43306,17'd43307,17'd43442,17'd43443,17'd43444,17'd43445,17'd43446,17'd43447,17'd43448,17'd43449,17'd36572,17'd23607,17'd43450,17'd29587,17'd43451,17'd38435,17'd43452,17'd19985,17'd19087,17'd37940,17'd18021,17'd40244,17'd43453,17'd43454,17'd38439,17'd22767,17'd28186,17'd12905,17'd13800,17'd6220,17'd30333,17'd28536,17'd5144,17'd5757,17'd5155,17'd33992,17'd4362,17'd4672,17'd42772,17'd39468,17'd6067,17'd4683,17'd4841,17'd5144,17'd5604,17'd32550,17'd42628,17'd5476,17'd4988,17'd43455,17'd43456,17'd43457,17'd33198,17'd43458,17'd43321,17'd43459,17'd40851,17'd43460,17'd3529,17'd43324,17'd43188,17'd43325,17'd3044,17'd43461,17'd43190,17'd43191,17'd39480,17'd43056,17'd43057,17'd43329,17'd42477,17'd3378,17'd41479,17'd9530,17'd5493,17'd43462,17'd11587,17'd39033,17'd38580,17'd38581,17'd16492,17'd16623,17'd6418,17'd6418,17'd6418,17'd7878,17'd9124,17'd7705,17'd8187,17'd6416,17'd7365,17'd5194,17'd3744,17'd3895,17'd1261,17'd1401,17'd2417,17'd3742,17'd7210,17'd781,17'd1408,17'd1382,17'd42786,17'd1951
},
'{
17'd3903,17'd3903,17'd4244,17'd4891,17'd3902,17'd3902,17'd4892,17'd14743,17'd3252,17'd4247,17'd466,17'd2,17'd18,17'd19,17'd18,17'd3905,17'd18,17'd1128,17'd980,17'd980,17'd4430,17'd3595,17'd2941,17'd2263,17'd1974,17'd1839,17'd1559,17'd1137,17'd992,17'd18275,17'd2790,17'd14451,17'd43332,17'd2614,17'd32732,17'd2445,17'd21798,17'd43333,17'd43463,17'd18767,17'd43192,17'd32891,17'd43464,17'd43336,17'd19893,17'd19006,17'd20292,17'd18884,17'd19755,17'd21039,17'd18300,17'd40261,17'd43065,17'd38878,17'd38346,17'd40110,17'd40112,17'd42205,17'd42491,17'd43341,17'd42207,17'd40112,17'd40112,17'd41014,17'd43465,17'd41914,17'd41487,17'd42656,17'd43344,17'd34528,17'd43466,17'd43467,17'd9844,17'd10696,17'd43468,17'd43469,17'd42499,17'd6306,17'd4924,17'd43069,17'd40730,17'd42501,17'd43470,17'd6153,17'd42934,17'd43351,17'd43471,17'd43352,17'd42936,17'd42936,17'd43472,17'd43354,17'd43355,17'd43473,17'd43210,17'd43356,17'd43357,17'd43474,17'd43475,17'd43476,17'd7281,17'd43477,17'd43478,17'd43479,17'd43218,17'd13888,17'd9196,17'd8572,17'd8569,17'd9194,17'd8874,17'd15944,17'd8873,17'd8873,17'd14811,17'd9042,17'd17600,17'd9346,17'd10742,17'd26152,17'd24029,17'd21505,17'd27004,17'd28460,17'd28461,17'd28818,17'd28816,17'd26370,17'd24856,17'd24707,17'd24362,17'd16442,17'd21985,17'd19533,17'd11275,17'd11275,17'd11808,17'd11808,17'd18326,17'd18326,17'd28821,17'd11525,17'd29335,17'd19278,17'd10024,17'd9885,17'd9479,17'd9479,17'd15187,17'd9345,17'd10743,17'd10743,17'd12116,17'd11276,17'd11670,17'd11527,17'd19532,17'd11132,17'd27743,17'd25144,17'd18447,17'd41659,17'd42676,17'd31450,17'd33736,17'd33735,17'd33581,17'd30085,17'd30086,17'd32603,17'd30684,17'd41659,17'd43480,17'd43363,17'd43364,17'd43364,17'd43481,17'd43482,17'd42368,17'd40891,17'd40751,17'd42234,17'd43483,17'd43366,17'd43484,17'd43485,17'd43486,17'd40895,17'd43487,17'd43488,17'd43489,17'd42819,17'd43490,17'd43491,17'd43492,17'd43493,17'd43494,17'd43495,17'd43496,17'd43497,17'd43498,17'd40636,17'd43499,17'd43500,17'd43501,17'd41814,17'd43502,17'd43503,17'd43504,17'd43505,17'd43506,17'd43507,17'd43508,17'd43509,17'd43510,17'd43511,17'd43512,17'd43513,17'd43514,17'd43515,17'd43516,17'd43517,17'd43518,17'd43519,17'd43520,17'd43521,17'd41371,17'd41223,17'd43522,17'd43523,17'd40175,17'd40910,17'd43524,17'd43525,17'd43526,17'd43527,17'd43528,17'd42858,17'd43529,17'd43530,17'd43531,17'd43532,17'd39407,17'd33282,17'd43003,17'd38644,17'd43533,17'd43273,17'd43410,17'd43534,17'd36384,17'd39262,17'd38393,17'd43535,17'd43536,17'd43537,17'd43538,17'd43539,17'd42430,17'd43013,17'd43540,17'd43013,17'd43541,17'd43542,17'd43421,17'd43543,17'd43422,17'd43544,17'd43545,17'd43546,17'd41997,17'd43547,17'd43289,17'd43548,17'd43549,17'd43550,17'd43020,17'd43020,17'd25317,17'd25030,17'd24416,17'd28852,17'd28849,17'd23731,17'd30424,17'd23733,17'd29975,17'd29827,17'd30275,17'd24249,17'd30431,17'd24252,17'd33951,17'd33000,17'd27511,17'd25709,17'd28594,17'd27767,17'd25833,17'd43551,17'd43552,17'd39276,17'd32356,17'd32507,17'd32507,17'd32018,17'd32018,17'd32507,17'd32193,17'd32354,17'd31352,17'd33163,17'd26902,17'd33815,17'd27515,17'd43553,17'd43554,17'd43555,17'd33796,17'd32663,17'd43556,17'd43557,17'd43558,17'd36846,17'd22328,17'd23386,17'd24745,17'd29970,17'd25565,17'd27515,17'd35304,17'd33963,17'd28725,17'd28481,17'd34300,17'd43432,17'd33815,17'd27371,17'd33963,17'd28726,17'd34768,17'd35441,17'd33791,17'd38153,17'd43297,17'd43559,17'd43560,17'd33308,17'd42891,17'd43561,17'd36868,17'd43160,17'd43562,17'd36551,17'd43435,17'd43563,17'd43564,17'd43565,17'd43566,17'd43567,17'd43440,17'd38171,17'd43568,17'd23384,17'd23560,17'd23913,17'd25567,17'd25566,17'd25708,17'd25565,17'd33333,17'd27765,17'd27509,17'd24894,17'd30895,17'd43569,17'd39144,17'd43570,17'd43571,17'd21403,17'd43572,17'd43573,17'd43574,17'd43575,17'd42764,17'd43576,17'd43577,17'd43578,17'd20369,17'd43579,17'd43451,17'd43580,17'd43452,17'd19985,17'd19087,17'd43581,17'd21772,17'd43582,17'd43583,17'd43317,17'd38438,17'd37556,17'd38701,17'd13046,17'd13800,17'd6219,17'd31553,17'd31716,17'd4997,17'd4839,17'd41459,17'd4998,17'd4362,17'd4832,17'd41455,17'd33839,17'd6067,17'd4683,17'd4841,17'd5145,17'd43584,17'd43585,17'd42628,17'd42630,17'd36022,17'd5321,17'd43586,17'd43587,17'd43588,17'd43589,17'd43321,17'd43459,17'd40851,17'd43052,17'd43590,17'd43591,17'd43592,17'd43593,17'd43594,17'd43461,17'd42329,17'd43595,17'd39480,17'd43056,17'd43057,17'd42921,17'd42477,17'd42334,17'd3561,17'd41001,17'd41625,17'd43462,17'd39790,17'd39033,17'd38580,17'd38581,17'd43596,17'd16623,17'd6418,17'd6417,17'd6418,17'd7705,17'd38460,17'd9124,17'd7537,17'd6416,17'd7365,17'd4869,17'd3744,17'd3895,17'd1261,17'd1401,17'd2417,17'd6407,17'd7210,17'd10911,17'd203,17'd201,17'd1813,17'd1951
},
'{
17'd6420,17'd4892,17'd4244,17'd3902,17'd29756,17'd31905,17'd4892,17'd4245,17'd2422,17'd2594,17'd1416,17'd3905,17'd20404,17'd3905,17'd3905,17'd3905,17'd11,17'd11,17'd980,17'd652,17'd289,17'd3595,17'd2941,17'd2601,17'd2266,17'd1839,17'd1559,17'd991,17'd992,17'd18275,17'd483,17'd668,17'd2613,17'd835,17'd2795,17'd37577,17'd43597,17'd20876,17'd32734,17'd14879,17'd16018,17'd33855,17'd43598,17'd43336,17'd19128,17'd12681,17'd22630,17'd16658,17'd43599,17'd40864,17'd17450,17'd43600,17'd38344,17'd15390,17'd40721,17'd39956,17'd40420,17'd42654,17'd42491,17'd41636,17'd40725,17'd40420,17'd40726,17'd42930,17'd42931,17'd41914,17'd42203,17'd43601,17'd41327,17'd41921,17'd43466,17'd43346,17'd10120,17'd22635,17'd11233,17'd6466,17'd11089,17'd43348,17'd5086,17'd7089,17'd6473,17'd42501,17'd43602,17'd43201,17'd43603,17'd43604,17'd43605,17'd43606,17'd42936,17'd43607,17'd43608,17'd43354,17'd43609,17'd43610,17'd43611,17'd43211,17'd43612,17'd43613,17'd43614,17'd43615,17'd43616,17'd43617,17'd43618,17'd43619,17'd43620,17'd43621,17'd8573,17'd10027,17'd9621,17'd15684,17'd17480,17'd17480,17'd9194,17'd15684,17'd14811,17'd10175,17'd15682,17'd9346,17'd10743,17'd17719,17'd11274,17'd22992,17'd26872,17'd29923,17'd28571,17'd28462,17'd28230,17'd28107,17'd24856,17'd24707,17'd24209,17'd21361,17'd18327,17'd24029,17'd11275,17'd11275,17'd19533,17'd24029,17'd18326,17'd12583,17'd43622,17'd12423,17'd34826,17'd11671,17'd17965,17'd17965,17'd9479,17'd9479,17'd9479,17'd9479,17'd10743,17'd9341,17'd9741,17'd11135,17'd12863,17'd12863,17'd10476,17'd11132,17'd10474,17'd29203,17'd15810,17'd41510,17'd42676,17'd31140,17'd33885,17'd33735,17'd32936,17'd30233,17'd29340,17'd13518,17'd30684,17'd14002,17'd43480,17'd29342,17'd16907,17'd43623,17'd43624,17'd43482,17'd41938,17'd42522,17'd42813,17'd42951,17'd43625,17'd43626,17'd43627,17'd43628,17'd42080,17'd43629,17'd36088,17'd43630,17'd43631,17'd43632,17'd43633,17'd43634,17'd43635,17'd42961,17'd43636,17'd43637,17'd43638,17'd43639,17'd40174,17'd43640,17'd43641,17'd43642,17'd43643,17'd43644,17'd43645,17'd43646,17'd43647,17'd43648,17'd43649,17'd43650,17'd43651,17'd43652,17'd43653,17'd43654,17'd43108,17'd43655,17'd43656,17'd43657,17'd43658,17'd43659,17'd43660,17'd43661,17'd43662,17'd40914,17'd41370,17'd43663,17'd43664,17'd43665,17'd43666,17'd43667,17'd43668,17'd43669,17'd43670,17'd43671,17'd43672,17'd43673,17'd43674,17'd42130,17'd43675,17'd40800,17'd43676,17'd43677,17'd43678,17'd43679,17'd34076,17'd35552,17'd35962,17'd40350,17'd35971,17'd39887,17'd43680,17'd43681,17'd38265,17'd43682,17'd43683,17'd43684,17'd43685,17'd43013,17'd43278,17'd43686,17'd43687,17'd43688,17'd43421,17'd43689,17'd43423,17'd43690,17'd43691,17'd41862,17'd43692,17'd43434,17'd43693,17'd42885,17'd43549,17'd43694,17'd33156,17'd43695,17'd42749,17'd24898,17'd24416,17'd29102,17'd23562,17'd23916,17'd30431,17'd23565,17'd29975,17'd29686,17'd34137,17'd23917,17'd30431,17'd24416,17'd27637,17'd25177,17'd25177,17'd28369,17'd27767,17'd27639,17'd25707,17'd43019,17'd43433,17'd43696,17'd40367,17'd33654,17'd29380,17'd28728,17'd28372,17'd29380,17'd29247,17'd27884,17'd31352,17'd26901,17'd28853,17'd25949,17'd26174,17'd43553,17'd23739,17'd31499,17'd31346,17'd43697,17'd41275,17'd43698,17'd43699,17'd31500,17'd37116,17'd29827,17'd32007,17'd28484,17'd25565,17'd26530,17'd27371,17'd26901,17'd27259,17'd28482,17'd28481,17'd28481,17'd27514,17'd27640,17'd26902,17'd26901,17'd29245,17'd31352,17'd33941,17'd40824,17'd43700,17'd43701,17'd43702,17'd43703,17'd42891,17'd43704,17'd43705,17'd33508,17'd43706,17'd36551,17'd43707,17'd43708,17'd43709,17'd43710,17'd43711,17'd43024,17'd43712,17'd42612,17'd23739,17'd29242,17'd33672,17'd24245,17'd25709,17'd26402,17'd26287,17'd25565,17'd28130,17'd24079,17'd43713,17'd43714,17'd43715,17'd43716,17'd43717,17'd43718,17'd40971,17'd43719,17'd43720,17'd43721,17'd43722,17'd43723,17'd43724,17'd41881,17'd40387,17'd29137,17'd23961,17'd43725,17'd43726,17'd43727,17'd36885,17'd19714,17'd16955,17'd43581,17'd41452,17'd43728,17'd43729,17'd43730,17'd38438,17'd38845,17'd37429,17'd38316,17'd11578,17'd6554,17'd5162,17'd4526,17'd4998,17'd4836,17'd4999,17'd34157,17'd4358,17'd4515,17'd41612,17'd41458,17'd4189,17'd4689,17'd4684,17'd4999,17'd42462,17'd42631,17'd42631,17'd42630,17'd4988,17'd36438,17'd33833,17'd33198,17'd43731,17'd43732,17'd43733,17'd33528,17'd43734,17'd42324,17'd43323,17'd43591,17'd43735,17'd43736,17'd42918,17'd42919,17'd43737,17'd36595,17'd39026,17'd43738,17'd42781,17'd43739,17'd42194,17'd43740,17'd43741,17'd42043,17'd43742,17'd10790,17'd11048,17'd38202,17'd38580,17'd38203,17'd43596,17'd16492,17'd6258,17'd6416,17'd7537,17'd7705,17'd9124,17'd7364,17'd8187,17'd8186,17'd4882,17'd4713,17'd3391,17'd3895,17'd1261,17'd1261,17'd6407,17'd2905,17'd24323,17'd1408,17'd43743,17'd43744,17'd1530,17'd1951
},
'{
17'd6420,17'd4892,17'd4244,17'd4891,17'd29756,17'd29756,17'd4244,17'd4245,17'd2422,17'd4247,17'd1416,17'd3905,17'd20404,17'd18,17'd17,17'd3905,17'd11,17'd11,17'd652,17'd29,17'd809,17'd31,17'd2941,17'd2943,17'd2785,17'd1839,17'd1559,17'd991,17'd992,17'd481,17'd483,17'd64,17'd43745,17'd835,17'd2620,17'd37577,17'd43597,17'd20876,17'd43463,17'd18646,17'd43746,17'd33855,17'd43598,17'd42485,17'd19382,17'd12681,17'd22630,17'd12532,17'd43747,17'd40864,17'd43748,17'd43600,17'd38344,17'd15390,17'd43749,17'd43750,17'd40420,17'd42654,17'd42654,17'd41636,17'd40725,17'd43342,17'd40726,17'd39803,17'd39639,17'd41914,17'd42203,17'd43601,17'd41327,17'd34190,17'd43466,17'd43467,17'd10120,17'd7581,17'd6466,17'd10695,17'd43068,17'd6306,17'd4924,17'd7253,17'd6473,17'd42662,17'd42663,17'd43201,17'd43751,17'd43752,17'd43605,17'd43606,17'd42936,17'd43206,17'd43753,17'd43354,17'd43754,17'd43610,17'd43611,17'd43755,17'd39064,17'd43756,17'd7773,17'd43757,17'd43758,17'd43759,17'd43760,17'd43761,17'd43762,17'd43763,17'd8571,17'd8883,17'd15682,17'd8874,17'd17480,17'd17848,17'd9194,17'd15684,17'd14811,17'd10175,17'd9043,17'd9346,17'd10743,17'd17719,17'd25280,17'd24363,17'd27621,17'd29923,17'd28571,17'd28461,17'd35376,17'd28347,17'd27004,17'd24030,17'd24209,17'd21361,17'd18327,17'd24029,17'd11275,17'd11275,17'd19533,17'd24029,17'd18326,17'd12583,17'd43622,17'd12423,17'd34826,17'd17847,17'd10170,17'd17965,17'd9479,17'd9479,17'd9479,17'd9479,17'd10743,17'd11136,17'd9884,17'd11135,17'd12863,17'd12863,17'd11132,17'd11132,17'd10474,17'd10474,17'd10737,17'd28938,17'd42676,17'd33736,17'd33885,17'd33100,17'd39662,17'd31138,17'd30231,17'd14526,17'd12995,17'd12113,17'd18682,17'd18915,17'd43764,17'd42366,17'd43765,17'd42233,17'd43766,17'd42522,17'd43767,17'd43768,17'd43769,17'd43626,17'd43770,17'd43771,17'd42080,17'd43629,17'd43772,17'd35254,17'd43773,17'd43774,17'd43775,17'd43491,17'd43776,17'd43777,17'd43778,17'd43779,17'd43780,17'd43781,17'd43125,17'd43782,17'd42251,17'd43783,17'd43784,17'd43785,17'd43786,17'd43787,17'd43788,17'd43789,17'd43790,17'd43791,17'd43792,17'd43793,17'd43794,17'd43795,17'd43796,17'd43797,17'd43798,17'd43799,17'd43800,17'd43801,17'd43802,17'd43803,17'd43804,17'd43805,17'd41072,17'd43806,17'd43807,17'd43808,17'd43809,17'd43810,17'd43811,17'd43812,17'd43813,17'd43814,17'd43815,17'd43816,17'd43817,17'd43818,17'd43819,17'd43820,17'd43821,17'd43822,17'd43823,17'd43824,17'd35407,17'd36522,17'd43825,17'd40350,17'd35972,17'd39887,17'd43826,17'd43827,17'd43828,17'd43829,17'd43683,17'd43684,17'd43142,17'd43013,17'd43278,17'd42734,17'd43830,17'd43831,17'd43150,17'd43283,17'd42296,17'd43153,17'd43832,17'd43833,17'd43692,17'd43559,17'd43834,17'd42885,17'd43835,17'd43836,17'd43837,17'd43838,17'd43022,17'd24898,17'd23916,17'd23563,17'd23562,17'd24252,17'd24249,17'd23565,17'd32191,17'd30128,17'd34137,17'd23917,17'd23916,17'd24416,17'd27637,17'd25177,17'd25320,17'd28369,17'd41999,17'd28009,17'd28252,17'd40825,17'd40366,17'd37777,17'd32506,17'd33654,17'd28372,17'd28857,17'd28372,17'd29380,17'd29247,17'd27884,17'd29379,17'd26901,17'd28724,17'd26062,17'd27766,17'd43553,17'd43839,17'd43840,17'd23041,17'd21693,17'd43841,17'd34757,17'd43842,17'd43843,17'd23569,17'd28976,17'd25180,17'd28484,17'd25565,17'd26530,17'd27371,17'd26901,17'd27371,17'd28009,17'd28482,17'd28482,17'd27883,17'd43290,17'd26781,17'd28726,17'd29246,17'd31352,17'd32005,17'd42600,17'd41997,17'd43844,17'd43702,17'd43703,17'd42891,17'd43561,17'd36868,17'd33508,17'd43845,17'd43846,17'd43707,17'd43847,17'd43848,17'd43849,17'd26068,17'd43850,17'd43851,17'd25440,17'd23739,17'd29827,17'd43852,17'd23559,17'd33484,17'd33333,17'd32364,17'd26287,17'd28130,17'd24080,17'd25027,17'd43853,17'd43715,17'd43716,17'd43854,17'd43855,17'd43856,17'd43857,17'd43858,17'd43859,17'd43860,17'd43861,17'd43862,17'd43863,17'd41603,17'd43864,17'd43865,17'd43866,17'd43726,17'd43867,17'd36885,17'd19480,17'd16955,17'd17534,17'd41297,17'd43728,17'd43868,17'd43730,17'd38438,17'd38845,17'd37557,17'd38316,17'd11578,17'd27935,17'd34921,17'd4525,17'd33691,17'd4524,17'd4524,17'd34157,17'd34157,17'd33691,17'd41458,17'd33533,17'd4189,17'd4689,17'd4684,17'd5155,17'd4515,17'd42631,17'd42631,17'd42630,17'd4988,17'd5908,17'd33833,17'd33362,17'd43731,17'd43869,17'd43733,17'd33528,17'd43734,17'd43870,17'd43871,17'd43872,17'd42778,17'd43873,17'd43874,17'd42919,17'd43737,17'd36595,17'd41310,17'd43875,17'd43876,17'd3056,17'd42194,17'd43740,17'd43741,17'd41906,17'd41002,17'd10790,17'd11048,17'd38202,17'd38580,17'd38580,17'd43596,17'd16492,17'd6258,17'd6416,17'd11336,17'd7705,17'd43877,17'd8506,17'd7537,17'd8186,17'd4882,17'd4713,17'd3391,17'd3895,17'd1261,17'd1261,17'd6407,17'd2905,17'd412,17'd939,17'd1102,17'd43878,17'd1530,17'd1530
},
'{
17'd6420,17'd25384,17'd4892,17'd4891,17'd32728,17'd31905,17'd4892,17'd4245,17'd2422,17'd4247,17'd1416,17'd3905,17'd1128,17'd1128,17'd3905,17'd3905,17'd11,17'd11,17'd652,17'd652,17'd289,17'd30,17'd3254,17'd2601,17'd2266,17'd1839,17'd1559,17'd1137,17'd992,17'd481,17'd62,17'd43745,17'd833,17'd835,17'd43879,17'd37577,17'd21798,17'd43880,17'd43881,17'd43882,17'd16018,17'd33855,17'd43598,17'd43883,17'd19006,17'd12681,17'd16658,17'd16658,17'd43599,17'd40864,17'd17450,17'd43600,17'd38344,17'd37315,17'd42047,17'd43750,17'd40420,17'd43195,17'd41635,17'd41636,17'd40573,17'd43342,17'd40726,17'd42930,17'd42931,17'd41914,17'd42203,17'd43884,17'd43885,17'd34190,17'd43466,17'd20032,17'd10120,17'd22635,17'd11233,17'd6467,17'd43886,17'd43348,17'd5086,17'd7253,17'd6632,17'd42662,17'd43887,17'd6153,17'd43888,17'd6325,17'd43889,17'd43890,17'd42936,17'd42936,17'd43891,17'd43892,17'd43609,17'd43610,17'd43893,17'd43894,17'd43895,17'd43896,17'd43897,17'd37062,17'd43898,17'd43899,17'd43900,17'd43901,17'd43902,17'd43763,17'd8728,17'd8881,17'd9044,17'd10174,17'd14811,17'd14811,17'd9194,17'd15684,17'd14811,17'd9189,17'd21984,17'd19415,17'd9471,17'd17124,17'd11274,17'd24995,17'd27123,17'd29923,17'd28571,17'd28462,17'd28103,17'd28107,17'd24537,17'd24030,17'd24209,17'd22472,17'd18327,17'd24029,17'd11275,17'd11275,17'd24029,17'd24029,17'd36206,17'd12583,17'd43622,17'd12423,17'd34826,17'd17847,17'd10169,17'd9885,17'd9479,17'd9479,17'd9479,17'd9479,17'd10743,17'd9341,17'd12116,17'd11135,17'd12863,17'd12863,17'd11132,17'd11132,17'd10472,17'd27738,17'd32137,17'd28938,17'd30984,17'd33583,17'd33885,17'd43903,17'd32936,17'd31138,17'd30231,17'd13760,17'd13365,17'd12259,17'd21822,17'd43219,17'd43904,17'd43905,17'd42367,17'd43906,17'd42368,17'd43907,17'd43908,17'd43909,17'd43769,17'd43626,17'd43910,17'd43771,17'd43911,17'd43629,17'd43912,17'd43913,17'd43914,17'd43915,17'd43916,17'd43634,17'd43917,17'd43918,17'd43919,17'd43920,17'd43921,17'd43922,17'd40646,17'd43923,17'd43924,17'd43925,17'd43926,17'd43927,17'd43928,17'd43929,17'd43930,17'd43931,17'd43932,17'd43933,17'd43934,17'd43935,17'd43936,17'd43937,17'd43938,17'd43939,17'd43940,17'd43941,17'd43942,17'd41832,17'd43943,17'd43944,17'd43945,17'd43946,17'd43947,17'd43522,17'd43948,17'd40471,17'd43949,17'd43950,17'd43951,17'd43922,17'd43952,17'd43953,17'd43954,17'd43955,17'd43956,17'd43957,17'd43958,17'd43959,17'd43821,17'd43960,17'd43961,17'd33452,17'd36247,17'd35835,17'd43825,17'd40349,17'd36385,17'd39887,17'd43962,17'd43963,17'd43964,17'd43965,17'd43966,17'd43684,17'd43967,17'd43968,17'd43141,17'd43969,17'd43970,17'd43971,17'd43150,17'd43972,17'd43423,17'd41861,17'd43832,17'd43973,17'd43974,17'd43559,17'd43975,17'd42742,17'd43976,17'd43977,17'd43978,17'd43979,17'd43836,17'd24898,17'd34467,17'd28849,17'd28852,17'd24415,17'd24087,17'd29376,17'd29828,17'd30128,17'd34137,17'd24087,17'd30431,17'd24416,17'd25180,17'd25178,17'd25177,17'd25567,17'd28481,17'd28482,17'd33642,17'd43980,17'd40366,17'd34275,17'd31354,17'd33654,17'd28372,17'd28857,17'd28372,17'd28257,17'd28370,17'd27761,17'd29379,17'd26901,17'd28724,17'd28481,17'd28602,17'd43553,17'd43839,17'd43981,17'd43982,17'd21693,17'd43983,17'd43984,17'd43985,17'd43986,17'd29829,17'd28976,17'd25180,17'd28600,17'd25565,17'd26530,17'd27371,17'd27027,17'd28725,17'd33815,17'd26530,17'd26530,17'd27883,17'd43290,17'd26781,17'd28726,17'd29246,17'd31352,17'd32005,17'd43433,17'd41416,17'd43974,17'd43987,17'd43703,17'd42891,17'd43988,17'd43989,17'd43990,17'd43991,17'd29703,17'd43992,17'd43993,17'd42757,17'd43994,17'd43995,17'd43996,17'd43997,17'd43303,17'd34277,17'd23923,17'd24248,17'd23560,17'd28719,17'd25951,17'd33970,17'd25708,17'd24410,17'd24080,17'd23547,17'd43998,17'd36854,17'd43716,17'd43999,17'd44000,17'd44001,17'd44002,17'd44003,17'd44004,17'd31692,17'd44005,17'd44006,17'd44007,17'd41603,17'd43312,17'd43865,17'd22235,17'd17030,17'd44008,17'd36732,17'd21310,17'd18022,17'd17779,17'd22088,17'd43728,17'd43729,17'd43728,17'd38438,17'd38845,17'd39014,17'd38440,17'd12307,17'd27935,17'd34921,17'd33841,17'd44009,17'd4359,17'd4189,17'd33991,17'd33991,17'd33839,17'd41612,17'd33533,17'd4189,17'd44010,17'd5156,17'd4525,17'd42462,17'd42772,17'd42631,17'd42630,17'd4988,17'd5908,17'd44011,17'd33362,17'd5906,17'd43869,17'd44012,17'd33528,17'd43734,17'd43870,17'd43871,17'd44013,17'd44014,17'd42779,17'd44015,17'd44016,17'd43737,17'd44017,17'd41310,17'd43875,17'd43876,17'd3056,17'd44018,17'd43740,17'd3561,17'd42043,17'd40100,17'd10906,17'd11048,17'd38202,17'd38580,17'd44019,17'd43596,17'd16492,17'd6258,17'd6416,17'd11336,17'd11336,17'd9124,17'd7878,17'd8187,17'd8186,17'd4882,17'd4713,17'd3391,17'd3895,17'd1261,17'd445,17'd6407,17'd24323,17'd951,17'd202,17'd201,17'd44020,17'd1530,17'd1530
},
'{
17'd6420,17'd4892,17'd3902,17'd4891,17'd32728,17'd29756,17'd4244,17'd4245,17'd2422,17'd4247,17'd1416,17'd3905,17'd1128,17'd18,17'd17,17'd17,17'd19,17'd1128,17'd652,17'd29,17'd809,17'd1129,17'd2940,17'd3253,17'd2785,17'd1839,17'd1559,17'd1137,17'd992,17'd827,17'd16637,17'd483,17'd831,17'd998,17'd43879,17'd37577,17'd21798,17'd15250,17'd43881,17'd44021,17'd16018,17'd33855,17'd43598,17'd44022,17'd19006,17'd12532,17'd16658,17'd12531,17'd14472,17'd21346,17'd17211,17'd42045,17'd15266,17'd37315,17'd41631,17'd44023,17'd42653,17'd43195,17'd41635,17'd41634,17'd41170,17'd43342,17'd40726,17'd42930,17'd42931,17'd41914,17'd42342,17'd44024,17'd44025,17'd44026,17'd44027,17'd12067,17'd10119,17'd7581,17'd6466,17'd6305,17'd43068,17'd6306,17'd4924,17'd7253,17'd6632,17'd42662,17'd43602,17'd6153,17'd43888,17'd6325,17'd43889,17'd44028,17'd43074,17'd42938,17'd44029,17'd42354,17'd43754,17'd43610,17'd43893,17'd43894,17'd43895,17'd43896,17'd44030,17'd44031,17'd7774,17'd44032,17'd44033,17'd43901,17'd43902,17'd44034,17'd30672,17'd15297,17'd8720,17'd10174,17'd14811,17'd14811,17'd9194,17'd15684,17'd14811,17'd10175,17'd9043,17'd9339,17'd9341,17'd17719,17'd25280,17'd29488,17'd28105,17'd29923,17'd28571,17'd28462,17'd28103,17'd28107,17'd24537,17'd24030,17'd23170,17'd22472,17'd18327,17'd24029,17'd11808,17'd11808,17'd24029,17'd24029,17'd36481,17'd36481,17'd35799,17'd28821,17'd34956,17'd17847,17'd10024,17'd9885,17'd9479,17'd9479,17'd9479,17'd9479,17'd10743,17'd11136,17'd9884,17'd11135,17'd12863,17'd12863,17'd11132,17'd11132,17'd10472,17'd10474,17'd10853,17'd28938,17'd34391,17'd33737,17'd33885,17'd33100,17'd39662,17'd38368,17'd30231,17'd14809,17'd12995,17'd12113,17'd15810,17'd44035,17'd43904,17'd44036,17'd42367,17'd44037,17'd44038,17'd44039,17'd44040,17'd44041,17'd42952,17'd43089,17'd43910,17'd43771,17'd43911,17'd40148,17'd44042,17'd44043,17'd44044,17'd44045,17'd44046,17'd44047,17'd44048,17'd44049,17'd44050,17'd44051,17'd44052,17'd44053,17'd44054,17'd44055,17'd44056,17'd41061,17'd44057,17'd41066,17'd44058,17'd44059,17'd44060,17'd44061,17'd44062,17'd44063,17'd44064,17'd44065,17'd44066,17'd44067,17'd44068,17'd44069,17'd44070,17'd44071,17'd44072,17'd44073,17'd44057,17'd44074,17'd43927,17'd41535,17'd44075,17'd44076,17'd40327,17'd44077,17'd44078,17'd44079,17'd44080,17'd44081,17'd44082,17'd44083,17'd44084,17'd44085,17'd42130,17'd44086,17'd44087,17'd44088,17'd42863,17'd44089,17'd44090,17'd44091,17'd36247,17'd36522,17'd35406,17'd40349,17'd36384,17'd39887,17'd40946,17'd44092,17'd44093,17'd44094,17'd44095,17'd43684,17'd44096,17'd43686,17'd43540,17'd44097,17'd44098,17'd44099,17'd43283,17'd44100,17'd41861,17'd41861,17'd44101,17'd44102,17'd43844,17'd44103,17'd44104,17'd42597,17'd44105,17'd39591,17'd32996,17'd44106,17'd43694,17'd24895,17'd24249,17'd28722,17'd28975,17'd24090,17'd31033,17'd29530,17'd23216,17'd23215,17'd29099,17'd31033,17'd24249,17'd24416,17'd25030,17'd25178,17'd25177,17'd25567,17'd26062,17'd26530,17'd42147,17'd43298,17'd40366,17'd34105,17'd27642,17'd33654,17'd28372,17'd28857,17'd28728,17'd30587,17'd29104,17'd27761,17'd29379,17'd26901,17'd26903,17'd28481,17'd26064,17'd29825,17'd44107,17'd44108,17'd44109,17'd21693,17'd34881,17'd32664,17'd42601,17'd44110,17'd29829,17'd29689,17'd29976,17'd25435,17'd25565,17'd27514,17'd27371,17'd26901,17'd26782,17'd27883,17'd26530,17'd26530,17'd27883,17'd43290,17'd26781,17'd38537,17'd37513,17'd31352,17'd32005,17'd43434,17'd43692,17'd43974,17'd43987,17'd44111,17'd42605,17'd43561,17'd43989,17'd33508,17'd31855,17'd44112,17'd43992,17'd43993,17'd44113,17'd25441,17'd43849,17'd43996,17'd44114,17'd44115,17'd37533,17'd29686,17'd44116,17'd24744,17'd44117,17'd44118,17'd33174,17'd27766,17'd24410,17'd25028,17'd44119,17'd44120,17'd36854,17'd43716,17'd23392,17'd44121,17'd44122,17'd44123,17'd44124,17'd44125,17'd31692,17'd20196,17'd44126,17'd44127,17'd44128,17'd44129,17'd44130,17'd22214,17'd44131,17'd44132,17'd36025,17'd18375,17'd26710,17'd17654,17'd40985,17'd43728,17'd43729,17'd43728,17'd38439,17'd38845,17'd39014,17'd38440,17'd12307,17'd27935,17'd5157,17'd33992,17'd41299,17'd4515,17'd33838,17'd33838,17'd33991,17'd33839,17'd41612,17'd33533,17'd4189,17'd4689,17'd4847,17'd5155,17'd4358,17'd42772,17'd42772,17'd4830,17'd4988,17'd6206,17'd44011,17'd33362,17'd5906,17'd44133,17'd44012,17'd3527,17'd44134,17'd44135,17'd44136,17'd44137,17'd44138,17'd44139,17'd44140,17'd44141,17'd41309,17'd44017,17'd20706,17'd38328,17'd43876,17'd42476,17'd44018,17'd43740,17'd3561,17'd7849,17'd39947,17'd10906,17'd38458,17'd38334,17'd38580,17'd44019,17'd43596,17'd16492,17'd6258,17'd8186,17'd11335,17'd7537,17'd43877,17'd43877,17'd8507,17'd8186,17'd4882,17'd4713,17'd3391,17'd3895,17'd1261,17'd445,17'd6407,17'd24323,17'd951,17'd11445,17'd1247,17'd199,17'd1530,17'd1673
},
'{
17'd6420,17'd25384,17'd4243,17'd4891,17'd32728,17'd31905,17'd4892,17'd4245,17'd2422,17'd4247,17'd1416,17'd3905,17'd1128,17'd1128,17'd3905,17'd3905,17'd1128,17'd1128,17'd652,17'd29,17'd809,17'd1129,17'd2940,17'd2602,17'd2266,17'd1839,17'd1559,17'd1135,17'd16967,17'd827,17'd16637,17'd831,17'd1145,17'd998,17'd43879,17'd37577,17'd43597,17'd15250,17'd43881,17'd18526,17'd16018,17'd44142,17'd44143,17'd44022,17'd19006,17'd12532,17'd12531,17'd12531,17'd14472,17'd42340,17'd17211,17'd44144,17'd16174,17'd38594,17'd40866,17'd44145,17'd42653,17'd44146,17'd41916,17'd40725,17'd40572,17'd44147,17'd44148,17'd41014,17'd43343,17'd44149,17'd44150,17'd44151,17'd44152,17'd34189,17'd44027,17'd12067,17'd10119,17'd22635,17'd11233,17'd6626,17'd44153,17'd6306,17'd4924,17'd7253,17'd42796,17'd6313,17'd43602,17'd42797,17'd44154,17'd44155,17'd44156,17'd44028,17'd43074,17'd42936,17'd43891,17'd43892,17'd43355,17'd42670,17'd43893,17'd43894,17'd43895,17'd44157,17'd44158,17'd44159,17'd44160,17'd44161,17'd44162,17'd44163,17'd44164,17'd44165,17'd30672,17'd15297,17'd8720,17'd9039,17'd14811,17'd14811,17'd15684,17'd15684,17'd14811,17'd9189,17'd21984,17'd9337,17'd9471,17'd17124,17'd14673,17'd24995,17'd25927,17'd28343,17'd28818,17'd28345,17'd28103,17'd27121,17'd24537,17'd23512,17'd23170,17'd22472,17'd18327,17'd24029,17'd11808,17'd11274,17'd11397,17'd21985,17'd21985,17'd11397,17'd25280,17'd11399,17'd11400,17'd10329,17'd9884,17'd9741,17'd10742,17'd10742,17'd9479,17'd9479,17'd10742,17'd10743,17'd9741,17'd11135,17'd12863,17'd12863,17'd10991,17'd11133,17'd10472,17'd10474,17'd10853,17'd28938,17'd29937,17'd31140,17'd33885,17'd33735,17'd31449,17'd38368,17'd30231,17'd13760,17'd13136,17'd14002,17'd16548,17'd44035,17'd43904,17'd44036,17'd44166,17'd44037,17'd44038,17'd44167,17'd44168,17'd44169,17'd42952,17'd42680,17'd43628,17'd44170,17'd44171,17'd44172,17'd44173,17'd44174,17'd44175,17'd44176,17'd44177,17'd44178,17'd44179,17'd44180,17'd44181,17'd44182,17'd44183,17'd44184,17'd44185,17'd44186,17'd44187,17'd44188,17'd43804,17'd44189,17'd44190,17'd44191,17'd44192,17'd44193,17'd44194,17'd44195,17'd44196,17'd44197,17'd44198,17'd44199,17'd44200,17'd40322,17'd44201,17'd44202,17'd41235,17'd43926,17'd44203,17'd44204,17'd42544,17'd42116,17'd44205,17'd41240,17'd40471,17'd43126,17'd44206,17'd44207,17'd44208,17'd44209,17'd44210,17'd44211,17'd44212,17'd42999,17'd43245,17'd44213,17'd44214,17'd44215,17'd44216,17'd44217,17'd35542,17'd43824,17'd35834,17'd36522,17'd38392,17'd35551,17'd36384,17'd39262,17'd43962,17'd39117,17'd44218,17'd44219,17'd44095,17'd43684,17'd44220,17'd43280,17'd44221,17'd44222,17'd41580,17'd44223,17'd44224,17'd44225,17'd43153,17'd42881,17'd39128,17'd44226,17'd43701,17'd44227,17'd44228,17'd42597,17'd44105,17'd39443,17'd44229,17'd44230,17'd43291,17'd24895,17'd24249,17'd28722,17'd28975,17'd23731,17'd23920,17'd23388,17'd30425,17'd23215,17'd29099,17'd24086,17'd23917,17'd32659,17'd25030,17'd27637,17'd25177,17'd25567,17'd26062,17'd27514,17'd44231,17'd41417,17'd39584,17'd33790,17'd29379,17'd32192,17'd28372,17'd28857,17'd28372,17'd29247,17'd28370,17'd26276,17'd29246,17'd26781,17'd26903,17'd27767,17'd26064,17'd43553,17'd33971,17'd44232,17'd31498,17'd22864,17'd35015,17'd43984,17'd33479,17'd44233,17'd23387,17'd23564,17'd29976,17'd25435,17'd25833,17'd27883,17'd33963,17'd26901,17'd26782,17'd27883,17'd26530,17'd26530,17'd27883,17'd43290,17'd26781,17'd28979,17'd29379,17'd31352,17'd32004,17'd44234,17'd39129,17'd43974,17'd44235,17'd39585,17'd42891,17'd43561,17'd43989,17'd37266,17'd44236,17'd44112,17'd44237,17'd44238,17'd44239,17'd33513,17'd44240,17'd44241,17'd44242,17'd44243,17'd39747,17'd32351,17'd44244,17'd42012,17'd24896,17'd25835,17'd27638,17'd25566,17'd24244,17'd27509,17'd23727,17'd25031,17'd36854,17'd44245,17'd23392,17'd44246,17'd44247,17'd44248,17'd44249,17'd44125,17'd43573,17'd44250,17'd44251,17'd44252,17'd44253,17'd44254,17'd44255,17'd27688,17'd44131,17'd44256,17'd35753,17'd18261,17'd17904,17'd16371,17'd22250,17'd41297,17'd44257,17'd41452,17'd39012,17'd37555,17'd36444,17'd16615,17'd13679,17'd28185,17'd5157,17'd42180,17'd44258,17'd4017,17'd4358,17'd4359,17'd4833,17'd33839,17'd4356,17'd4017,17'd33841,17'd4689,17'd4847,17'd5155,17'd4358,17'd4185,17'd42772,17'd4671,17'd36022,17'd35190,17'd44011,17'd43588,17'd33199,17'd44259,17'd44012,17'd3527,17'd44134,17'd44260,17'd44261,17'd44262,17'd44263,17'd44264,17'd44265,17'd44266,17'd43737,17'd44017,17'd44267,17'd39026,17'd44268,17'd42476,17'd44018,17'd3378,17'd41624,17'd6081,17'd44269,17'd10906,17'd38458,17'd38334,17'd44019,17'd44019,17'd43596,17'd16492,17'd6258,17'd8186,17'd8507,17'd7537,17'd8506,17'd7364,17'd6416,17'd8186,17'd4713,17'd4713,17'd3391,17'd3895,17'd229,17'd3895,17'd5372,17'd2575,17'd951,17'd1382,17'd200,17'd199,17'd1951,17'd1813
},
'{
17'd6420,17'd4892,17'd3902,17'd4425,17'd32728,17'd32728,17'd4244,17'd4245,17'd2422,17'd4247,17'd1416,17'd3905,17'd1128,17'd20404,17'd3905,17'd3905,17'd1128,17'd18,17'd288,17'd981,17'd31,17'd469,17'd2943,17'd2262,17'd1973,17'd1839,17'd1559,17'd1135,17'd16967,17'd827,17'd18275,17'd62,17'd994,17'd2950,17'd43879,17'd44270,17'd3767,17'd15250,17'd44271,17'd18526,17'd16018,17'd44272,17'd44273,17'd44022,17'd18884,17'd12532,17'd12531,17'd12531,17'd10815,17'd42340,17'd17211,17'd44274,17'd43600,17'd15648,17'd38469,17'd44275,17'd44276,17'd44277,17'd41774,17'd40573,17'd43342,17'd40110,17'd39957,17'd42930,17'd39495,17'd44149,17'd44278,17'd44279,17'd44280,17'd34189,17'd44027,17'd12067,17'd10119,17'd7581,17'd6466,17'd11089,17'd43348,17'd6306,17'd5250,17'd7253,17'd42796,17'd44281,17'd43602,17'd6154,17'd44282,17'd6325,17'd43889,17'd44283,17'd43074,17'd42938,17'd44029,17'd44284,17'd44285,17'd42670,17'd41650,17'd44286,17'd43895,17'd7601,17'd44287,17'd44288,17'd44289,17'd44290,17'd44291,17'd44292,17'd44293,17'd44294,17'd30672,17'd15297,17'd8720,17'd10174,17'd14811,17'd14811,17'd15684,17'd9194,17'd17480,17'd10336,17'd9189,17'd9339,17'd9341,17'd9883,17'd11523,17'd29488,17'd28105,17'd30218,17'd35372,17'd28345,17'd28230,17'd28107,17'd24537,17'd23512,17'd23170,17'd22472,17'd18327,17'd11397,17'd11274,17'd11397,17'd18327,17'd21985,17'd21985,17'd18327,17'd23337,17'd11398,17'd11525,17'd11526,17'd11671,17'd9741,17'd9885,17'd10742,17'd9479,17'd11809,17'd10742,17'd10743,17'd9741,17'd11276,17'd12863,17'd12863,17'd10991,17'd11133,17'd26374,17'd10473,17'd10853,17'd15186,17'd29937,17'd34393,17'd33583,17'd32447,17'd32294,17'd30983,17'd13643,17'd14809,17'd15685,17'd12858,17'd15810,17'd43219,17'd44295,17'd44036,17'd44166,17'd44296,17'd44297,17'd44298,17'd44168,17'd44169,17'd44299,17'd42525,17'd44300,17'd44170,17'd44171,17'd44301,17'd44302,17'd35822,17'd44303,17'd44304,17'd44305,17'd44306,17'd44307,17'd44308,17'd44309,17'd44310,17'd44311,17'd44312,17'd44313,17'd44314,17'd44315,17'd40638,17'd44316,17'd44317,17'd41069,17'd41069,17'd44318,17'd44319,17'd44320,17'd44321,17'd44322,17'd44323,17'd44324,17'd44325,17'd44326,17'd43785,17'd44327,17'd43946,17'd41067,17'd44328,17'd44329,17'd44330,17'd44331,17'd41694,17'd40642,17'd44332,17'd44333,17'd44334,17'd44207,17'd44335,17'd44336,17'd44337,17'd44338,17'd44339,17'd44340,17'd44341,17'd44342,17'd44343,17'd44344,17'd44345,17'd34582,17'd38775,17'd44346,17'd44347,17'd33620,17'd33620,17'd38392,17'd35972,17'd38958,17'd38958,17'd43826,17'd38959,17'd44218,17'd44348,17'd44349,17'd44350,17'd40949,17'd44351,17'd44352,17'd44353,17'd42145,17'd44224,17'd44354,17'd44355,17'd43153,17'd43545,17'd43546,17'd44356,17'd44357,17'd43289,17'd44358,17'd42597,17'd43291,17'd39443,17'd42749,17'd44359,17'd43157,17'd24745,17'd23917,17'd24902,17'd24902,17'd31033,17'd23734,17'd32191,17'd32830,17'd22501,17'd35865,17'd23918,17'd31033,17'd32659,17'd24898,17'd27512,17'd25709,17'd27638,17'd26530,17'd26903,17'd42437,17'd42600,17'd38974,17'd36264,17'd33952,17'd33654,17'd28372,17'd28857,17'd28372,17'd29247,17'd28854,17'd26276,17'd28980,17'd33963,17'd27515,17'd28481,17'd30606,17'd39443,17'd36152,17'd39282,17'd34455,17'd21694,17'd32187,17'd42887,17'd44360,17'd31501,17'd23387,17'd24902,17'd25320,17'd28723,17'd25833,17'd27640,17'd26781,17'd28726,17'd33963,17'd33499,17'd27883,17'd26530,17'd27640,17'd43290,17'd26781,17'd28980,17'd33952,17'd31352,17'd32495,17'd44361,17'd39434,17'd44362,17'd44227,17'd33475,17'd42605,17'd43561,17'd43989,17'd37266,17'd44236,17'd44112,17'd44363,17'd42164,17'd33347,17'd25035,17'd25441,17'd44364,17'd44365,17'd44366,17'd33674,17'd23215,17'd23919,17'd24590,17'd24417,17'd34127,17'd25567,17'd28723,17'd24244,17'd27509,17'd23727,17'd25031,17'd36854,17'd44367,17'd44368,17'd44369,17'd44247,17'd44370,17'd44371,17'd44372,17'd43573,17'd44373,17'd44374,17'd41748,17'd44375,17'd44376,17'd44377,17'd21759,17'd44378,17'd44379,17'd36306,17'd18621,17'd16847,17'd16247,17'd39162,17'd40985,17'd44380,17'd22088,17'd41754,17'd37427,17'd36444,17'd16615,17'd13800,17'd5335,17'd4529,17'd33691,17'd40548,17'd41455,17'd33839,17'd4359,17'd4359,17'd33839,17'd4356,17'd4356,17'd33841,17'd4847,17'd37153,17'd5155,17'd4358,17'd4185,17'd4185,17'd4671,17'd42179,17'd44381,17'd4665,17'd43588,17'd33199,17'd44259,17'd44012,17'd33201,17'd44382,17'd44260,17'd44383,17'd44384,17'd44385,17'd44264,17'd44265,17'd39322,17'd41309,17'd44017,17'd44267,17'd44386,17'd44268,17'd42476,17'd42477,17'd42334,17'd3702,17'd7849,17'd39789,17'd39032,17'd38458,17'd38334,17'd44019,17'd44019,17'd44387,17'd37959,17'd6258,17'd6416,17'd7537,17'd7537,17'd8506,17'd8506,17'd8507,17'd7365,17'd4713,17'd4729,17'd3391,17'd3895,17'd229,17'd4880,17'd2409,17'd2575,17'd780,17'd11445,17'd1103,17'd198,17'd1951,17'd1813
},
'{
17'd4428,17'd4892,17'd3902,17'd5646,17'd44388,17'd35063,17'd4892,17'd4245,17'd2422,17'd4247,17'd1416,17'd3905,17'd20404,17'd20404,17'd3905,17'd3905,17'd980,17'd980,17'd28,17'd29,17'd30,17'd1129,17'd2940,17'd2602,17'd2266,17'd19608,17'd1703,17'd19499,17'd16967,17'd827,17'd18275,17'd993,17'd1287,17'd1146,17'd43879,17'd37577,17'd44389,17'd15250,17'd44271,17'd18526,17'd44390,17'd44272,17'd44273,17'd44022,17'd18884,17'd11764,17'd12532,17'd12531,17'd10815,17'd21487,17'd20430,17'd16990,17'd42045,17'd44391,17'd44392,17'd39800,17'd44393,17'd44394,17'd40725,17'd40419,17'd40110,17'd39496,17'd41014,17'd41488,17'd39337,17'd39800,17'd44395,17'd44279,17'd42791,17'd44396,17'd44027,17'd12067,17'd10119,17'd7579,17'd7251,17'd6626,17'd44153,17'd6627,17'd5250,17'd7253,17'd42796,17'd44281,17'd43602,17'd43887,17'd44397,17'd44155,17'd44156,17'd44283,17'd43074,17'd42936,17'd43891,17'd43892,17'd43355,17'd44398,17'd41650,17'd44399,17'd44400,17'd44401,17'd44402,17'd44403,17'd44404,17'd44405,17'd44406,17'd44407,17'd44293,17'd44408,17'd36932,17'd9348,17'd8720,17'd10174,17'd15944,17'd15944,17'd15684,17'd9194,17'd17480,17'd8874,17'd9192,17'd9338,17'd9472,17'd10166,17'd14673,17'd24995,17'd25927,17'd28816,17'd28460,17'd28345,17'd28230,17'd28107,17'd24537,17'd24030,17'd21505,17'd16442,17'd18327,17'd11397,17'd11397,17'd11397,17'd18327,17'd21985,17'd24994,17'd18327,17'd23337,17'd25280,17'd12423,17'd19280,17'd11671,17'd9741,17'd9885,17'd10992,17'd10742,17'd17011,17'd10742,17'd10743,17'd9885,17'd11276,17'd12863,17'd12863,17'd10991,17'd11133,17'd10165,17'd27743,17'd25144,17'd11665,17'd40286,17'd44409,17'd33583,17'd33885,17'd31449,17'd38368,17'd30378,17'd13760,17'd13519,17'd12858,17'd11665,17'd43364,17'd44295,17'd44410,17'd44411,17'd40751,17'd44412,17'd44413,17'd44414,17'd41939,17'd44415,17'd42369,17'd44416,17'd44417,17'd44418,17'd44419,17'd44420,17'd44421,17'd44422,17'd44423,17'd44424,17'd44425,17'd44426,17'd44427,17'd44428,17'd44429,17'd44430,17'd44431,17'd44432,17'd44433,17'd44434,17'd41549,17'd43803,17'd41954,17'd44057,17'd44435,17'd43501,17'd43235,17'd44436,17'd44437,17'd44438,17'd44439,17'd44440,17'd44441,17'd44442,17'd44443,17'd44444,17'd44445,17'd44446,17'd43501,17'd41816,17'd44447,17'd41699,17'd44448,17'd44449,17'd44450,17'd44334,17'd44451,17'd44452,17'd44053,17'd44453,17'd44454,17'd44455,17'd44456,17'd44457,17'd44458,17'd44459,17'd44460,17'd44461,17'd44462,17'd44463,17'd44464,17'd44465,17'd36674,17'd35273,17'd36247,17'd36245,17'd35972,17'd38958,17'd39567,17'd42868,17'd44466,17'd44467,17'd44468,17'd44095,17'd44350,17'd44469,17'd44351,17'd44470,17'd44471,17'd42880,17'd44472,17'd44473,17'd44355,17'd42881,17'd44474,17'd44475,17'd44476,17'd44357,17'd42298,17'd44477,17'd42597,17'd44105,17'd39591,17'd29970,17'd44229,17'd38282,17'd24745,17'd34467,17'd24902,17'd24902,17'd29241,17'd31190,17'd23217,17'd33316,17'd22501,17'd35865,17'd23565,17'd31033,17'd23916,17'd24898,17'd27512,17'd28597,17'd30606,17'd27515,17'd28978,17'd44478,17'd43433,17'd41109,17'd35570,17'd29977,17'd32017,17'd28372,17'd28857,17'd28372,17'd29104,17'd32354,17'd29977,17'd28980,17'd33963,17'd27515,17'd30606,17'd27638,17'd31034,17'd23923,17'd36009,17'd33649,17'd31831,17'd22510,17'd43158,17'd40523,17'd31195,17'd29827,17'd30879,17'd29244,17'd28723,17'd25707,17'd27371,17'd26781,17'd28486,17'd26782,17'd43290,17'd27640,17'd27883,17'd27640,17'd43290,17'd34767,17'd28980,17'd33952,17'd31352,17'd32495,17'd41863,17'd44479,17'd39434,17'd44227,17'd33475,17'd42605,17'd44480,17'd44481,17'd33669,17'd44236,17'd31046,17'd44482,17'd44483,17'd44484,17'd44485,17'd44486,17'd44487,17'd44488,17'd25182,17'd44489,17'd23389,17'd44490,17'd23382,17'd24743,17'd25320,17'd28597,17'd25435,17'd27026,17'd23726,17'd23727,17'd25031,17'd37267,17'd23738,17'd44491,17'd44492,17'd44247,17'd33676,17'd44493,17'd44494,17'd44495,17'd43574,17'd44496,17'd44497,17'd44498,17'd42172,17'd44499,17'd44500,17'd44501,17'd44502,17'd44503,17'd18023,17'd15340,17'd18134,17'd39012,17'd44504,17'd44505,17'd44504,17'd37555,17'd22767,17'd41141,17'd12906,17'd15990,17'd5160,17'd4529,17'd39468,17'd42464,17'd39313,17'd39468,17'd4833,17'd4359,17'd4357,17'd4831,17'd4356,17'd33841,17'd4689,17'd4847,17'd4526,17'd4358,17'd4185,17'd4830,17'd36022,17'd42773,17'd35188,17'd42774,17'd44506,17'd33199,17'd44259,17'd44012,17'd44507,17'd44508,17'd44509,17'd44510,17'd40091,17'd39320,17'd44511,17'd44512,17'd39322,17'd41154,17'd36743,17'd44267,17'd44386,17'd44268,17'd44513,17'd44514,17'd42334,17'd3702,17'd5493,17'd39789,17'd39032,17'd38458,17'd38334,17'd44019,17'd12913,17'd44387,17'd37959,17'd6258,17'd6094,17'd7537,17'd7537,17'd8506,17'd6418,17'd6416,17'd7365,17'd4713,17'd4729,17'd3391,17'd3895,17'd4881,17'd4880,17'd2409,17'd2575,17'd413,17'd1526,17'd44020,17'd198,17'd1951,17'd14587
},
'{
17'd4428,17'd3903,17'd4087,17'd5646,17'd44388,17'd32728,17'd4244,17'd4245,17'd2422,17'd4247,17'd1416,17'd3905,17'd20404,17'd20404,17'd3905,17'd3905,17'd980,17'd28,17'd288,17'd981,17'd31,17'd469,17'd2943,17'd2262,17'd1973,17'd1839,17'd1559,17'd19499,17'd16967,17'd992,17'd828,17'd16637,17'd2612,17'd1146,17'd43879,17'd37577,17'd36184,17'd20416,17'd44515,17'd44516,17'd44390,17'd44272,17'd44273,17'd44517,17'd12532,17'd11764,17'd12532,17'd12531,17'd10815,17'd21487,17'd20588,17'd16990,17'd44144,17'd43600,17'd15648,17'd42047,17'd44518,17'd44519,17'd42488,17'd40111,17'd43750,17'd40722,17'd39496,17'd43465,17'd39337,17'd39800,17'd44395,17'd44520,17'd42791,17'd44396,17'd44027,17'd12067,17'd10119,17'd7581,17'd6466,17'd5253,17'd6306,17'd4610,17'd44521,17'd7090,17'd6474,17'd44281,17'd43602,17'd6154,17'd44282,17'd6325,17'd42665,17'd44283,17'd44522,17'd42938,17'd44029,17'd44284,17'd44285,17'd44523,17'd44524,17'd44525,17'd44526,17'd44401,17'd44527,17'd44528,17'd44529,17'd44530,17'd44531,17'd44532,17'd44533,17'd44165,17'd23341,17'd9348,17'd8873,17'd10173,17'd15807,17'd15807,17'd17480,17'd9194,17'd17480,17'd10336,17'd9189,17'd9339,17'd9341,17'd10329,17'd11523,17'd29488,17'd28105,17'd29778,17'd28460,17'd28818,17'd28230,17'd28107,17'd24537,17'd24030,17'd21505,17'd16442,17'd18327,17'd11397,17'd11397,17'd11396,17'd18327,17'd18327,17'd23169,17'd23169,17'd14382,17'd23337,17'd28821,17'd13647,17'd17847,17'd9884,17'd9885,17'd10992,17'd10742,17'd17011,17'd10742,17'd10743,17'd10992,17'd11671,17'd11670,17'd12863,17'd10991,17'd11133,17'd10165,17'd19281,17'd14263,17'd29341,17'd39514,17'd44409,17'd32608,17'd32447,17'd32294,17'd29205,17'd14523,17'd12418,17'd12106,17'd13135,17'd11519,17'd14926,17'd44295,17'd44534,17'd44535,17'd42813,17'd43365,17'd44168,17'd44536,17'd41939,17'd44537,17'd44538,17'd44539,17'd44540,17'd44418,17'd44541,17'd44542,17'd44543,17'd44544,17'd44545,17'd44546,17'd44547,17'd44548,17'd44549,17'd44550,17'd44551,17'd44552,17'd44553,17'd44554,17'd44555,17'd44556,17'd40787,17'd40479,17'd44188,17'd41384,17'd43946,17'd42251,17'd41229,17'd44327,17'd44557,17'd44558,17'd44559,17'd44560,17'd44561,17'd44562,17'd44443,17'd43944,17'd44563,17'd41374,17'd41071,17'd42543,17'd44564,17'd44565,17'd44332,17'd40646,17'd44566,17'd43239,17'd40168,17'd44567,17'd44568,17'd44569,17'd44570,17'd44571,17'd43673,17'd44572,17'd44573,17'd44574,17'd44214,17'd44575,17'd44576,17'd44577,17'd44578,17'd34076,17'd36825,17'd36247,17'd33620,17'd38645,17'd36385,17'd38958,17'd39568,17'd44579,17'd44580,17'd44467,17'd44581,17'd43966,17'd44582,17'd44583,17'd44351,17'd44584,17'd44585,17'd43423,17'd44586,17'd44587,17'd44355,17'd44588,17'd43832,17'd39903,17'd43974,17'd44234,17'd42298,17'd41418,17'd44589,17'd43694,17'd29825,17'd29970,17'd42749,17'd43553,17'd24745,17'd23916,17'd24902,17'd30275,17'd29241,17'd38980,17'd41273,17'd41272,17'd30277,17'd35865,17'd23565,17'd24086,17'd23916,17'd24898,17'd27512,17'd28597,17'd30606,17'd27515,17'd31827,17'd44590,17'd42740,17'd37114,17'd35707,17'd30279,17'd32355,17'd28372,17'd28728,17'd28371,17'd29104,17'd33319,17'd29977,17'd28980,17'd26782,17'd26174,17'd30606,17'd28598,17'd29103,17'd23387,17'd22857,17'd32013,17'd32997,17'd22864,17'd32012,17'd44591,17'd31195,17'd29827,17'd29100,17'd25438,17'd25566,17'd26903,17'd27371,17'd26901,17'd28979,17'd26781,17'd27371,17'd27259,17'd27640,17'd27640,17'd43290,17'd34767,17'd28980,17'd29977,17'd31352,17'd42598,17'd41997,17'd44592,17'd44593,17'd44103,17'd44594,17'd42605,17'd44480,17'd44481,17'd41424,17'd44236,17'd37121,17'd44595,17'd44596,17'd44597,17'd44598,17'd44599,17'd44600,17'd44601,17'd44602,17'd33972,17'd37533,17'd31190,17'd44603,17'd34884,17'd29976,17'd27882,17'd28600,17'd25173,17'd24245,17'd23559,17'd25031,17'd29688,17'd36152,17'd38296,17'd44604,17'd44247,17'd38686,17'd25956,17'd44605,17'd44606,17'd44607,17'd44608,17'd44609,17'd44498,17'd42172,17'd44499,17'd21447,17'd44501,17'd44610,17'd44611,17'd27198,17'd24803,17'd19590,17'd41754,17'd38844,17'd44612,17'd38844,17'd37555,17'd22943,17'd36310,17'd13046,17'd44613,17'd5329,17'd44614,17'd39468,17'd42464,17'd40395,17'd4356,17'd4833,17'd4359,17'd4515,17'd4356,17'd4356,17'd33841,17'd4847,17'd37153,17'd5155,17'd4358,17'd4185,17'd4830,17'd36022,17'd36166,17'd34327,17'd42774,17'd44506,17'd33199,17'd44259,17'd44012,17'd4350,17'd44508,17'd44509,17'd44510,17'd40091,17'd39320,17'd44615,17'd44512,17'd39322,17'd41154,17'd36743,17'd44267,17'd44386,17'd44268,17'd42476,17'd42477,17'd42334,17'd41905,17'd5493,17'd39789,17'd39032,17'd38458,17'd38334,17'd44019,17'd12913,17'd38581,17'd44387,17'd16492,17'd6094,17'd7537,17'd7364,17'd44616,17'd15484,17'd6094,17'd7365,17'd4713,17'd4729,17'd3391,17'd3895,17'd4881,17'd4880,17'd2409,17'd2575,17'd413,17'd939,17'd1103,17'd198,17'd1951,17'd14587
},
'{
17'd4088,17'd4892,17'd3902,17'd4426,17'd44617,17'd44388,17'd4244,17'd4245,17'd2422,17'd4247,17'd1416,17'd3905,17'd20404,17'd20404,17'd3905,17'd3905,17'd652,17'd652,17'd288,17'd29,17'd30,17'd1129,17'd2940,17'd3253,17'd2263,17'd19874,17'd1423,17'd1135,17'd1138,17'd992,17'd667,17'd828,17'd1141,17'd3264,17'd2953,17'd37577,17'd44618,17'd44619,17'd44620,17'd28436,17'd44390,17'd31418,17'd44273,17'd44621,17'd16658,17'd11913,17'd11913,17'd11913,17'd12531,17'd19756,17'd20429,17'd17211,17'd14480,17'd44144,17'd44622,17'd42047,17'd44623,17'd44624,17'd41169,17'd40110,17'd39337,17'd40570,17'd43465,17'd43343,17'd42048,17'd44625,17'd44626,17'd44627,17'd42791,17'd42659,17'd44628,17'd21190,17'd7579,17'd7579,17'd44629,17'd44630,17'd44153,17'd6627,17'd4924,17'd7253,17'd42796,17'd6313,17'd43602,17'd42663,17'd42211,17'd44631,17'd44632,17'd44283,17'd42938,17'd43206,17'd44029,17'd44633,17'd44285,17'd44634,17'd44635,17'd44636,17'd44637,17'd44638,17'd44639,17'd44640,17'd44641,17'd44642,17'd44643,17'd44644,17'd44645,17'd44408,17'd44646,17'd9348,17'd9043,17'd9346,17'd15807,17'd10173,17'd10336,17'd15684,17'd14811,17'd8874,17'd9192,17'd20175,17'd21820,17'd10165,17'd11274,17'd15055,17'd24856,17'd28343,17'd28460,17'd28104,17'd27121,17'd24991,17'd24537,17'd23512,17'd21505,17'd16442,17'd18327,17'd11396,17'd11522,17'd11396,17'd17478,17'd23513,17'd23513,17'd23513,17'd14382,17'd12583,17'd11668,17'd11525,17'd10331,17'd10024,17'd9885,17'd9885,17'd10742,17'd17011,17'd17011,17'd9341,17'd9885,17'd12116,17'd10479,17'd12863,17'd14518,17'd10991,17'd10326,17'd10166,17'd10474,17'd29341,17'd39514,17'd33250,17'd33583,17'd33735,17'd30085,17'd29791,17'd44647,17'd13518,17'd13136,17'd12260,17'd11665,17'd29073,17'd44648,17'd44534,17'd42812,17'd44649,17'd44650,17'd44414,17'd41940,17'd41940,17'd44651,17'd44651,17'd41353,17'd44418,17'd44652,17'd44653,17'd44654,17'd44655,17'd44656,17'd44657,17'd44658,17'd44659,17'd44660,17'd44661,17'd44662,17'd44663,17'd44664,17'd44665,17'd44666,17'd44667,17'd44668,17'd44669,17'd40785,17'd44670,17'd41538,17'd41072,17'd41682,17'd41071,17'd41375,17'd43946,17'd41066,17'd41067,17'd43945,17'd44317,17'd44317,17'd44671,17'd41228,17'd41954,17'd41377,17'd42406,17'd44672,17'd44673,17'd40644,17'd44674,17'd44675,17'd40488,17'd44676,17'd44677,17'd44678,17'd44679,17'd44680,17'd44681,17'd40021,17'd44682,17'd44683,17'd44684,17'd44685,17'd39995,17'd44686,17'd44687,17'd44688,17'd44689,17'd41716,17'd38134,17'd38263,17'd44690,17'd38645,17'd35971,17'd38958,17'd39415,17'd39416,17'd44691,17'd44692,17'd44693,17'd44694,17'd43010,17'd44695,17'd43010,17'd43142,17'd44696,17'd43151,17'd44587,17'd44473,17'd44101,17'd44355,17'd44697,17'd44226,17'd44698,17'd44234,17'd42436,17'd41418,17'd44699,17'd43836,17'd38156,17'd28484,17'd27511,17'd31034,17'd25032,17'd24252,17'd28722,17'd24086,17'd33950,17'd41587,17'd33316,17'd33799,17'd23215,17'd29829,17'd31502,17'd24086,17'd34467,17'd25030,17'd25177,17'd28598,17'd26062,17'd28724,17'd28978,17'd44700,17'd42740,17'd34450,17'd31354,17'd29977,17'd32355,17'd29248,17'd29248,17'd32017,17'd33654,17'd32354,17'd37513,17'd34767,17'd26782,17'd26174,17'd28598,17'd25567,17'd33483,17'd35865,17'd22857,17'd35292,17'd44701,17'd34457,17'd32012,17'd44702,17'd24592,17'd29099,17'd24090,17'd27511,17'd25708,17'd26903,17'd27371,17'd28726,17'd28727,17'd26901,17'd27371,17'd27259,17'd27640,17'd33815,17'd43290,17'd44703,17'd44704,17'd29977,17'd38025,17'd41271,17'd43974,17'd44705,17'd39583,17'd44103,17'd33475,17'd35707,17'd31503,17'd30586,17'd41424,17'd44236,17'd44706,17'd43166,17'd44707,17'd44708,17'd44709,17'd44599,17'd44710,17'd44711,17'd44712,17'd44713,17'd32015,17'd38980,17'd23210,17'd24090,17'd25180,17'd28717,17'd25317,17'd44714,17'd24245,17'd25030,17'd25032,17'd34883,17'd44715,17'd44716,17'd44717,17'd44718,17'd33676,17'd44719,17'd44720,17'd44721,17'd44722,17'd44723,17'd44609,17'd44724,17'd42316,17'd44725,17'd21447,17'd44726,17'd44610,17'd44611,17'd24802,17'd17655,17'd16955,17'd37555,17'd39012,17'd44727,17'd44504,17'd22767,17'd36029,17'd38701,17'd13046,17'd29296,17'd5334,17'd5000,17'd41458,17'd39313,17'd44728,17'd41612,17'd4357,17'd4833,17'd4017,17'd4016,17'd4356,17'd33841,17'd4689,17'd4684,17'd4526,17'd4833,17'd42772,17'd42630,17'd42179,17'd35332,17'd44729,17'd42774,17'd44730,17'd33199,17'd44259,17'd44731,17'd44507,17'd44732,17'd44733,17'd44734,17'd40406,17'd44735,17'd44736,17'd41899,17'd44737,17'd44738,17'd44739,17'd44267,17'd44386,17'd44740,17'd44741,17'd2533,17'd43740,17'd41480,17'd5493,17'd39789,17'd39032,17'd44742,17'd41481,17'd44019,17'd38580,17'd43330,17'd44387,17'd16623,17'd6890,17'd7537,17'd7537,17'd7364,17'd6418,17'd8186,17'd4869,17'd4729,17'd4713,17'd4085,17'd3895,17'd4880,17'd5371,17'd2409,17'd412,17'd413,17'd1669,17'd43878,17'd196,17'd1530,17'd14587
},
'{
17'd4088,17'd4244,17'd4087,17'd5646,17'd44617,17'd44388,17'd4244,17'd4245,17'd2422,17'd4247,17'd1416,17'd3905,17'd20404,17'd20404,17'd3905,17'd3905,17'd652,17'd652,17'd288,17'd981,17'd31,17'd469,17'd2943,17'd2262,17'd2122,17'd1972,17'd1557,17'd1135,17'd16967,17'd992,17'd667,17'd828,17'd1142,17'd3264,17'd2953,17'd37577,17'd44618,17'd44619,17'd44743,17'd28436,17'd44390,17'd44744,17'd44745,17'd44621,17'd16658,17'd11913,17'd11913,17'd11913,17'd12532,17'd19388,17'd44746,17'd17450,17'd17099,17'd16990,17'd15014,17'd44747,17'd44748,17'd44749,17'd44750,17'd39801,17'd39191,17'd44751,17'd40570,17'd39337,17'd38879,17'd44625,17'd44626,17'd44752,17'd44753,17'd44754,17'd44755,17'd21190,17'd8685,17'd7411,17'd6140,17'd5254,17'd6306,17'd6627,17'd4924,17'd7253,17'd42796,17'd6313,17'd43602,17'd6154,17'd44282,17'd44756,17'd44757,17'd44758,17'd42938,17'd43472,17'd44759,17'd44760,17'd41787,17'd44761,17'd44762,17'd44763,17'd44764,17'd44765,17'd44766,17'd34951,17'd44767,17'd44768,17'd44769,17'd44532,17'd44770,17'd44771,17'd35930,17'd9040,17'd9043,17'd9346,17'd10334,17'd15807,17'd10175,17'd9194,17'd17480,17'd10336,17'd9189,17'd9191,17'd10744,17'd10330,17'd25280,17'd29488,17'd26371,17'd28343,17'd28460,17'd28104,17'd27121,17'd24991,17'd24537,17'd23515,17'd21505,17'd22472,17'd18327,17'd11396,17'd11522,17'd18327,17'd23513,17'd23167,17'd23167,17'd23513,17'd36348,17'd44772,17'd18326,17'd12423,17'd29335,17'd13522,17'd10169,17'd9741,17'd10742,17'd17011,17'd17011,17'd9341,17'd9885,17'd12116,17'd10479,17'd12863,17'd10991,17'd10991,17'd10326,17'd19281,17'd14132,17'd10736,17'd40137,17'd33250,17'd32608,17'd33416,17'd29936,17'd29205,17'd16799,17'd13252,17'd11958,17'd12996,17'd11519,17'd44773,17'd44648,17'd44774,17'd44775,17'd44649,17'd44776,17'd44414,17'd41940,17'd42527,17'd44651,17'd44651,17'd41352,17'd42081,17'd44777,17'd44778,17'd44779,17'd44780,17'd38123,17'd44781,17'd44782,17'd44783,17'd44784,17'd44785,17'd44786,17'd44787,17'd42725,17'd44788,17'd43953,17'd44789,17'd44790,17'd44791,17'd42120,17'd42408,17'd42099,17'd44792,17'd44793,17'd44331,17'd40635,17'd41547,17'd41225,17'd41373,17'd41384,17'd41817,17'd44794,17'd43924,17'd40915,17'd44795,17'd44796,17'd44797,17'd44798,17'd44799,17'd44800,17'd42122,17'd44801,17'd44451,17'd44802,17'd44803,17'd44804,17'd44805,17'd44806,17'd44807,17'd44808,17'd44809,17'd44810,17'd44811,17'd44812,17'd43133,17'd33911,17'd44813,17'd34420,17'd37637,17'd35972,17'd38009,17'd38389,17'd44690,17'd35972,17'd36384,17'd39567,17'd39416,17'd38006,17'd44814,17'd44467,17'd44815,17'd44816,17'd43010,17'd44817,17'd44818,17'd44819,17'd44820,17'd43151,17'd44472,17'd44473,17'd44821,17'd44821,17'd39128,17'd44356,17'd44822,17'd43434,17'd42298,17'd43548,17'd44106,17'd44229,17'd43977,17'd25317,17'd25438,17'd29244,17'd25032,17'd24252,17'd28975,17'd23732,17'd33794,17'd37116,17'd31495,17'd31495,17'd32351,17'd23388,17'd29376,17'd24086,17'd24252,17'd24898,17'd33484,17'd30734,17'd26530,17'd28853,17'd27260,17'd44823,17'd43434,17'd41110,17'd27885,17'd30279,17'd33165,17'd32355,17'd29248,17'd32017,17'd32192,17'd32354,17'd37513,17'd34767,17'd28725,17'd25565,17'd25567,17'd28597,17'd30432,17'd29530,17'd23573,17'd22683,17'd44824,17'd34457,17'd44825,17'd34453,17'd33673,17'd23565,17'd24415,17'd27511,17'd25708,17'd26903,17'd27371,17'd28726,17'd28980,17'd28726,17'd35023,17'd27371,17'd27640,17'd33815,17'd43290,17'd44703,17'd44826,17'd29977,17'd37908,17'd44827,17'd39434,17'd44828,17'd39738,17'd44103,17'd33475,17'd35570,17'd31503,17'd30586,17'd41424,17'd31681,17'd29994,17'd42610,17'd38419,17'd44829,17'd39756,17'd44830,17'd44831,17'd44832,17'd44833,17'd44834,17'd44835,17'd31341,17'd23210,17'd29100,17'd24895,17'd25177,17'd25317,17'd27510,17'd23727,17'd25030,17'd24895,17'd34883,17'd29829,17'd32346,17'd44836,17'd44837,17'd38686,17'd44838,17'd44839,17'd44840,17'd44722,17'd44841,17'd44842,17'd44843,17'd42316,17'd44844,17'd21447,17'd44726,17'd44845,17'd44846,17'd29297,17'd15094,17'd26710,17'd37427,17'd41754,17'd44504,17'd39012,17'd36734,17'd36170,17'd36171,17'd13046,17'd30179,17'd5334,17'd5000,17'd4356,17'd42772,17'd44728,17'd41612,17'd4357,17'd4833,17'd4357,17'd4831,17'd4356,17'd33841,17'd5156,17'd4684,17'd4526,17'd4833,17'd4185,17'd42630,17'd42179,17'd4669,17'd44729,17'd42774,17'd44730,17'd33199,17'd44259,17'd44012,17'd33201,17'd44732,17'd44509,17'd44734,17'd40406,17'd44735,17'd44615,17'd44847,17'd44737,17'd44738,17'd44848,17'd44267,17'd44386,17'd44740,17'd44849,17'd42784,17'd43740,17'd41905,17'd41907,17'd18629,17'd39181,17'd38859,17'd41481,17'd44019,17'd38580,17'd43330,17'd44387,17'd16623,17'd6094,17'd7537,17'd7364,17'd44850,17'd15484,17'd6258,17'd4869,17'd4729,17'd4713,17'd4085,17'd3895,17'd4880,17'd5371,17'd412,17'd412,17'd1383,17'd421,17'd43878,17'd196,17'd1530,17'd1811
},
'{
17'd4428,17'd4892,17'd3902,17'd5646,17'd44617,17'd44388,17'd4244,17'd4245,17'd2422,17'd4247,17'd1416,17'd3905,17'd20404,17'd20404,17'd3905,17'd3905,17'd980,17'd652,17'd29,17'd29,17'd30,17'd1129,17'd16866,17'd3253,17'd2263,17'd19874,17'd1423,17'd1559,17'd44851,17'd16967,17'd826,17'd828,17'd1142,17'd3264,17'd44852,17'd37577,17'd36184,17'd44619,17'd44743,17'd44853,17'd44854,17'd44744,17'd44855,17'd44621,17'd16765,17'd12361,17'd11913,17'd11913,17'd12532,17'd19513,17'd21039,17'd35354,17'd20431,17'd37177,17'd16524,17'd44856,17'd44857,17'd44023,17'd44145,17'd39494,17'd44858,17'd44859,17'd44751,17'd44751,17'd44859,17'd41631,17'd37315,17'd44860,17'd44861,17'd44862,17'd44628,17'd12816,17'd8685,17'd7579,17'd7417,17'd11479,17'd5254,17'd6627,17'd5250,17'd4923,17'd7754,17'd6314,17'd44863,17'd42663,17'd42211,17'd44756,17'd42665,17'd44864,17'd42938,17'd43206,17'd44029,17'd44760,17'd44865,17'd44761,17'd44762,17'd44763,17'd44866,17'd44867,17'd44868,17'd44869,17'd44870,17'd44871,17'd44872,17'd44873,17'd44645,17'd44874,17'd44646,17'd9040,17'd9043,17'd10335,17'd9480,17'd15807,17'd10175,17'd10175,17'd17480,17'd9189,17'd9191,17'd20175,17'd44875,17'd10165,17'd11274,17'd24995,17'd24856,17'd28816,17'd28460,17'd28104,17'd25528,17'd18200,17'd24537,17'd23515,17'd23170,17'd21361,17'd18327,17'd18327,17'd17478,17'd17478,17'd18443,17'd16325,17'd21361,17'd18443,17'd23513,17'd17478,17'd23337,17'd11668,17'd19280,17'd19278,17'd10024,17'd9741,17'd10742,17'd17011,17'd10742,17'd9341,17'd10992,17'd12116,17'd11134,17'd11528,17'd10991,17'd10991,17'd10326,17'd10166,17'd10474,17'd18445,17'd34709,17'd33250,17'd32608,17'd33885,17'd30085,17'd29791,17'd44647,17'd21506,17'd13519,17'd12114,17'd11665,17'd44773,17'd44648,17'd44774,17'd44775,17'd44876,17'd42679,17'd41798,17'd44877,17'd42527,17'd44651,17'd44651,17'd44878,17'd42081,17'd44777,17'd44879,17'd44880,17'd44881,17'd44882,17'd44883,17'd44306,17'd44884,17'd41086,17'd44885,17'd44886,17'd44887,17'd44808,17'd44888,17'd44889,17'd43814,17'd44890,17'd44891,17'd44892,17'd44893,17'd44894,17'd44895,17'd42119,17'd44896,17'd44897,17'd44898,17'd44795,17'd41698,17'd40777,17'd40777,17'd40923,17'd44899,17'd44898,17'd44900,17'd44901,17'd41240,17'd44902,17'd44903,17'd44904,17'd44905,17'd44906,17'd44907,17'd44908,17'd44568,17'd44909,17'd44910,17'd42724,17'd44911,17'd44912,17'd44913,17'd44914,17'd44915,17'd44916,17'd44917,17'd44918,17'd44919,17'd44920,17'd44921,17'd35972,17'd38009,17'd38645,17'd36245,17'd35972,17'd36384,17'd39567,17'd39415,17'd44922,17'd44923,17'd44924,17'd44925,17'd44926,17'd44927,17'd44817,17'd44350,17'd44928,17'd44929,17'd44930,17'd44472,17'd44931,17'd44931,17'd44932,17'd43833,17'd44356,17'd44933,17'd44227,17'd43289,17'd44934,17'd44230,17'd38156,17'd39591,17'd29101,17'd25320,17'd25180,17'd25032,17'd24252,17'd28852,17'd23732,17'd31190,17'd22328,17'd39911,17'd31495,17'd22501,17'd30128,17'd29827,17'd30879,17'd24416,17'd24897,17'd33484,17'd27767,17'd27640,17'd27146,17'd43551,17'd44935,17'd44234,17'd41731,17'd27885,17'd32832,17'd33165,17'd32017,17'd32355,17'd33654,17'd32192,17'd33319,17'd29246,17'd26781,17'd28853,17'd28483,17'd28369,17'd25709,17'd25031,17'd23387,17'd23573,17'd22683,17'd21847,17'd31660,17'd44825,17'd24094,17'd33673,17'd23565,17'd23916,17'd27511,17'd25708,17'd27259,17'd35023,17'd28726,17'd28727,17'd26901,17'd26782,17'd27259,17'd27640,17'd26530,17'd43290,17'd44703,17'd37513,17'd29977,17'd37908,17'd44700,17'd44479,17'd44936,17'd44937,17'd44938,17'd33475,17'd35570,17'd31503,17'd30586,17'd26174,17'd33008,17'd37122,17'd24422,17'd43854,17'd44939,17'd44940,17'd44941,17'd42165,17'd44942,17'd24256,17'd44943,17'd44944,17'd31828,17'd23918,17'd28975,17'd24745,17'd25320,17'd28850,17'd26399,17'd24740,17'd24895,17'd30126,17'd44945,17'd29829,17'd32013,17'd44946,17'd44947,17'd38552,17'd44948,17'd44949,17'd44950,17'd44722,17'd44951,17'd44952,17'd44953,17'd44954,17'd24126,17'd21447,17'd44726,17'd44845,17'd44955,17'd24945,17'd14971,17'd26585,17'd22767,17'd37555,17'd38314,17'd37802,17'd36029,17'd36444,17'd38440,17'd12905,17'd35194,17'd5334,17'd5001,17'd4017,17'd4185,17'd44728,17'd41455,17'd4357,17'd4362,17'd4357,17'd4831,17'd41612,17'd33992,17'd5156,17'd4684,17'd4526,17'd4359,17'd4185,17'd42630,17'd4670,17'd5475,17'd44956,17'd42774,17'd44957,17'd44958,17'd33200,17'd44012,17'd33201,17'd44732,17'd44959,17'd44960,17'd40091,17'd44961,17'd44511,17'd40711,17'd44962,17'd44963,17'd3194,17'd22095,17'd44964,17'd43056,17'd44965,17'd2535,17'd43740,17'd3702,17'd7849,17'd39789,17'd39032,17'd11867,17'd41481,17'd12635,17'd44966,17'd43330,17'd44387,17'd16623,17'd6094,17'd7537,17'd7537,17'd7364,17'd6418,17'd8186,17'd4869,17'd4713,17'd4713,17'd4729,17'd5193,17'd4880,17'd5372,17'd2393,17'd14178,17'd779,17'd421,17'd43878,17'd196,17'd946,17'd196
},
'{
17'd4428,17'd3902,17'd4087,17'd5646,17'd44617,17'd44388,17'd4244,17'd4245,17'd2422,17'd4247,17'd1416,17'd3905,17'd20404,17'd20404,17'd3905,17'd3905,17'd980,17'd652,17'd29,17'd981,17'd31,17'd982,17'd3253,17'd2262,17'd2122,17'd1972,17'd1557,17'd1135,17'd991,17'd992,17'd667,17'd829,17'd1142,17'd3264,17'd44852,17'd37577,17'd36184,17'd44619,17'd44743,17'd44853,17'd44854,17'd44744,17'd44855,17'd44621,17'd16765,17'd12362,17'd11913,17'd11913,17'd12532,17'd19755,17'd21652,17'd18299,17'd20429,17'd20429,17'd41486,17'd38877,17'd40417,17'd44967,17'd44968,17'd44859,17'd38595,17'd42047,17'd44275,17'd38879,17'd39800,17'd42203,17'd44969,17'd44970,17'd44971,17'd44972,17'd44973,17'd12816,17'd7579,17'd7411,17'd6140,17'd5254,17'd6627,17'd5088,17'd5250,17'd7253,17'd42796,17'd6313,17'd43470,17'd6154,17'd44282,17'd44756,17'd42665,17'd44864,17'd43608,17'd43472,17'd44759,17'd44760,17'd44865,17'd44761,17'd44974,17'd44763,17'd44975,17'd44976,17'd44977,17'd44869,17'd44870,17'd44978,17'd44872,17'd44979,17'd44645,17'd44980,17'd44981,17'd9195,17'd9042,17'd10335,17'd9480,17'd10334,17'd16682,17'd10175,17'd17480,17'd10175,17'd9190,17'd15295,17'd13255,17'd10330,17'd25280,17'd29488,17'd26371,17'd28816,17'd28460,17'd28104,17'd24991,17'd18200,17'd24537,17'd23515,17'd23170,17'd21361,17'd23169,17'd18327,17'd14264,17'd14264,17'd18443,17'd22992,17'd22992,17'd14258,17'd44982,17'd23167,17'd14382,17'd43622,17'd19919,17'd17847,17'd9884,17'd10024,17'd9885,17'd10742,17'd10742,17'd10743,17'd10992,17'd9741,17'd11134,17'd11528,17'd10991,17'd10991,17'd11133,17'd10166,17'd10473,17'd10737,17'd17837,17'd33250,17'd32608,17'd32447,17'd29936,17'd44983,17'd29204,17'd21506,17'd13519,17'd12114,17'd29341,17'd28697,17'd44648,17'd44984,17'd44985,17'd44876,17'd42524,17'd41798,17'd44418,17'd44877,17'd44651,17'd44651,17'd44878,17'd44418,17'd44652,17'd44986,17'd44987,17'd44988,17'd44989,17'd44990,17'd44991,17'd44992,17'd44993,17'd44885,17'd44994,17'd44995,17'd39544,17'd41084,17'd44996,17'd44997,17'd43814,17'd44998,17'd44999,17'd45000,17'd44198,17'd40173,17'd45001,17'd45002,17'd45003,17'd40786,17'd45004,17'd45005,17'd44896,17'd41075,17'd45006,17'd45007,17'd45008,17'd45009,17'd45010,17'd45011,17'd45012,17'd42720,17'd40169,17'd45013,17'd45014,17'd45015,17'd45016,17'd45017,17'd45018,17'd41083,17'd45019,17'd45020,17'd45021,17'd44914,17'd45022,17'd45023,17'd45024,17'd45025,17'd45026,17'd33617,17'd45027,17'd45028,17'd36385,17'd43412,17'd36384,17'd36385,17'd35972,17'd36385,17'd39567,17'd39568,17'd39416,17'd45029,17'd44924,17'd45030,17'd45031,17'd45032,17'd44817,17'd43684,17'd45033,17'd45034,17'd45035,17'd44354,17'd44821,17'd44587,17'd44936,17'd44102,17'd44476,17'd44933,17'd43426,17'd43552,17'd44106,17'd45036,17'd43977,17'd29101,17'd28850,17'd25178,17'd24898,17'd25032,17'd24743,17'd24902,17'd23733,17'd39133,17'd33311,17'd35711,17'd45037,17'd22501,17'd32191,17'd23386,17'd23731,17'd28851,17'd25029,17'd31366,17'd26530,17'd28725,17'd27146,17'd40826,17'd44103,17'd43434,17'd36403,17'd32354,17'd28258,17'd32831,17'd28373,17'd32355,17'd33654,17'd33319,17'd29977,17'd28980,17'd26781,17'd28978,17'd28253,17'd28369,17'd25709,17'd25032,17'd29686,17'd22859,17'd22158,17'd23222,17'd33648,17'd31833,17'd43986,17'd35877,17'd23565,17'd24416,17'd27882,17'd25708,17'd27259,17'd33963,17'd28979,17'd28980,17'd28726,17'd33963,17'd27371,17'd27640,17'd26530,17'd43290,17'd38537,17'd33952,17'd29977,17'd35426,17'd42741,17'd45038,17'd45039,17'd44937,17'd44938,17'd33475,17'd35570,17'd27642,17'd30586,17'd26174,17'd25835,17'd37122,17'd45040,17'd43999,17'd45041,17'd45042,17'd45043,17'd42017,17'd45044,17'd45045,17'd40065,17'd44944,17'd44233,17'd29099,17'd24902,17'd24417,17'd25178,17'd29103,17'd43714,17'd24740,17'd24745,17'd24416,17'd35036,17'd29829,17'd32013,17'd45046,17'd34776,17'd45047,17'd45048,17'd45049,17'd45050,17'd45051,17'd45052,17'd45053,17'd45054,17'd44954,17'd25870,17'd45055,17'd44726,17'd45056,17'd45057,17'd24945,17'd14970,17'd26585,17'd45058,17'd37555,17'd38056,17'd37693,17'd36170,17'd41141,17'd38316,17'd11710,17'd25084,17'd33692,17'd34155,17'd4017,17'd4185,17'd42463,17'd39313,17'd4017,17'd43183,17'd42462,17'd4831,17'd41455,17'd4998,17'd4526,17'd4684,17'd5000,17'd4362,17'd4185,17'd42630,17'd4829,17'd36165,17'd45059,17'd42774,17'd44957,17'd44958,17'd33200,17'd44012,17'd33201,17'd45060,17'd45061,17'd44960,17'd45062,17'd39621,17'd44511,17'd45063,17'd45064,17'd45065,17'd3194,17'd45066,17'd44964,17'd43056,17'd44965,17'd2535,17'd43740,17'd3561,17'd45067,17'd18629,17'd11188,17'd38859,17'd41481,17'd44966,17'd44966,17'd43330,17'd44387,17'd16623,17'd6094,17'd8507,17'd7537,17'd7364,17'd6418,17'd6258,17'd7365,17'd4713,17'd4882,17'd4713,17'd3744,17'd4880,17'd5372,17'd14178,17'd2098,17'd779,17'd1529,17'd44020,17'd417,17'd946,17'd197
},
'{
17'd3903,17'd3902,17'd4426,17'd5646,17'd45068,17'd44388,17'd4244,17'd4088,17'd2422,17'd4247,17'd1416,17'd3905,17'd20404,17'd20404,17'd3905,17'd3905,17'd980,17'd980,17'd652,17'd289,17'd3595,17'd3256,17'd16866,17'd3253,17'd2263,17'd1973,17'd1839,17'd1559,17'd19499,17'd991,17'd826,17'd828,17'd1426,17'd24509,17'd44852,17'd37577,17'd3929,17'd41910,17'd44743,17'd44853,17'd44854,17'd44744,17'd44855,17'd45069,17'd14622,17'd12218,17'd11913,17'd11913,17'd16765,17'd28925,17'd45070,17'd20294,17'd35778,17'd20295,17'd36612,17'd40568,17'd45071,17'd45072,17'd45073,17'd44625,17'd37455,17'd45074,17'd45075,17'd45075,17'd40721,17'd38735,17'd37714,17'd36190,17'd45076,17'd45077,17'd45078,17'd7749,17'd7579,17'd7415,17'd7417,17'd11479,17'd5254,17'd5088,17'd5250,17'd6933,17'd7754,17'd6314,17'd44863,17'd6154,17'd44282,17'd44756,17'd43606,17'd44864,17'd45079,17'd43472,17'd45080,17'd45081,17'd44865,17'd45082,17'd45083,17'd45084,17'd45085,17'd44976,17'd45086,17'd45087,17'd45088,17'd44978,17'd45089,17'd45090,17'd44645,17'd45091,17'd37334,17'd9046,17'd9041,17'd9743,17'd9620,17'd9345,17'd9189,17'd10175,17'd17480,17'd8874,17'd9191,17'd20175,17'd21820,17'd10326,17'd11274,17'd24995,17'd24537,17'd28816,17'd28104,17'd26629,17'd24991,17'd18200,17'd24856,17'd23515,17'd23170,17'd21361,17'd23169,17'd18327,17'd14264,17'd14379,17'd18443,17'd22992,17'd22992,17'd14258,17'd25143,17'd14259,17'd24540,17'd12583,17'd12423,17'd10331,17'd11671,17'd12116,17'd10742,17'd10742,17'd17011,17'd10743,17'd10992,17'd9741,17'd9883,17'd10479,17'd11527,17'd11527,17'd11133,17'd10165,17'd27864,17'd42810,17'd34709,17'd33103,17'd33102,17'd45092,17'd39073,17'd32604,17'd45093,17'd21506,17'd13519,17'd12114,17'd29341,17'd28697,17'd44648,17'd45094,17'd45095,17'd42078,17'd44651,17'd41353,17'd45096,17'd45097,17'd45098,17'd45099,17'd44878,17'd44418,17'd45100,17'd44986,17'd45101,17'd45102,17'd45103,17'd45104,17'd45105,17'd44087,17'd45106,17'd45107,17'd45108,17'd45109,17'd45110,17'd45111,17'd45112,17'd45113,17'd45114,17'd45115,17'd45116,17'd45117,17'd45118,17'd45119,17'd45120,17'd45121,17'd45122,17'd45123,17'd40929,17'd45124,17'd45125,17'd45126,17'd45127,17'd40644,17'd44669,17'd45128,17'd40646,17'd45129,17'd45130,17'd45131,17'd45132,17'd45133,17'd45134,17'd45135,17'd44805,17'd45136,17'd40336,17'd42725,17'd45137,17'd45138,17'd39856,17'd45139,17'd39387,17'd45140,17'd45141,17'd45142,17'd45143,17'd45144,17'd41988,17'd40350,17'd36244,17'd44922,17'd38391,17'd35972,17'd40350,17'd36244,17'd39415,17'd39416,17'd38006,17'd45145,17'd45146,17'd45147,17'd45148,17'd45149,17'd44583,17'd42430,17'd45150,17'd45151,17'd45035,17'd44354,17'd44931,17'd44472,17'd45152,17'd39583,17'd43974,17'd44933,17'd43426,17'd44103,17'd43156,17'd44359,17'd29825,17'd31034,17'd29103,17'd25180,17'd24744,17'd30126,17'd24415,17'd28849,17'd23734,17'd39280,17'd22333,17'd31657,17'd22857,17'd22329,17'd29828,17'd23386,17'd23731,17'd28851,17'd25029,17'd33000,17'd27514,17'd26902,17'd30586,17'd32495,17'd43701,17'd43297,17'd35707,17'd32354,17'd28258,17'd32832,17'd28373,17'd28373,17'd32354,17'd33001,17'd33952,17'd38537,17'd33963,17'd28724,17'd33643,17'd28850,17'd27511,17'd24745,17'd36987,17'd31656,17'd22158,17'd22156,17'd31832,17'd45153,17'd45154,17'd36700,17'd23565,17'd24416,17'd27882,17'd26174,17'd27259,17'd33963,17'd28727,17'd29245,17'd26901,17'd26902,17'd28725,17'd27883,17'd26530,17'd27259,17'd28979,17'd29977,17'd29379,17'd36542,17'd45155,17'd45156,17'd44932,17'd45157,17'd44938,17'd43696,17'd35570,17'd27642,17'd25560,17'd27766,17'd34127,17'd37253,17'd43986,17'd34905,17'd45158,17'd45159,17'd40686,17'd45160,17'd45161,17'd44941,17'd44708,17'd45162,17'd45154,17'd23566,17'd45163,17'd24418,17'd25180,17'd25320,17'd24081,17'd23914,17'd24744,17'd23916,17'd45164,17'd45165,17'd31497,17'd45166,17'd34640,17'd45167,17'd45048,17'd45168,17'd45169,17'd45051,17'd45170,17'd45171,17'd45172,17'd45173,17'd23960,17'd45055,17'd44501,17'd45174,17'd45057,17'd24945,17'd14971,17'd26585,17'd20847,17'd37693,17'd38056,17'd37693,17'd36170,17'd41141,17'd38316,17'd11710,17'd25084,17'd27570,17'd4836,17'd4017,17'd4016,17'd45175,17'd40395,17'd4356,17'd4358,17'd42462,17'd4831,17'd39313,17'd34157,17'd4526,17'd4684,17'd5000,17'd4362,17'd4671,17'd4670,17'd4829,17'd35889,17'd45176,17'd42774,17'd44957,17'd44958,17'd33200,17'd44731,17'd4350,17'd45177,17'd40991,17'd45178,17'd45179,17'd45180,17'd45181,17'd45063,17'd45182,17'd44963,17'd3194,17'd45066,17'd45183,17'd45184,17'd44514,17'd42194,17'd43740,17'd3561,17'd7849,17'd45185,17'd45186,17'd11867,17'd39033,17'd44966,17'd44966,17'd43330,17'd44387,17'd16623,17'd6094,17'd8507,17'd7537,17'd7364,17'd6418,17'd6258,17'd6095,17'd4713,17'd4882,17'd4713,17'd3744,17'd35907,17'd8185,17'd2393,17'd1383,17'd778,17'd1529,17'd44020,17'd418,17'd946,17'd198
},
'{
17'd4244,17'd3902,17'd4426,17'd5646,17'd45068,17'd4889,17'd4427,17'd4088,17'd2422,17'd4247,17'd1416,17'd3905,17'd20404,17'd20404,17'd3905,17'd3905,17'd980,17'd652,17'd29,17'd809,17'd3255,17'd2940,17'd3253,17'd2262,17'd2122,17'd1972,17'd1557,17'd1281,17'd1137,17'd824,17'd667,17'd828,17'd1426,17'd24509,17'd44852,17'd37577,17'd45187,17'd41910,17'd44743,17'd18287,17'd45188,17'd44744,17'd45189,17'd45190,17'd12362,17'd12218,17'd11913,17'd11913,17'd16765,17'd20886,17'd43062,17'd45191,17'd21346,17'd40864,17'd20431,17'd14899,17'd39492,17'd39955,17'd42342,17'd38595,17'd37714,17'd38734,17'd40417,17'd39493,17'd44858,17'd45192,17'd45193,17'd32105,17'd45194,17'd45077,17'd45078,17'd8684,17'd7414,17'd7087,17'd6468,17'd5254,17'd6627,17'd5088,17'd5250,17'd7253,17'd42796,17'd42350,17'd43602,17'd6154,17'd44282,17'd45195,17'd43471,17'd45196,17'd45079,17'd45197,17'd45198,17'd45199,17'd42219,17'd40432,17'd45200,17'd38358,17'd45085,17'd45201,17'd45086,17'd45087,17'd45088,17'd45202,17'd45203,17'd45204,17'd45205,17'd45206,17'd10993,17'd9046,17'd9041,17'd9189,17'd9344,17'd15807,17'd10336,17'd10336,17'd17480,17'd10336,17'd9743,17'd23679,17'd11136,17'd12863,17'd11523,17'd29488,17'd26371,17'd29778,17'd28104,17'd26629,17'd24991,17'd18200,17'd24856,17'd23512,17'd23170,17'd22992,17'd23513,17'd18327,17'd14264,17'd28112,17'd22472,17'd21363,17'd21505,17'd20608,17'd33084,17'd24706,17'd29783,17'd45207,17'd45208,17'd29335,17'd17847,17'd9884,17'd9885,17'd10742,17'd17011,17'd10743,17'd10992,17'd9741,17'd9883,17'd10479,17'd11527,17'd11527,17'd11133,17'd10165,17'd27864,17'd10988,17'd17837,17'd33250,17'd37071,17'd32607,17'd31449,17'd32604,17'd45209,17'd21506,17'd13519,17'd12114,17'd29341,17'd29332,17'd44648,17'd45094,17'd45095,17'd42078,17'd44651,17'd41352,17'd42681,17'd42681,17'd45210,17'd45211,17'd45212,17'd42081,17'd45100,17'd45213,17'd33751,17'd45214,17'd45215,17'd45216,17'd45217,17'd45218,17'd45219,17'd42280,17'd45220,17'd45221,17'd42726,17'd45222,17'd45223,17'd45224,17'd45225,17'd42724,17'd44553,17'd45226,17'd45227,17'd45228,17'd45118,17'd45229,17'd45230,17'd45231,17'd45232,17'd41974,17'd45233,17'd45234,17'd45235,17'd45236,17'd45237,17'd45238,17'd45239,17'd45240,17'd45241,17'd45242,17'd45243,17'd45244,17'd45245,17'd45246,17'd45247,17'd45248,17'd45249,17'd45250,17'd39858,17'd45251,17'd45252,17'd45253,17'd39405,17'd45254,17'd39258,17'd45255,17'd45256,17'd45257,17'd41988,17'd36813,17'd36670,17'd39567,17'd36385,17'd36385,17'd36512,17'd39116,17'd37634,17'd39416,17'd45258,17'd45145,17'd45259,17'd45147,17'd39891,17'd45260,17'd41259,17'd43142,17'd45261,17'd45262,17'd45035,17'd45263,17'd44473,17'd44587,17'd45264,17'd44362,17'd44698,17'd44938,17'd43426,17'd44227,17'd43018,17'd43694,17'd39443,17'd29103,17'd29244,17'd25180,17'd24742,17'd35159,17'd24090,17'd23564,17'd40960,17'd39588,17'd22158,17'd31829,17'd32344,17'd32827,17'd37117,17'd28976,17'd23731,17'd24744,17'd27764,17'd28598,17'd27640,17'd27027,17'd30586,17'd33308,17'd41997,17'd44235,17'd35570,17'd33654,17'd28373,17'd32832,17'd28373,17'd28373,17'd32354,17'd40681,17'd37513,17'd44703,17'd35023,17'd28724,17'd25435,17'd27511,17'd28850,17'd24744,17'd32352,17'd31656,17'd22158,17'd22156,17'd45265,17'd31347,17'd45154,17'd42449,17'd30275,17'd24416,17'd28369,17'd26174,17'd27259,17'd26781,17'd28727,17'd29246,17'd28726,17'd26781,17'd26782,17'd27883,17'd26530,17'd28725,17'd28979,17'd29977,17'd29379,17'd36690,17'd45266,17'd45267,17'd44931,17'd45157,17'd44938,17'd43696,17'd36127,17'd27642,17'd26400,17'd27766,17'd32688,17'd45268,17'd43843,17'd45269,17'd37268,17'd45270,17'd45271,17'd39145,17'd44248,17'd45043,17'd44708,17'd45162,17'd43843,17'd23387,17'd34126,17'd24590,17'd24898,17'd25178,17'd24894,17'd24744,17'd24251,17'd24415,17'd24084,17'd45272,17'd34455,17'd45166,17'd45273,17'd38421,17'd45048,17'd45274,17'd45169,17'd45275,17'd45276,17'd45277,17'd45278,17'd45279,17'd23960,17'd45055,17'd45280,17'd45281,17'd45282,17'd36443,17'd45283,17'd15607,17'd22942,17'd37802,17'd38314,17'd37693,17'd39467,17'd41141,17'd38316,17'd11710,17'd6392,17'd4845,17'd4524,17'd4017,17'd4016,17'd41755,17'd42464,17'd4356,17'd4358,17'd33839,17'd4356,17'd39313,17'd34157,17'd4526,17'd4684,17'd5000,17'd4362,17'd4671,17'd4670,17'd35332,17'd45284,17'd45176,17'd45285,17'd44957,17'd44958,17'd43869,17'd45286,17'd42634,17'd33529,17'd44135,17'd45287,17'd45288,17'd45289,17'd45181,17'd40711,17'd45064,17'd45065,17'd3194,17'd45066,17'd45183,17'd42781,17'd2532,17'd42194,17'd45290,17'd3561,17'd45067,17'd10247,17'd11587,17'd45291,17'd39033,17'd44966,17'd39182,17'd43330,17'd44387,17'd16623,17'd6094,17'd8507,17'd7537,17'd6418,17'd6418,17'd6258,17'd6095,17'd4882,17'd4882,17'd4713,17'd3744,17'd35907,17'd5630,17'd2393,17'd1383,17'd778,17'd1529,17'd44020,17'd418,17'd946,17'd198
},
'{
17'd4244,17'd4891,17'd4426,17'd4734,17'd45068,17'd44388,17'd4244,17'd4088,17'd2422,17'd4247,17'd1416,17'd3905,17'd20404,17'd20404,17'd3905,17'd3905,17'd980,17'd980,17'd652,17'd289,17'd3433,17'd3256,17'd16866,17'd3253,17'd2263,17'd1973,17'd1839,17'd1282,17'd1135,17'd991,17'd992,17'd828,17'd1425,17'd3263,17'd2953,17'd35064,17'd45187,17'd41910,17'd44743,17'd18287,17'd45188,17'd45292,17'd45293,17'd45069,17'd14470,17'd12218,17'd11913,17'd11913,17'd16658,17'd12532,17'd19621,17'd34360,17'd19622,17'd20024,17'd18780,17'd39333,17'd39954,17'd40866,17'd44626,17'd44626,17'd45294,17'd38878,17'd39955,17'd39955,17'd41487,17'd38595,17'd36760,17'd45295,17'd45296,17'd13974,17'd13604,17'd8684,17'd8218,17'd30658,17'd44629,17'd11479,17'd5254,17'd6627,17'd5250,17'd4923,17'd7914,17'd42060,17'd44863,17'd6154,17'd44282,17'd44756,17'd43890,17'd45196,17'd43353,17'd45197,17'd45198,17'd45199,17'd42219,17'd45297,17'd45200,17'd45298,17'd45299,17'd45300,17'd45301,17'd45302,17'd33870,17'd45202,17'd45303,17'd45304,17'd45305,17'd45306,17'd45307,17'd23517,17'd9040,17'd9189,17'd9346,17'd9345,17'd9189,17'd10336,17'd17480,17'd8874,17'd9191,17'd9338,17'd9472,17'd11133,17'd14673,17'd15055,17'd25925,17'd26370,17'd28104,17'd26629,17'd24991,17'd18200,17'd25927,17'd23512,17'd23170,17'd22992,17'd23513,17'd23169,17'd23167,17'd28112,17'd21361,17'd21505,17'd21505,17'd21363,17'd26258,17'd24706,17'd29783,17'd14382,17'd12423,17'd12585,17'd11276,17'd9884,17'd9885,17'd9885,17'd17011,17'd10742,17'd11136,17'd9885,17'd9883,17'd10479,17'd12863,17'd11527,17'd11133,17'd10326,17'd27864,17'd42810,17'd34709,17'd33103,17'd32773,17'd32938,17'd33579,17'd32604,17'd45209,17'd30684,17'd12259,17'd12114,17'd43363,17'd17009,17'd45308,17'd45309,17'd45310,17'd45311,17'd45098,17'd41799,17'd45312,17'd42681,17'd45210,17'd41664,17'd41519,17'd45313,17'd45096,17'd45314,17'd45315,17'd45316,17'd45317,17'd45318,17'd45319,17'd45320,17'd45321,17'd45322,17'd40339,17'd40339,17'd45323,17'd45107,17'd45107,17'd41983,17'd40796,17'd44682,17'd45324,17'd45325,17'd45326,17'd45327,17'd45328,17'd45329,17'd45330,17'd45331,17'd44313,17'd45332,17'd45333,17'd45334,17'd45335,17'd45336,17'd45337,17'd45338,17'd45339,17'd45340,17'd45341,17'd45342,17'd45343,17'd45344,17'd45345,17'd45346,17'd45347,17'd45348,17'd45349,17'd45350,17'd39249,17'd45351,17'd45352,17'd45353,17'd45354,17'd45355,17'd45356,17'd45357,17'd45358,17'd45359,17'd45360,17'd45361,17'd38391,17'd38958,17'd36244,17'd38391,17'd36512,17'd39116,17'd37634,17'd36669,17'd38006,17'd45362,17'd45259,17'd45363,17'd45364,17'd45365,17'd45366,17'd45367,17'd45368,17'd45369,17'd45035,17'd45263,17'd44473,17'd45370,17'd45038,17'd43974,17'd44933,17'd44938,17'd44227,17'd43426,17'd43018,17'd38156,17'd31034,17'd30432,17'd29976,17'd25032,17'd34467,17'd30431,17'd23731,17'd30275,17'd34894,17'd22327,17'd32345,17'd36984,17'd22506,17'd22679,17'd37117,17'd23565,17'd24249,17'd24417,17'd27512,17'd28720,17'd28725,17'd26901,17'd34637,17'd38975,17'd41997,17'd42436,17'd31354,17'd33654,17'd28373,17'd28258,17'd28134,17'd28373,17'd33319,17'd40681,17'd44826,17'd34767,17'd27371,17'd28252,17'd25435,17'd25438,17'd27511,17'd24252,17'd38976,17'd34458,17'd22158,17'd23040,17'd43158,17'd32009,17'd43986,17'd38669,17'd23732,17'd24742,17'd28369,17'd25833,17'd27259,17'd26781,17'd29245,17'd29245,17'd28486,17'd27027,17'd28725,17'd27883,17'd26530,17'd28853,17'd28727,17'd29977,17'd27642,17'd33790,17'd45371,17'd45372,17'd44931,17'd43546,17'd44938,17'd43696,17'd36127,17'd31352,17'd25699,17'd28602,17'd25710,17'd38542,17'd24094,17'd23220,17'd45373,17'd45374,17'd45375,17'd45376,17'd45167,17'd45377,17'd40834,17'd45378,17'd45379,17'd30128,17'd45380,17'd44116,17'd24745,17'd25180,17'd26900,17'd23915,17'd24742,17'd24090,17'd23209,17'd45381,17'd31659,17'd45382,17'd45383,17'd39452,17'd45384,17'd45385,17'd45169,17'd45386,17'd45387,17'd45388,17'd45389,17'd38832,17'd45390,17'd23441,17'd45280,17'd45391,17'd36441,17'd37027,17'd45283,17'd15725,17'd37940,17'd38056,17'd45392,17'd37693,17'd39467,17'd37557,17'd38316,17'd11710,17'd6392,17'd4687,17'd4524,17'd45393,17'd41890,17'd45175,17'd42631,17'd4017,17'd4358,17'd4357,17'd45393,17'd39313,17'd34157,17'd5000,17'd5156,17'd4525,17'd43183,17'd4671,17'd4670,17'd35332,17'd45394,17'd45395,17'd45285,17'd44957,17'd45396,17'd43869,17'd44731,17'd4350,17'd33689,17'd43870,17'd45397,17'd45398,17'd45180,17'd45399,17'd45400,17'd45401,17'd45065,17'd3194,17'd45066,17'd45183,17'd42781,17'd2532,17'd42194,17'd45290,17'd3702,17'd45402,17'd18755,17'd45403,17'd11720,17'd39033,17'd39182,17'd39182,17'd43330,17'd37959,17'd6094,17'd6416,17'd4714,17'd8187,17'd6418,17'd6418,17'd6258,17'd6095,17'd4882,17'd5958,17'd4713,17'd3744,17'd35907,17'd5630,17'd14178,17'd779,17'd778,17'd1529,17'd44020,17'd418,17'd946,17'd44020
},
'{
17'd4244,17'd4891,17'd5201,17'd4734,17'd45068,17'd4889,17'd4244,17'd4245,17'd2422,17'd4247,17'd1416,17'd3905,17'd3905,17'd3905,17'd3905,17'd3905,17'd980,17'd652,17'd29,17'd809,17'd3254,17'd2940,17'd3253,17'd2262,17'd2263,17'd1973,17'd1839,17'd1282,17'd1135,17'd19244,17'd827,17'd827,17'd45404,17'd1427,17'd2953,17'd28197,17'd45187,17'd41910,17'd44743,17'd45405,17'd45188,17'd25394,17'd45189,17'd45406,17'd20885,17'd12362,17'd11913,17'd11764,17'd22630,17'd19006,17'd10816,17'd8214,17'd19513,17'd19388,17'd38211,17'd39044,17'd43065,17'd45407,17'd15390,17'd15390,17'd37178,17'd38594,17'd40108,17'd39955,17'd41487,17'd45408,17'd35355,17'd32264,17'd45296,17'd45409,17'd45410,17'd8684,17'd8218,17'd8368,17'd6468,17'd9302,17'd7088,17'd6627,17'd4924,17'd7253,17'd6475,17'd42060,17'd6312,17'd42663,17'd44282,17'd44756,17'd44757,17'd6329,17'd43353,17'd45197,17'd43075,17'd45411,17'd45412,17'd45413,17'd39506,17'd45298,17'd45414,17'd45415,17'd45416,17'd45417,17'd45418,17'd45419,17'd45420,17'd44032,17'd45421,17'd45422,17'd45423,17'd23517,17'd11402,17'd9043,17'd10335,17'd10173,17'd9189,17'd10175,17'd17480,17'd8874,17'd9190,17'd23679,17'd11136,17'd12863,17'd11522,17'd15055,17'd25925,17'd26370,17'd28104,17'd26629,17'd24991,17'd24856,17'd25927,17'd23856,17'd24209,17'd21505,17'd14258,17'd23169,17'd23167,17'd24995,17'd21363,17'd23170,17'd24209,17'd23170,17'd26150,17'd26258,17'd33572,17'd14382,17'd28821,17'd34826,17'd10331,17'd9884,17'd9885,17'd9885,17'd17011,17'd10742,17'd11136,17'd9885,17'd9883,17'd11134,17'd12863,17'd11527,17'd11133,17'd10326,17'd27739,17'd10852,17'd40746,17'd38912,17'd32773,17'd37071,17'd33416,17'd33247,17'd45209,17'd13518,17'd12259,17'd11957,17'd10735,17'd17009,17'd45308,17'd45309,17'd45310,17'd45311,17'd45099,17'd45424,17'd45312,17'd45312,17'd41354,17'd44878,17'd45424,17'd45313,17'd45425,17'd45426,17'd45427,17'd45428,17'd45429,17'd45430,17'd45431,17'd45432,17'd43820,17'd45433,17'd45434,17'd45435,17'd45436,17'd45106,17'd45437,17'd45438,17'd45439,17'd45440,17'd45441,17'd45442,17'd45443,17'd45444,17'd44570,17'd45445,17'd45446,17'd45447,17'd45448,17'd44998,17'd45449,17'd45450,17'd45451,17'd45452,17'd45453,17'd45454,17'd45455,17'd45456,17'd45457,17'd45458,17'd45459,17'd45460,17'd45461,17'd42417,17'd45462,17'd45463,17'd45464,17'd45465,17'd45466,17'd45467,17'd45468,17'd45469,17'd45470,17'd42284,17'd45471,17'd35678,17'd45472,17'd45473,17'd36513,17'd45474,17'd36670,17'd39415,17'd44922,17'd36385,17'd39116,17'd39116,17'd37634,17'd36669,17'd38006,17'd45475,17'd45259,17'd45363,17'd45476,17'd45365,17'd44220,17'd45477,17'd45478,17'd45479,17'd43972,17'd45263,17'd44473,17'd45480,17'd45481,17'd44698,17'd44938,17'd44227,17'd45482,17'd45483,17'd44699,17'd29825,17'd32353,17'd29533,17'd25032,17'd24895,17'd24252,17'd24415,17'd23917,17'd23918,17'd31655,17'd22504,17'd41867,17'd36984,17'd22333,17'd39131,17'd37386,17'd23920,17'd32659,17'd24896,17'd28717,17'd25708,17'd27027,17'd31035,17'd35011,17'd40958,17'd41863,17'd45484,17'd31503,17'd32017,17'd28258,17'd32831,17'd32354,17'd28134,17'd33319,17'd37513,17'd28980,17'd34767,17'd26782,17'd31351,17'd25435,17'd25438,17'd29244,17'd24743,17'd38976,17'd23038,17'd22158,17'd22163,17'd45485,17'd39745,17'd43986,17'd38668,17'd31033,17'd24417,17'd27765,17'd25707,17'd27259,17'd26781,17'd29246,17'd29246,17'd28979,17'd27027,17'd28725,17'd27514,17'd26062,17'd28978,17'd31035,17'd27642,17'd39437,17'd39741,17'd45486,17'd45487,17'd44931,17'd45157,17'd44227,17'd33308,17'd36127,17'd31352,17'd26400,17'd28602,17'd31521,17'd45488,17'd45379,17'd32009,17'd38173,17'd45489,17'd23744,17'd45490,17'd38421,17'd34484,17'd40834,17'd45491,17'd45492,17'd23215,17'd29827,17'd24087,17'd24416,17'd24082,17'd26900,17'd24742,17'd37388,17'd45493,17'd23208,17'd23390,17'd43982,17'd45494,17'd45495,17'd45496,17'd45497,17'd45498,17'd45169,17'd45499,17'd45500,17'd45501,17'd45502,17'd45503,17'd45504,17'd22387,17'd45505,17'd45506,17'd45507,17'd37027,17'd23116,17'd15725,17'd43581,17'd38314,17'd45392,17'd45508,17'd39467,17'd37557,17'd38316,17'd11710,17'd6392,17'd4687,17'd4524,17'd4017,17'd45393,17'd42463,17'd39165,17'd4017,17'd4358,17'd4515,17'd4017,17'd39165,17'd34157,17'd5156,17'd5156,17'd4525,17'd4833,17'd4016,17'd42630,17'd35332,17'd35602,17'd45509,17'd42774,17'd45510,17'd43731,17'd6537,17'd44731,17'd4350,17'd45511,17'd42324,17'd45397,17'd40709,17'd45180,17'd45512,17'd45400,17'd45513,17'd45065,17'd3194,17'd45066,17'd44964,17'd42781,17'd44849,17'd2536,17'd45514,17'd3702,17'd9789,17'd10523,17'd45515,17'd11720,17'd39033,17'd39182,17'd38860,17'd38861,17'd37959,17'd6094,17'd6416,17'd6416,17'd6416,17'd8507,17'd6418,17'd6258,17'd6095,17'd4882,17'd5958,17'd4713,17'd3744,17'd35907,17'd5630,17'd14178,17'd779,17'd13573,17'd941,17'd44020,17'd418,17'd599,17'd43878
},
'{
17'd4428,17'd4891,17'd5202,17'd6263,17'd6263,17'd4888,17'd3903,17'd15746,17'd10535,17'd2595,17'd17,17'd1416,17'd468,17'd2938,17'd653,17'd652,17'd980,17'd980,17'd652,17'd981,17'd31,17'd2259,17'd45516,17'd2262,17'd2263,17'd1973,17'd1839,17'd1282,17'd1135,17'd824,17'd666,17'd480,17'd45404,17'd3266,17'd45517,17'd3447,17'd13443,17'd44619,17'd45518,17'd29619,17'd24516,17'd25394,17'd45519,17'd30057,17'd45520,17'd12362,17'd12361,17'd13969,17'd12681,17'd19006,17'd11087,17'd22464,17'd19512,17'd19513,17'd36611,17'd45521,17'd45522,17'd45523,17'd45524,17'd45525,17'd16414,17'd42045,17'd42202,17'd44747,17'd38595,17'd37455,17'd32419,17'd33862,17'd31577,17'd45526,17'd45527,17'd7413,17'd8536,17'd12220,17'd8370,17'd11479,17'd5254,17'd6627,17'd4924,17'd4463,17'd6630,17'd6314,17'd42350,17'd45528,17'd45529,17'd45530,17'd43889,17'd43204,17'd45196,17'd45531,17'd42354,17'd40430,17'd45532,17'd45533,17'd45534,17'd45535,17'd45536,17'd45537,17'd45538,17'd45539,17'd45540,17'd45541,17'd45542,17'd45543,17'd45544,17'd45545,17'd45546,17'd29919,17'd19033,17'd9189,17'd10335,17'd10173,17'd9189,17'd8874,17'd10174,17'd8874,17'd9190,17'd23679,17'd10169,17'd13647,17'd17478,17'd24362,17'd25925,17'd26872,17'd28343,17'd29778,17'd27347,17'd25672,17'd26370,17'd23856,17'd22818,17'd20314,17'd18197,17'd18806,17'd18557,17'd24995,17'd25926,17'd24705,17'd24705,17'd26494,17'd26151,17'd26258,17'd24706,17'd24540,17'd27350,17'd11525,17'd19280,17'd10330,17'd10169,17'd9885,17'd17011,17'd10742,17'd10742,17'd9885,17'd17719,17'd10479,17'd11133,17'd11133,17'd19532,17'd10326,17'd27236,17'd24703,17'd23164,17'd33419,17'd32609,17'd33102,17'd33416,17'd33247,17'd45547,17'd45548,17'd12260,17'd17598,17'd10604,17'd45549,17'd28698,17'd45550,17'd45310,17'd45551,17'd44414,17'd45424,17'd42953,17'd45552,17'd42953,17'd45553,17'd44878,17'd41352,17'd45554,17'd45555,17'd45556,17'd45428,17'd45557,17'd45558,17'd45320,17'd45559,17'd45560,17'd39714,17'd40026,17'd45561,17'd45562,17'd44213,17'd43675,17'd45563,17'd45564,17'd44662,17'd45565,17'd45566,17'd45567,17'd45568,17'd45569,17'd45570,17'd45571,17'd45456,17'd45572,17'd45573,17'd45574,17'd45226,17'd45575,17'd45576,17'd45577,17'd45578,17'd45579,17'd45580,17'd45581,17'd45582,17'd45583,17'd45584,17'd45585,17'd45586,17'd45587,17'd45588,17'd45589,17'd45590,17'd45591,17'd45592,17'd45593,17'd45594,17'd45595,17'd45596,17'd35973,17'd45597,17'd38645,17'd38391,17'd37227,17'd36812,17'd36669,17'd39415,17'd39567,17'd36384,17'd45598,17'd45599,17'd37228,17'd37367,17'd45600,17'd45601,17'd45602,17'd45603,17'd41258,17'd45604,17'd45605,17'd45606,17'd45607,17'd45608,17'd44100,17'd44354,17'd44472,17'd45609,17'd39583,17'd43974,17'd43434,17'd44235,17'd45610,17'd45610,17'd43979,17'd25317,17'd25179,17'd32668,17'd32007,17'd24897,17'd28718,17'd24743,17'd23731,17'd23734,17'd39280,17'd23573,17'd41729,17'd23222,17'd22334,17'd39131,17'd29829,17'd23920,17'd28975,17'd28254,17'd27638,17'd26530,17'd32016,17'd26901,17'd33942,17'd45611,17'd45612,17'd40520,17'd32356,17'd40051,17'd45613,17'd40367,17'd27884,17'd28370,17'd25697,17'd25828,17'd28727,17'd26781,17'd26902,17'd26903,17'd27638,17'd25709,17'd30432,17'd23731,17'd45614,17'd40523,17'd32346,17'd38041,17'd45615,17'd22334,17'd45616,17'd35865,17'd24086,17'd28851,17'd25317,17'd26174,17'd27371,17'd28726,17'd40371,17'd45617,17'd28726,17'd27146,17'd33478,17'd33642,17'd25565,17'd27260,17'd36542,17'd36264,17'd35152,17'd44827,17'd45618,17'd45619,17'd45620,17'd45621,17'd43552,17'd42890,17'd38025,17'd28727,17'd26902,17'd26064,17'd29548,17'd41123,17'd44702,17'd33649,17'd38173,17'd45622,17'd45623,17'd45624,17'd45625,17'd45626,17'd45627,17'd45628,17'd39441,17'd22679,17'd32191,17'd23920,17'd43852,17'd23915,17'd24900,17'd30431,17'd45629,17'd42161,17'd31341,17'd22680,17'd22166,17'd22686,17'd45630,17'd45631,17'd45047,17'd45632,17'd45633,17'd31529,17'd45634,17'd45635,17'd45636,17'd45637,17'd45638,17'd22387,17'd45639,17'd45640,17'd45641,17'd29297,17'd15340,17'd18260,17'd24152,17'd39162,17'd45642,17'd45643,17'd39771,17'd36310,17'd36031,17'd12905,17'd6392,17'd4687,17'd4838,17'd33041,17'd4364,17'd45644,17'd39773,17'd4017,17'd4833,17'd4515,17'd4356,17'd33534,17'd38058,17'd4995,17'd4526,17'd4526,17'd4189,17'd33533,17'd42772,17'd4669,17'd6206,17'd45645,17'd45285,17'd4178,17'd44506,17'd44133,17'd45646,17'd45647,17'd42633,17'd45648,17'd45287,17'd45649,17'd45650,17'd39024,17'd3192,17'd45651,17'd45652,17'd44739,17'd45066,17'd45653,17'd45654,17'd42476,17'd3057,17'd45655,17'd41905,17'd45656,17'd10247,17'd45657,17'd11720,17'd11867,17'd39483,17'd38334,17'd38072,17'd13176,17'd16492,17'd6258,17'd6418,17'd8507,17'd35769,17'd7537,17'd35769,17'd8186,17'd5789,17'd5789,17'd4423,17'd4085,17'd8185,17'd2393,17'd15233,17'd15233,17'd1672,17'd940,17'd198,17'd946,17'd195,17'd201
},
'{
17'd4428,17'd4891,17'd5202,17'd6263,17'd6263,17'd4888,17'd4892,17'd15746,17'd17917,17'd2595,17'd17,17'd1416,17'd468,17'd468,17'd653,17'd652,17'd980,17'd652,17'd29,17'd981,17'd31,17'd32,17'd3103,17'd2262,17'd2263,17'd1973,17'd1839,17'd1282,17'd1135,17'd824,17'd666,17'd482,17'd45404,17'd3266,17'd45658,17'd2801,17'd13443,17'd44619,17'd45518,17'd29619,17'd24516,17'd30204,17'd45519,17'd30057,17'd45520,17'd20885,17'd12361,17'd13969,17'd12681,17'd17204,17'd11915,17'd12533,17'd16518,17'd19755,17'd45659,17'd18661,17'd45660,17'd43600,17'd45661,17'd45662,17'd41486,17'd45663,17'd39954,17'd40866,17'd45408,17'd45664,17'd35496,17'd45665,17'd31422,17'd45666,17'd13847,17'd6931,17'd8536,17'd12220,17'd8370,17'd4927,17'd4926,17'd6627,17'd4924,17'd6934,17'd6776,17'd6315,17'd42350,17'd45667,17'd45529,17'd45530,17'd44156,17'd43204,17'd6162,17'd45668,17'd45669,17'd40430,17'd45670,17'd45671,17'd45672,17'd45673,17'd45674,17'd45675,17'd45676,17'd8866,17'd45677,17'd45678,17'd45679,17'd45680,17'd45681,17'd45545,17'd45682,17'd29919,17'd19033,17'd9189,17'd26153,17'd16552,17'd9743,17'd8874,17'd10174,17'd10174,17'd9743,17'd22812,17'd10332,17'd34205,17'd23513,17'd24362,17'd25925,17'd27123,17'd26757,17'd29778,17'd29640,17'd27483,17'd26370,17'd23856,17'd23514,17'd20314,17'd17722,17'd18806,17'd18557,17'd19408,17'd23170,17'd24031,17'd25526,17'd41187,17'd45683,17'd24993,17'd24706,17'd45684,17'd45207,17'd34205,17'd13647,17'd19280,17'd10169,17'd9885,17'd17011,17'd10742,17'd10743,17'd10743,17'd10856,17'd11134,17'd12863,17'd11133,17'd19532,17'd10165,17'd41194,17'd24703,17'd28938,17'd33419,17'd32940,17'd31778,17'd33582,17'd33099,17'd45547,17'd14526,17'd12260,17'd11666,17'd10604,17'd16908,17'd45685,17'd45550,17'd45310,17'd40892,17'd45686,17'd45687,17'd40895,17'd45688,17'd45689,17'd45690,17'd45691,17'd44878,17'd45692,17'd45693,17'd45556,17'd45694,17'd45695,17'd45696,17'd45320,17'd45697,17'd41850,17'd45698,17'd45699,17'd42282,17'd45700,17'd42420,17'd45701,17'd45702,17'd45703,17'd45021,17'd45704,17'd45705,17'd45705,17'd45706,17'd41394,17'd45707,17'd45708,17'd45709,17'd45710,17'd45711,17'd44910,17'd45018,17'd45712,17'd45713,17'd45714,17'd45715,17'd45716,17'd45717,17'd45718,17'd43242,17'd45719,17'd45720,17'd45721,17'd39242,17'd45722,17'd45723,17'd45724,17'd45725,17'd45726,17'd45727,17'd45728,17'd45729,17'd45730,17'd45731,17'd45732,17'd45733,17'd36244,17'd38391,17'd36812,17'd37634,17'd44922,17'd39415,17'd43680,17'd36385,17'd45734,17'd45735,17'd37092,17'd45258,17'd45736,17'd45737,17'd45738,17'd45739,17'd45740,17'd44583,17'd45741,17'd45742,17'd45743,17'd45744,17'd44473,17'd44472,17'd44587,17'd38971,17'd39583,17'd43844,17'd42740,17'd44235,17'd45745,17'd45745,17'd43979,17'd27765,17'd25179,17'd29533,17'd25180,17'd24898,17'd28595,17'd28718,17'd30879,17'd40960,17'd45746,17'd35429,17'd45615,17'd30727,17'd30426,17'd32827,17'd23567,17'd23918,17'd24743,17'd27512,17'd27513,17'd27259,17'd30735,17'd33163,17'd40959,17'd45747,17'd45748,17'd33790,17'd35707,17'd39438,17'd39743,17'd32356,17'd27884,17'd27884,17'd25555,17'd25828,17'd28979,17'd26781,17'd26782,17'd26903,17'd27513,17'd25709,17'd25179,17'd24086,17'd34482,17'd40523,17'd32346,17'd38041,17'd41423,17'd22333,17'd36543,17'd35865,17'd24086,17'd24745,17'd28130,17'd26174,17'd27371,17'd28726,17'd40371,17'd45617,17'd28486,17'd33154,17'd42437,17'd45749,17'd43837,17'd33155,17'd33309,17'd33476,17'd37658,17'd43693,17'd45750,17'd45751,17'd45752,17'd45753,17'd42600,17'd34105,17'd38025,17'd31035,17'd26782,17'd41588,17'd37252,17'd41741,17'd45754,17'd45755,17'd45756,17'd45757,17'd45758,17'd45759,17'd45490,17'd45760,17'd45761,17'd45762,17'd35319,17'd22332,17'd32513,17'd30127,17'd24590,17'd42012,17'd32659,17'd45763,17'd41123,17'd25181,17'd45764,17'd22677,17'd45765,17'd40522,17'd45766,17'd45767,17'd41285,17'd45768,17'd45633,17'd45769,17'd45770,17'd45635,17'd45771,17'd45772,17'd45773,17'd45774,17'd45775,17'd23281,17'd24801,17'd12622,17'd15340,17'd18620,17'd24152,17'd22250,17'd45776,17'd45643,17'd39771,17'd36310,17'd36031,17'd12905,17'd6392,17'd5005,17'd5144,17'd4186,17'd42462,17'd40395,17'd39469,17'd4017,17'd4833,17'd4358,17'd4356,17'd33534,17'd33532,17'd4995,17'd5156,17'd4526,17'd33841,17'd44009,17'd42772,17'd4669,17'd6206,17'd45645,17'd45285,17'd4178,17'd44506,17'd44133,17'd45646,17'd45647,17'd42633,17'd45777,17'd45287,17'd45778,17'd39172,17'd39024,17'd45779,17'd45780,17'd44738,17'd45781,17'd45782,17'd45653,17'd45654,17'd45783,17'd3056,17'd45784,17'd45785,17'd45786,17'd45787,17'd45657,17'd11866,17'd39790,17'd39483,17'd41481,17'd38072,17'd13176,17'd16492,17'd16492,17'd6418,17'd6418,17'd35769,17'd7537,17'd35769,17'd35769,17'd6258,17'd5789,17'd4423,17'd4085,17'd8185,17'd5940,17'd14586,17'd15233,17'd2560,17'd45788,17'd198,17'd946,17'd600,17'd45789
},
'{
17'd4428,17'd4891,17'd5201,17'd6263,17'd6263,17'd4888,17'd4892,17'd15746,17'd17917,17'd2595,17'd17,17'd1416,17'd1416,17'd1416,17'd653,17'd652,17'd980,17'd980,17'd652,17'd809,17'd1129,17'd2259,17'd45516,17'd2262,17'd2785,17'd2785,17'd19608,17'd1282,17'd19499,17'd824,17'd666,17'd667,17'd45404,17'd3437,17'd2798,17'd2801,17'd13443,17'd45790,17'd24680,17'd29619,17'd24516,17'd25394,17'd45519,17'd30057,17'd45520,17'd12361,17'd12530,17'd13969,17'd19006,17'd17689,17'd11915,17'd11087,17'd19893,17'd39797,17'd35212,17'd45791,17'd18302,17'd14630,17'd45792,17'd45793,17'd17211,17'd45794,17'd45795,17'd38469,17'd38345,17'd45796,17'd45797,17'd45798,17'd31270,17'd45799,17'd45800,17'd7250,17'd8536,17'd8687,17'd12219,17'd44630,17'd5254,17'd6627,17'd4924,17'd6933,17'd6630,17'd6314,17'd6480,17'd45667,17'd45529,17'd45530,17'd42504,17'd44028,17'd45196,17'd45668,17'd45669,17'd45801,17'd45802,17'd45671,17'd45803,17'd45673,17'd45674,17'd45675,17'd45804,17'd45805,17'd45806,17'd45807,17'd45808,17'd45809,17'd45681,17'd45810,17'd45811,17'd45812,17'd19285,17'd9192,17'd9743,17'd16552,17'd10335,17'd10335,17'd15944,17'd10174,17'd9743,17'd9340,17'd13522,17'd11525,17'd17478,17'd24362,17'd25925,17'd27123,17'd26757,17'd26370,17'd29640,17'd27483,17'd25927,17'd23512,17'd22818,17'd20314,17'd17722,17'd18806,17'd18557,17'd19408,17'd24992,17'd24538,17'd24857,17'd25526,17'd26628,17'd24993,17'd24363,17'd28112,17'd13367,17'd13368,17'd11525,17'd19280,17'd10024,17'd9885,17'd17011,17'd10743,17'd10743,17'd10743,17'd9885,17'd9883,17'd11670,17'd11670,17'd10165,17'd10165,17'd41194,17'd45813,17'd18683,17'd33419,17'd32940,17'd31451,17'd33736,17'd31139,17'd45814,17'd14809,17'd12260,17'd11520,17'd10604,17'd16908,17'd45815,17'd45816,17'd45817,17'd45818,17'd45819,17'd45820,17'd40895,17'd45821,17'd41665,17'd45822,17'd45823,17'd45691,17'd45692,17'd45824,17'd45825,17'd45826,17'd45827,17'd45828,17'd45431,17'd45829,17'd41714,17'd41850,17'd45830,17'd45831,17'd42421,17'd45434,17'd45832,17'd45437,17'd45833,17'd45834,17'd45835,17'd45836,17'd45836,17'd45837,17'd45838,17'd45567,17'd45839,17'd45840,17'd45841,17'd45842,17'd45843,17'd45844,17'd45845,17'd45846,17'd39548,17'd45847,17'd45848,17'd45837,17'd40937,17'd45109,17'd45849,17'd39241,17'd45850,17'd45851,17'd45852,17'd45853,17'd45854,17'd45855,17'd45856,17'd45857,17'd45858,17'd45859,17'd45860,17'd35834,17'd35972,17'd36670,17'd38391,17'd38391,17'd36812,17'd37228,17'd37366,17'd39568,17'd43274,17'd43412,17'd45861,17'd45862,17'd37096,17'd39412,17'd45863,17'd45864,17'd45865,17'd45866,17'd45867,17'd45868,17'd45869,17'd45478,17'd45870,17'd45871,17'd44473,17'd44472,17'd45370,17'd45872,17'd44362,17'd43844,17'd43433,17'd43560,17'd45873,17'd45745,17'd43979,17'd27765,17'd25178,17'd29976,17'd25030,17'd25029,17'd34283,17'd24252,17'd31033,17'd34894,17'd45874,17'd45875,17'd45615,17'd22861,17'd30427,17'd22503,17'd23736,17'd23564,17'd24744,17'd25177,17'd30606,17'd28853,17'd28727,17'd32016,17'd43021,17'd40217,17'd37657,17'd38025,17'd36541,17'd35425,17'd36403,17'd31354,17'd27761,17'd27761,17'd38537,17'd28726,17'd28486,17'd26782,17'd27259,17'd27515,17'd30734,17'd28717,17'd25031,17'd23732,17'd39278,17'd22677,17'd32666,17'd45876,17'd45877,17'd22856,17'd23569,17'd29099,17'd31033,17'd24895,17'd28600,17'd27515,17'd28725,17'd28726,17'd37513,17'd37513,17'd34637,17'd40826,17'd43548,17'd42885,17'd44934,17'd44478,17'd45878,17'd43696,17'd41108,17'd44822,17'd45879,17'd45870,17'd45880,17'd45881,17'd41582,17'd33790,17'd37908,17'd28486,17'd26782,17'd27513,17'd35735,17'd37922,17'd32190,17'd45882,17'd30620,17'd45883,17'd45884,17'd45885,17'd45886,17'd45887,17'd45496,17'd44718,17'd45888,17'd33645,17'd37533,17'd29099,17'd23382,17'd45889,17'd24901,17'd35999,17'd37407,17'd23738,17'd44110,17'd30427,17'd45890,17'd33314,17'd22339,17'd45891,17'd41285,17'd45892,17'd45893,17'd45894,17'd45895,17'd45896,17'd45897,17'd45898,17'd45899,17'd45900,17'd45901,17'd23281,17'd45902,17'd29297,17'd15476,17'd18620,17'd23463,17'd22250,17'd45776,17'd45903,17'd39771,17'd36310,17'd12761,17'd12622,17'd6221,17'd4687,17'd4838,17'd43584,17'd4363,17'd42631,17'd42464,17'd4357,17'd4359,17'd4358,17'd4017,17'd33534,17'd33532,17'd4995,17'd5156,17'd5156,17'd4999,17'd39468,17'd42772,17'd4669,17'd6206,17'd45645,17'd42774,17'd4178,17'd43588,17'd43869,17'd44133,17'd45904,17'd42633,17'd44135,17'd45905,17'd45906,17'd45907,17'd45908,17'd45909,17'd45780,17'd44963,17'd3047,17'd45910,17'd2881,17'd43327,17'd45911,17'd42333,17'd41770,17'd4552,17'd10071,17'd10523,17'd45657,17'd11587,17'd11048,17'd39948,17'd41481,17'd38072,17'd13176,17'd16492,17'd16492,17'd6418,17'd6418,17'd35769,17'd7537,17'd35769,17'd35769,17'd6258,17'd5789,17'd4423,17'd4085,17'd8185,17'd2393,17'd2394,17'd2394,17'd1950,17'd45788,17'd197,17'd599,17'd600,17'd45912
},
'{
17'd4428,17'd4891,17'd5201,17'd6263,17'd6263,17'd4888,17'd4892,17'd15746,17'd17917,17'd2595,17'd17,17'd17,17'd1416,17'd1416,17'd653,17'd653,17'd980,17'd653,17'd29,17'd809,17'd1129,17'd32,17'd3103,17'd2262,17'd2785,17'd1973,17'd1702,17'd1282,17'd19499,17'd825,17'd666,17'd667,17'd45404,17'd3437,17'd2798,17'd2801,17'd13443,17'd15123,17'd44620,17'd29619,17'd24516,17'd25394,17'd45519,17'd30057,17'd45520,17'd16765,17'd12361,17'd13969,17'd19382,17'd17689,17'd18533,17'd30356,17'd16766,17'd39797,17'd19623,17'd45913,17'd39333,17'd16524,17'd45914,17'd45915,17'd14349,17'd17099,17'd45916,17'd43884,17'd44626,17'd45917,17'd33064,17'd45918,17'd45919,17'd45920,17'd45921,17'd7250,17'd8687,17'd45922,17'd13212,17'd9302,17'd4926,17'd6627,17'd4924,17'd7089,17'd6776,17'd6314,17'd6480,17'd45667,17'd45529,17'd45530,17'd42504,17'd43073,17'd6162,17'd45668,17'd45669,17'd45801,17'd45802,17'd45923,17'd45803,17'd45924,17'd45925,17'd45926,17'd45927,17'd45805,17'd45928,17'd45929,17'd45930,17'd7935,17'd44407,17'd43902,17'd45931,17'd45932,17'd8566,17'd8873,17'd10336,17'd16552,17'd10173,17'd10173,17'd10173,17'd10335,17'd9743,17'd10026,17'd33725,17'd34205,17'd23513,17'd24362,17'd25925,17'd25927,17'd26872,17'd26370,17'd27483,17'd29640,17'd25927,17'd23512,17'd22818,17'd20314,17'd17722,17'd18806,17'd18557,17'd19408,17'd24208,17'd26493,17'd27483,17'd24857,17'd26871,17'd26372,17'd24539,17'd29488,17'd35801,17'd35799,17'd13368,17'd19280,17'd19278,17'd10024,17'd9741,17'd10743,17'd10743,17'd10743,17'd9885,17'd11277,17'd10479,17'd11670,17'd10330,17'd10165,17'd41194,17'd45813,17'd18683,17'd33419,17'd32774,17'd31451,17'd33583,17'd30085,17'd45933,17'd13643,17'd12260,17'd11395,17'd16320,17'd45934,17'd45935,17'd45816,17'd45817,17'd41039,17'd45936,17'd45820,17'd45690,17'd45821,17'd41665,17'd45937,17'd40610,17'd45823,17'd40895,17'd45938,17'd45939,17'd45940,17'd45941,17'd45942,17'd45943,17'd45944,17'd45945,17'd45946,17'd45947,17'd45948,17'd45949,17'd39881,17'd45950,17'd45951,17'd45952,17'd43531,17'd45833,17'd45953,17'd45587,17'd45954,17'd39693,17'd45955,17'd45956,17'd45957,17'd44682,17'd45958,17'd45959,17'd45960,17'd45961,17'd45962,17'd42576,17'd41212,17'd45223,17'd40797,17'd45963,17'd45964,17'd45965,17'd45966,17'd45967,17'd45968,17'd45969,17'd45970,17'd45971,17'd45972,17'd45973,17'd45974,17'd33915,17'd34076,17'd36385,17'd38391,17'd36244,17'd36384,17'd36670,17'd36669,17'd37227,17'd36661,17'd37368,17'd39720,17'd43826,17'd39720,17'd45975,17'd45976,17'd37096,17'd45258,17'd43411,17'd45977,17'd45978,17'd45979,17'd45980,17'd45981,17'd45982,17'd45151,17'd45983,17'd45871,17'd44354,17'd45984,17'd45152,17'd45481,17'd44362,17'd43701,17'd42600,17'd43298,17'd44823,17'd45873,17'd44106,17'd25567,17'd25568,17'd27637,17'd28254,17'd25029,17'd24896,17'd24742,17'd29241,17'd39133,17'd22860,17'd45985,17'd41586,17'd22157,17'd23573,17'd37116,17'd23566,17'd28722,17'd25030,17'd25709,17'd26064,17'd27146,17'd29379,17'd32016,17'd43289,17'd40822,17'd36983,17'd39437,17'd41429,17'd41110,17'd40367,17'd32832,17'd27761,17'd27761,17'd38537,17'd28726,17'd26901,17'd26782,17'd27259,17'd27515,17'd30734,17'd28717,17'd32007,17'd23732,17'd39278,17'd22677,17'd45986,17'd38041,17'd37659,17'd22680,17'd30128,17'd23565,17'd23731,17'd24898,17'd28720,17'd27515,17'd28725,17'd28486,17'd37513,17'd29246,17'd32496,17'd40959,17'd44358,17'd42299,17'd41864,17'd41418,17'd42886,17'd43560,17'd43434,17'd44593,17'd45987,17'd45369,17'd45988,17'd45989,17'd41417,17'd33790,17'd37908,17'd28486,17'd27259,17'd27638,17'd35735,17'd44367,17'd40523,17'd45990,17'd45991,17'd45992,17'd45993,17'd45994,17'd45995,17'd35321,17'd45996,17'd45997,17'd45998,17'd34638,17'd35455,17'd35865,17'd45999,17'd26528,17'd30879,17'd23922,17'd46000,17'd36139,17'd43986,17'd31496,17'd46001,17'd34879,17'd46002,17'd30620,17'd46003,17'd46004,17'd46005,17'd46006,17'd46007,17'd46008,17'd46009,17'd46010,17'd45899,17'd46011,17'd46012,17'd23281,17'd45902,17'd24802,17'd15476,17'd18620,17'd23463,17'd22250,17'd45776,17'd45903,17'd39771,17'd36310,17'd28186,17'd12622,17'd6221,17'd5005,17'd5145,17'd5604,17'd4363,17'd42631,17'd42464,17'd4357,17'd4359,17'd4358,17'd4017,17'd41458,17'd33532,17'd4683,17'd5156,17'd5156,17'd4999,17'd33839,17'd42772,17'd46013,17'd37147,17'd46014,17'd44011,17'd5600,17'd7320,17'd43589,17'd43869,17'd6061,17'd46015,17'd43870,17'd46016,17'd46017,17'd46018,17'd46019,17'd46020,17'd45651,17'd44963,17'd3047,17'd45910,17'd2881,17'd43327,17'd2531,17'd2892,17'd45514,17'd5772,17'd46021,17'd45787,17'd10649,17'd11188,17'd39181,17'd39483,17'd41481,17'd38072,17'd13176,17'd16492,17'd16492,17'd6418,17'd6418,17'd35769,17'd7537,17'd8507,17'd35769,17'd6258,17'd6258,17'd4713,17'd4085,17'd5630,17'd5940,17'd5631,17'd2394,17'd2560,17'd29440,17'd196,17'd947,17'd10396,17'd46022
},
'{
17'd46023,17'd31905,17'd5200,17'd10532,17'd6263,17'd4888,17'd4892,17'd15746,17'd17917,17'd466,17'd2,17'd2,17'd1416,17'd17,17'd653,17'd653,17'd980,17'd1278,17'd653,17'd809,17'd3254,17'd16866,17'd45516,17'd2262,17'd1973,17'd1973,17'd1702,17'd1282,17'd19499,17'd19609,17'd826,17'd667,17'd17079,17'd46024,17'd2797,17'd3447,17'd37173,17'd15123,17'd44620,17'd29619,17'd24516,17'd25394,17'd30656,17'd29763,17'd46025,17'd16765,17'd13969,17'd13969,17'd19382,17'd17689,17'd17205,17'd18174,17'd18774,17'd39797,17'd34359,17'd39490,17'd46026,17'd46027,17'd46028,17'd46029,17'd36917,17'd46030,17'd40568,17'd38344,17'd37315,17'd35355,17'd46031,17'd31421,17'd46032,17'd46033,17'd30958,17'd9701,17'd8687,17'd12535,17'd9006,17'd13212,17'd4927,17'd4926,17'd4127,17'd6933,17'd7093,17'd42060,17'd6480,17'd45667,17'd40581,17'd44631,17'd46034,17'd43073,17'd6162,17'd46035,17'd44284,17'd40278,17'd46036,17'd46037,17'd46038,17'd46039,17'd46040,17'd46041,17'd45927,17'd46042,17'd46043,17'd46044,17'd46045,17'd46046,17'd46047,17'd46048,17'd7944,17'd46049,17'd38496,17'd8720,17'd10175,17'd16552,17'd10173,17'd9344,17'd10173,17'd10335,17'd9743,17'd13370,17'd13522,17'd11525,17'd17478,17'd24362,17'd25925,17'd25927,17'd26872,17'd26370,17'd26493,17'd24857,17'd28105,17'd24031,17'd22818,17'd18198,17'd15053,17'd18806,17'd18557,17'd20314,17'd24208,17'd26149,17'd26371,17'd27483,17'd25526,17'd26494,17'd24539,17'd28109,17'd46050,17'd23337,17'd28821,17'd11525,17'd17847,17'd9741,17'd17011,17'd10742,17'd9479,17'd9480,17'd10992,17'd12116,17'd11135,17'd10479,17'd11134,17'd10741,17'd46051,17'd40139,17'd18561,17'd33419,17'd31141,17'd37858,17'd36492,17'd33415,17'd32445,17'd13512,17'd18447,17'd10736,17'd16320,17'd16908,17'd45935,17'd46052,17'd45817,17'd41039,17'd45936,17'd46053,17'd45690,17'd45821,17'd46054,17'd46055,17'd40452,17'd40610,17'd45822,17'd46056,17'd45825,17'd46057,17'd46058,17'd46059,17'd46060,17'd46061,17'd46062,17'd46063,17'd46064,17'd46065,17'd46066,17'd46067,17'd46068,17'd46069,17'd46070,17'd46071,17'd46072,17'd40654,17'd46073,17'd43531,17'd44427,17'd46074,17'd46075,17'd46076,17'd46077,17'd45585,17'd46078,17'd46079,17'd42130,17'd45223,17'd43268,17'd46080,17'd46081,17'd46082,17'd46083,17'd46084,17'd38946,17'd46085,17'd46085,17'd46086,17'd46087,17'd33911,17'd46088,17'd40501,17'd40033,17'd40945,17'd35406,17'd39116,17'd37634,17'd36669,17'd38391,17'd37634,17'd39720,17'd37366,17'd37094,17'd37229,17'd37634,17'd38958,17'd43274,17'd39567,17'd36812,17'd37092,17'd37366,17'd39415,17'd35971,17'd39568,17'd46089,17'd46090,17'd46091,17'd46092,17'd44820,17'd45262,17'd45035,17'd44100,17'd44354,17'd45984,17'd45264,17'd46093,17'd43974,17'd44357,17'd44235,17'd46094,17'd43021,17'd44823,17'd46095,17'd28369,17'd27512,17'd28254,17'd25029,17'd28254,17'd24896,17'd24742,17'd29241,17'd46096,17'd32660,17'd46097,17'd46098,17'd31496,17'd30276,17'd29974,17'd23385,17'd34467,17'd27637,17'd25567,17'd27766,17'd27146,17'd31503,17'd30735,17'd43559,17'd41863,17'd41731,17'd31503,17'd36983,17'd34450,17'd40367,17'd32832,17'd27885,17'd30279,17'd44703,17'd34767,17'd26901,17'd26782,17'd27259,17'd26174,17'd28599,17'd25177,17'd25032,17'd23732,17'd29973,17'd22332,17'd46099,17'd32345,17'd31343,17'd22680,17'd32191,17'd23565,17'd23731,17'd25030,17'd28723,17'd27515,17'd28725,17'd28486,17'd29246,17'd31352,17'd33309,17'd43016,17'd46100,17'd46101,17'd46102,17'd46103,17'd44104,17'd44938,17'd44698,17'd44828,17'd46104,17'd46105,17'd45988,17'd45989,17'd41417,17'd33790,17'd37908,17'd30586,17'd26903,17'd25567,17'd30446,17'd34124,17'd32350,17'd46106,17'd46107,17'd46108,17'd46109,17'd46110,17'd46111,17'd46112,17'd46113,17'd46114,17'd44939,17'd33479,17'd39747,17'd35865,17'd45163,17'd45999,17'd24902,17'd23565,17'd34298,17'd46115,17'd22502,17'd31829,17'd34878,17'd41727,17'd46116,17'd46117,17'd46118,17'd46119,17'd46120,17'd46121,17'd46122,17'd46008,17'd46123,17'd46124,17'd45899,17'd46125,17'd45901,17'd46126,17'd45641,17'd24802,17'd17904,17'd18620,17'd23463,17'd39162,17'd38438,17'd39013,17'd36734,17'd36028,17'd28059,17'd12622,17'd5919,17'd4687,17'd4681,17'd43584,17'd4363,17'd42772,17'd39313,17'd4357,17'd4359,17'd4833,17'd4357,17'd41612,17'd4997,17'd4683,17'd4683,17'd4839,17'd4836,17'd4515,17'd4185,17'd5475,17'd6206,17'd33526,17'd42465,17'd5600,17'd46127,17'd12439,17'd4664,17'd46128,17'd46015,17'd40851,17'd46129,17'd46130,17'd46131,17'd46132,17'd38712,17'd45651,17'd44963,17'd34927,17'd45910,17'd46133,17'd46134,17'd46135,17'd2890,17'd41903,17'd5772,17'd46136,17'd10523,17'd10649,17'd11188,17'd5355,17'd39948,17'd41481,17'd38072,17'd13176,17'd16492,17'd16492,17'd6418,17'd6418,17'd6417,17'd7364,17'd8507,17'd8507,17'd6416,17'd8186,17'd4713,17'd4729,17'd5630,17'd14178,17'd15233,17'd27094,17'd1671,17'd1671,17'd195,17'd42923,17'd2920,17'd42648
},
'{
17'd46023,17'd31905,17'd5200,17'd10532,17'd6263,17'd4888,17'd4428,17'd15746,17'd17917,17'd466,17'd0,17'd2,17'd17,17'd17,17'd653,17'd653,17'd980,17'd653,17'd289,17'd809,17'd3254,17'd45516,17'd3103,17'd3103,17'd1973,17'd1973,17'd1702,17'd1282,17'd19499,17'd825,17'd667,17'd827,17'd17079,17'd46024,17'd2797,17'd28434,17'd37173,17'd15123,17'd44620,17'd18526,17'd45188,17'd25394,17'd30656,17'd29621,17'd45406,17'd16765,17'd13969,17'd11764,17'd19382,17'd18774,17'd17205,17'd19891,17'd18774,17'd39797,17'd33859,17'd19389,17'd18780,17'd36053,17'd46137,17'd46137,17'd20295,17'd20430,17'd16415,17'd45523,17'd46138,17'd35496,17'd31920,17'd15013,17'd46139,17'd46140,17'd7410,17'd9701,17'd9158,17'd9005,17'd13212,17'd44630,17'd5254,17'd4926,17'd4127,17'd6933,17'd7094,17'd42060,17'd40874,17'd45667,17'd40581,17'd44631,17'd46034,17'd43073,17'd6162,17'd45668,17'd42354,17'd40278,17'd46141,17'd46037,17'd46038,17'd46142,17'd46143,17'd46041,17'd46144,17'd46042,17'd46043,17'd46145,17'd46146,17'd46147,17'd46148,17'd46149,17'd46150,17'd36932,17'd12118,17'd9040,17'd9194,17'd14811,17'd16328,17'd9480,17'd10334,17'd16328,17'd10026,17'd10172,17'd10332,17'd34205,17'd23513,17'd30229,17'd25925,17'd25927,17'd26872,17'd26370,17'd26493,17'd24857,17'd28105,17'd24031,17'd22818,17'd18198,17'd18917,17'd18806,17'd18557,17'd20314,17'd24208,17'd26493,17'd29196,17'd29196,17'd29640,17'd26756,17'd26372,17'd27985,17'd46151,17'd24540,17'd35799,17'd11525,17'd10331,17'd9884,17'd9741,17'd10742,17'd9479,17'd9480,17'd10992,17'd12116,17'd11276,17'd11276,17'd11134,17'd9883,17'd20044,17'd40602,17'd18446,17'd34049,17'd46152,17'd37858,17'd46153,17'd33579,17'd46154,17'd13512,17'd18447,17'd10736,17'd16320,17'd25812,17'd46155,17'd46156,17'd45817,17'd41039,17'd46157,17'd46053,17'd45690,17'd41665,17'd45822,17'd46158,17'd46159,17'd40452,17'd46160,17'd39675,17'd45825,17'd46161,17'd46162,17'd46163,17'd46164,17'd46165,17'd46166,17'd46167,17'd46168,17'd46169,17'd46170,17'd46171,17'd46172,17'd44088,17'd39881,17'd46173,17'd46173,17'd46174,17'd40800,17'd46175,17'd46176,17'd46177,17'd46178,17'd46179,17'd46180,17'd46181,17'd46180,17'd46182,17'd46183,17'd46073,17'd46184,17'd46185,17'd45724,17'd46186,17'd46187,17'd46188,17'd46189,17'd33283,17'd46190,17'd46191,17'd46192,17'd46193,17'd36238,17'd37235,17'd35551,17'd40349,17'd40350,17'd39116,17'd37634,17'd37367,17'd36670,17'd36384,17'd44922,17'd46194,17'd37494,17'd37093,17'd36669,17'd36385,17'd38958,17'd39415,17'd37227,17'd37229,17'd37368,17'd36384,17'd40349,17'd39415,17'd46195,17'd46196,17'd46197,17'd46198,17'd46199,17'd46104,17'd43972,17'd44224,17'd44224,17'd45370,17'd44592,17'd39129,17'd43844,17'd43559,17'd43289,17'd45484,17'd46200,17'd43021,17'd44230,17'd27882,17'd28480,17'd28719,17'd25029,17'd28254,17'd24896,17'd34467,17'd23734,17'd39588,17'd41867,17'd46097,17'd37385,17'd35429,17'd22326,17'd30128,17'd29972,17'd28851,17'd25177,17'd28598,17'd25833,17'd33163,17'd31354,17'd37908,17'd40822,17'd44357,17'd35707,17'd32832,17'd37114,17'd34877,17'd32356,17'd33319,17'd27885,17'd31503,17'd28726,17'd34767,17'd26901,17'd28725,17'd27515,17'd25949,17'd28599,17'd25177,17'd24895,17'd23732,17'd23216,17'd22678,17'd22682,17'd30580,17'd32344,17'd22679,17'd29374,17'd30275,17'd24415,17'd28254,17'd28723,17'd27515,17'd28853,17'd28486,17'd29379,17'd31352,17'd41111,17'd43975,17'd46201,17'd46202,17'd46203,17'd46204,17'd45745,17'd46205,17'd39738,17'd44931,17'd46105,17'd46105,17'd45988,17'd46206,17'd41417,17'd33941,17'd37908,17'd30586,17'd26903,17'd28597,17'd24251,17'd31664,17'd33944,17'd46207,17'd46208,17'd46209,17'd46210,17'd46211,17'd46212,17'd46213,17'd34777,17'd45490,17'd46214,17'd38296,17'd23572,17'd23567,17'd33813,17'd23383,17'd23564,17'd42449,17'd23738,17'd46215,17'd31500,17'd41867,17'd46216,17'd42003,17'd46217,17'd46218,17'd46219,17'd46220,17'd46221,17'd46222,17'd46223,17'd46008,17'd46224,17'd46225,17'd27406,17'd46226,17'd46227,17'd46126,17'd45641,17'd29297,17'd15476,17'd18620,17'd24152,17'd39162,17'd38439,17'd38845,17'd36029,17'd28059,17'd28186,17'd12622,17'd5615,17'd5005,17'd6067,17'd5604,17'd4364,17'd42772,17'd39165,17'd4357,17'd4359,17'd4833,17'd42462,17'd4356,17'd4997,17'd4683,17'd4840,17'd4683,17'd4525,17'd4358,17'd4016,17'd46228,17'd37147,17'd46229,17'd33833,17'd46230,17'd46127,17'd45647,17'd12439,17'd46231,17'd33529,17'd46232,17'd42036,17'd46233,17'd3361,17'd46234,17'd46235,17'd46236,17'd46237,17'd34927,17'd45910,17'd46133,17'd2717,17'd46135,17'd3057,17'd46238,17'd5024,17'd46021,17'd46239,17'd43462,17'd11188,17'd39181,17'd39483,17'd41481,17'd38072,17'd13176,17'd16492,17'd16492,17'd6418,17'd6418,17'd6417,17'd7364,17'd8507,17'd8507,17'd6416,17'd8186,17'd4713,17'd4729,17'd5630,17'd14178,17'd15233,17'd27094,17'd1671,17'd1671,17'd195,17'd42482,17'd9671,17'd46240
},
'{
17'd46023,17'd31905,17'd30047,17'd10532,17'd10532,17'd44617,17'd4428,17'd14743,17'd46241,17'd12647,17'd0,17'd2,17'd17,17'd17,17'd3905,17'd3905,17'd980,17'd980,17'd653,17'd809,17'd3254,17'd46242,17'd46243,17'd3103,17'd1973,17'd1973,17'd1702,17'd1282,17'd19499,17'd19609,17'd826,17'd827,17'd17079,17'd46024,17'd2797,17'd28434,17'd37173,17'd15123,17'd44620,17'd28666,17'd24010,17'd25800,17'd46244,17'd29621,17'd45406,17'd16765,17'd11764,17'd12532,17'd19892,17'd27461,17'd17205,17'd46245,17'd18655,17'd28925,17'd27458,17'd39043,17'd20026,17'd46246,17'd46247,17'd18889,17'd19894,17'd46248,17'd14631,17'd14898,17'd46249,17'd32418,17'd15142,17'd46250,17'd46139,17'd46251,17'd7248,17'd9573,17'd12219,17'd9006,17'd46252,17'd13212,17'd4927,17'd5254,17'd6306,17'd5085,17'd7914,17'd6474,17'd6633,17'd40580,17'd41329,17'd44631,17'd46034,17'd43073,17'd46253,17'd46254,17'd44284,17'd40278,17'd46255,17'd46256,17'd37844,17'd46257,17'd46258,17'd46259,17'd46260,17'd46261,17'd46262,17'd45806,17'd46263,17'd44529,17'd44873,17'd46264,17'd46265,17'd46266,17'd10607,17'd9348,17'd9041,17'd10174,17'd9480,17'd9480,17'd17232,17'd10334,17'd16328,17'd10333,17'd13522,17'd11525,17'd14382,17'd30229,17'd25925,17'd24856,17'd25927,17'd25927,17'd26149,17'd24538,17'd26371,17'd24031,17'd25926,17'd22992,17'd18917,17'd18806,17'd18557,17'd20314,17'd24030,17'd24856,17'd29065,17'd27621,17'd27483,17'd26756,17'd24705,17'd24992,17'd27860,17'd14259,17'd12583,17'd28463,17'd19280,17'd9883,17'd9741,17'd9885,17'd11809,17'd9480,17'd9620,17'd11809,17'd11277,17'd11277,17'd12116,17'd9740,17'd46267,17'd40288,17'd32137,17'd38370,17'd30381,17'd46268,17'd46269,17'd33582,17'd46154,17'd18807,17'd18447,17'd11519,17'd10739,17'd10606,17'd46270,17'd46271,17'd45817,17'd41039,17'd46272,17'd46273,17'd46274,17'd46275,17'd46276,17'd31972,17'd46159,17'd40147,17'd46277,17'd46278,17'd46279,17'd46280,17'd46281,17'd46282,17'd46283,17'd46284,17'd46285,17'd46286,17'd46287,17'd46288,17'd46285,17'd46289,17'd46290,17'd46291,17'd46292,17'd46293,17'd46294,17'd46295,17'd39230,17'd46296,17'd46297,17'd46298,17'd42421,17'd46299,17'd40304,17'd46300,17'd46301,17'd46302,17'd46303,17'd46304,17'd33281,17'd46305,17'd46306,17'd46307,17'd46308,17'd46309,17'd46310,17'd46311,17'd46312,17'd33913,17'd46313,17'd46314,17'd35406,17'd40349,17'd38391,17'd36670,17'd36669,17'd37634,17'd36669,17'd38391,17'd36660,17'd36819,17'd46315,17'd37494,17'd46316,17'd37092,17'd36813,17'd36384,17'd39720,17'd39416,17'd37366,17'd37096,17'd44922,17'd35971,17'd36813,17'd39416,17'd46317,17'd46318,17'd46319,17'd46320,17'd46321,17'd45879,17'd44100,17'd44224,17'd44224,17'd44936,17'd46093,17'd41416,17'd43844,17'd44103,17'd42436,17'd46200,17'd40825,17'd46200,17'd44230,17'd27511,17'd33803,17'd33803,17'd27764,17'd28254,17'd24896,17'd34467,17'd38980,17'd22325,17'd46322,17'd22167,17'd31829,17'd22857,17'd33158,17'd29374,17'd28722,17'd25030,17'd27511,17'd27638,17'd28978,17'd35011,17'd31353,17'd34451,17'd46323,17'd43552,17'd35570,17'd39910,17'd41274,17'd37658,17'd31354,17'd33319,17'd30279,17'd27642,17'd34767,17'd33963,17'd26902,17'd27259,17'd27515,17'd27766,17'd33000,17'd25178,17'd28851,17'd23918,17'd37117,17'd22678,17'd22505,17'd32660,17'd22332,17'd32827,17'd29374,17'd23732,17'd23916,17'd25178,17'd25566,17'd27515,17'd28853,17'd28486,17'd31352,17'd35426,17'd40959,17'd45745,17'd46324,17'd46325,17'd46326,17'd46324,17'd46327,17'd44226,17'd41862,17'd43972,17'd45262,17'd46105,17'd46328,17'd46329,17'd42889,17'd36264,17'd35426,17'd26901,17'd27515,17'd33000,17'd24088,17'd37673,17'd44491,17'd46330,17'd46331,17'd46332,17'd46333,17'd31228,17'd46334,17'd46335,17'd46336,17'd46337,17'd46338,17'd38296,17'd23572,17'd30579,17'd23212,17'd26656,17'd23565,17'd23566,17'd44715,17'd23570,17'd32999,17'd41865,17'd33947,17'd46339,17'd46340,17'd46341,17'd46342,17'd25839,17'd46343,17'd46344,17'd46345,17'd46346,17'd45771,17'd46347,17'd24631,17'd46348,17'd45901,17'd46126,17'd44955,17'd29297,17'd15476,17'd18620,17'd18619,17'd39161,17'd39013,17'd37556,17'd36030,17'd12761,17'd12761,17'd14301,17'd5614,17'd4686,17'd4681,17'd5604,17'd4364,17'd42772,17'd39165,17'd4357,17'd4359,17'd4362,17'd4364,17'd4356,17'd4997,17'd4840,17'd4840,17'd4839,17'd34155,17'd4833,17'd4016,17'd36165,17'd6206,17'd46229,17'd5473,17'd46230,17'd45510,17'd6061,17'd11826,17'd46231,17'd45177,17'd46349,17'd40708,17'd46350,17'd38065,17'd46351,17'd46352,17'd44962,17'd45652,17'd3194,17'd45910,17'd45183,17'd42475,17'd46353,17'd3057,17'd41904,17'd7680,17'd46136,17'd46354,17'd18629,17'd11188,17'd11048,17'd38202,17'd41481,17'd38072,17'd13420,17'd16492,17'd16492,17'd6418,17'd6418,17'd6417,17'd7364,17'd8507,17'd35769,17'd8186,17'd8186,17'd4713,17'd4729,17'd5630,17'd2098,17'd15233,17'd27094,17'd1671,17'd196,17'd195,17'd42335,17'd46355,17'd46356
},
'{
17'd46023,17'd46357,17'd30047,17'd10532,17'd10532,17'd4889,17'd4428,17'd14743,17'd46241,17'd12647,17'd0,17'd0,17'd17,17'd17,17'd3905,17'd3905,17'd980,17'd652,17'd289,17'd809,17'd2940,17'd45516,17'd46358,17'd3103,17'd1973,17'd1973,17'd1702,17'd1282,17'd19499,17'd825,17'd667,17'd827,17'd17079,17'd46024,17'd2797,17'd28434,17'd37173,17'd15123,17'd44620,17'd28666,17'd24010,17'd25800,17'd46244,17'd46359,17'd45406,17'd29048,17'd12532,17'd12532,17'd18655,17'd17206,17'd17318,17'd25395,17'd18655,17'd20886,17'd24347,17'd46360,17'd20152,17'd20294,17'd46361,17'd46362,17'd19514,17'd46363,17'd39044,17'd15014,17'd36918,17'd46364,17'd31576,17'd46365,17'd31919,17'd14627,17'd6929,17'd46366,17'd9159,17'd9006,17'd46252,17'd44630,17'd5254,17'd5254,17'd6306,17'd4924,17'd7584,17'd6474,17'd6639,17'd46367,17'd46368,17'd44631,17'd46034,17'd43073,17'd46253,17'd46369,17'd42354,17'd40278,17'd46255,17'd46370,17'd46371,17'd46372,17'd46373,17'd46259,17'd46260,17'd46374,17'd46375,17'd46376,17'd45540,17'd44529,17'd44979,17'd46377,17'd46378,17'd46379,17'd8572,17'd8878,17'd9041,17'd17480,17'd10334,17'd17965,17'd37607,17'd17232,17'd46380,17'd46381,17'd33725,17'd34205,17'd36348,17'd27985,17'd28110,17'd24856,17'd25927,17'd25927,17'd26149,17'd24538,17'd26371,17'd24031,17'd25926,17'd22992,17'd18917,17'd18806,17'd18557,17'd20314,17'd24707,17'd27004,17'd29327,17'd32435,17'd32759,17'd46382,17'd26756,17'd24538,17'd46383,17'd24363,17'd36481,17'd38499,17'd11525,17'd10329,17'd10024,17'd9885,17'd9479,17'd9620,17'd9620,17'd9479,17'd12116,17'd11277,17'd9741,17'd10856,17'd46267,17'd40288,17'd42677,17'd38370,17'd30381,17'd46384,17'd37858,17'd33736,17'd46154,17'd18807,17'd18447,17'd11519,17'd10739,17'd10479,17'd46385,17'd46271,17'd46386,17'd46387,17'd46272,17'd46273,17'd46274,17'd45822,17'd46388,17'd46389,17'd39838,17'd40147,17'd46390,17'd42083,17'd46391,17'd46280,17'd46392,17'd46282,17'd46164,17'd46393,17'd46394,17'd46395,17'd46396,17'd46397,17'd46398,17'd35125,17'd46399,17'd46400,17'd46401,17'd46402,17'd46403,17'd46404,17'd39563,17'd46405,17'd46406,17'd46407,17'd46065,17'd46171,17'd46408,17'd43822,17'd46409,17'd46191,17'd46410,17'd46411,17'd46310,17'd46412,17'd46413,17'd46413,17'd40347,17'd46414,17'd46415,17'd46416,17'd44578,17'd44689,17'd35962,17'd35551,17'd35962,17'd36244,17'd36669,17'd36244,17'd36670,17'd37634,17'd36670,17'd36244,17'd36668,17'd38130,17'd46417,17'd46417,17'd37095,17'd39569,17'd39116,17'd36384,17'd39567,17'd46418,17'd39412,17'd37096,17'd38006,17'd38645,17'd37227,17'd46419,17'd46420,17'd46421,17'd46422,17'd46423,17'd43420,17'd46424,17'd45263,17'd44354,17'd44224,17'd45609,17'd39434,17'd41997,17'd44357,17'd44227,17'd42741,17'd46425,17'd40959,17'd42886,17'd46426,17'd27511,17'd33803,17'd33803,17'd27764,17'd25030,17'd24744,17'd23917,17'd46427,17'd22681,17'd46428,17'd46428,17'd37659,17'd22680,17'd29974,17'd29529,17'd24252,17'd27637,17'd25317,17'd27513,17'd27258,17'd37908,17'd30735,17'd46429,17'd46430,17'd43560,17'd36127,17'd45613,17'd41274,17'd42890,17'd31503,17'd27885,17'd27642,17'd29379,17'd46431,17'd35023,17'd26782,17'd27640,17'd27514,17'd28602,17'd31366,17'd25178,17'd24416,17'd23918,17'd37117,17'd39131,17'd33311,17'd35296,17'd30276,17'd23389,17'd29686,17'd24086,17'd24416,17'd25568,17'd25708,17'd27259,17'd26782,17'd28486,17'd31352,17'd37908,17'd41271,17'd46432,17'd46433,17'd46434,17'd46435,17'd46436,17'd46437,17'd39903,17'd44697,17'd46438,17'd46439,17'd45369,17'd46440,17'd46441,17'd38975,17'd38025,17'd31352,17'd26781,17'd27514,17'd28717,17'd24089,17'd46442,17'd46443,17'd46444,17'd46445,17'd46446,17'd30015,17'd46447,17'd46448,17'd46449,17'd46450,17'd46113,17'd46451,17'd46443,17'd43292,17'd23569,17'd46452,17'd23211,17'd29099,17'd38668,17'd36139,17'd46453,17'd46454,17'd42001,17'd41727,17'd46455,17'd46456,17'd46457,17'd46342,17'd46458,17'd46459,17'd46460,17'd31865,17'd46461,17'd45771,17'd46462,17'd46463,17'd46348,17'd46464,17'd46126,17'd44955,17'd24945,17'd15476,17'd19590,17'd37940,17'd43581,17'd38845,17'd37428,17'd41141,17'd12906,17'd16615,17'd12467,17'd27935,17'd4842,17'd6067,17'd40079,17'd42462,17'd42772,17'd39165,17'd4357,17'd4359,17'd4359,17'd42462,17'd4356,17'd4997,17'd4840,17'd4840,17'd4683,17'd5000,17'd4833,17'd4831,17'd46228,17'd37147,17'd46229,17'd5473,17'd46465,17'd5318,17'd6061,17'd46466,17'd46467,17'd46468,17'd46469,17'd46470,17'd46471,17'd37950,17'd46351,17'd46472,17'd46473,17'd46474,17'd3194,17'd45782,17'd45183,17'd42475,17'd46475,17'd46476,17'd41904,17'd7680,17'd45786,17'd46477,17'd41003,17'd11188,17'd39790,17'd38859,17'd41481,17'd38203,17'd13420,17'd37959,17'd37959,17'd6418,17'd6418,17'd6417,17'd7364,17'd8507,17'd35769,17'd8186,17'd8186,17'd4882,17'd4729,17'd5940,17'd14586,17'd15233,17'd777,17'd196,17'd196,17'd195,17'd46478,17'd2117,17'd46479
},
'{
17'd46023,17'd46357,17'd30047,17'd5053,17'd46480,17'd4889,17'd4088,17'd15746,17'd15357,17'd15495,17'd2,17'd2,17'd17,17'd17,17'd3905,17'd3905,17'd27,17'd4430,17'd289,17'd30,17'd982,17'd1130,17'd46358,17'd3103,17'd1973,17'd2122,17'd1702,17'd1557,17'd19499,17'd19609,17'd992,17'd18991,17'd18150,17'd1561,17'd2797,17'd28434,17'd46481,17'd41910,17'd44743,17'd28666,17'd24010,17'd25800,17'd30954,17'd46482,17'd45406,17'd29048,17'd12532,17'd18884,17'd27461,17'd17206,17'd17572,17'd18656,17'd19511,17'd19006,17'd24347,17'd34181,17'd35068,17'd19134,17'd45070,17'd28925,17'd46483,17'd19624,17'd18537,17'd46484,17'd15904,17'd46485,17'd46486,17'd46487,17'd46488,17'd6134,17'd6929,17'd9702,17'd9159,17'd10694,17'd12534,17'd10430,17'd9302,17'd5254,17'd6306,17'd4924,17'd7253,17'd7754,17'd40873,17'd46489,17'd46490,17'd46491,17'd46492,17'd43204,17'd46493,17'd46494,17'd43892,17'd40124,17'd46495,17'd38101,17'd46496,17'd46497,17'd46498,17'd46499,17'd46500,17'd46501,17'd46375,17'd46502,17'd45806,17'd46503,17'd45304,17'd46504,17'd46505,17'd8417,17'd8571,17'd8725,17'd9348,17'd8874,17'd9742,17'd18556,17'd37607,17'd17717,17'd26875,17'd10333,17'd13369,17'd13368,17'd36348,17'd30229,17'd25925,17'd24537,17'd25927,17'd27123,17'd26149,17'd24031,17'd26149,17'd24208,17'd20450,17'd22992,17'd16325,17'd15185,17'd12582,17'd18559,17'd23512,17'd27004,17'd28816,17'd29923,17'd30369,17'd30219,17'd46382,17'd25526,17'd24538,17'd24362,17'd23513,17'd37196,17'd12423,17'd11526,17'd10169,17'd9885,17'd9479,17'd9480,17'd9620,17'd9480,17'd9619,17'd9619,17'd12116,17'd9473,17'd9611,17'd46051,17'd41511,17'd37859,17'd46506,17'd46507,17'd36356,17'd32608,17'd32604,17'd12717,17'd11805,17'd28696,17'd10477,17'd29199,17'd46508,17'd46509,17'd45310,17'd46387,17'd46272,17'd46273,17'd46274,17'd46054,17'd32153,17'd46510,17'd46511,17'd36224,17'd46512,17'd46513,17'd46279,17'd34413,17'd46514,17'd46282,17'd46515,17'd46516,17'd46517,17'd40500,17'd46518,17'd46519,17'd46398,17'd46520,17'd35396,17'd35396,17'd46521,17'd46522,17'd46523,17'd46524,17'd46525,17'd46526,17'd46526,17'd46527,17'd38936,17'd46528,17'd40660,17'd43135,17'd42580,17'd46529,17'd46530,17'd45859,17'd46531,17'd46532,17'd46533,17'd46534,17'd46535,17'd46536,17'd34591,17'd44689,17'd46537,17'd43004,17'd46538,17'd43411,17'd46539,17'd46540,17'd36670,17'd39262,17'd35971,17'd36244,17'd36669,17'd37634,17'd36818,17'd38007,17'd38128,17'd46315,17'd37634,17'd38391,17'd39116,17'd36244,17'd39416,17'd38259,17'd46541,17'd39412,17'd39567,17'd39720,17'd37366,17'd44923,17'd46542,17'd46543,17'd46544,17'd46545,17'd42295,17'd44223,17'd44354,17'd44224,17'd44587,17'd43833,17'd44479,17'd43844,17'd44933,17'd46546,17'd46547,17'd43424,17'd41270,17'd41418,17'd46548,17'd29103,17'd46549,17'd46549,17'd25568,17'd25030,17'd24252,17'd32186,17'd46550,17'd31496,17'd22009,17'd46551,17'd37510,17'd22328,17'd37386,17'd23564,17'd24895,17'd25568,17'd28484,17'd27513,17'd33163,17'd37908,17'd32004,17'd42297,17'd46552,17'd39907,17'd35570,17'd35990,17'd37248,17'd33790,17'd31503,17'd30279,17'd27642,17'd28727,17'd35023,17'd26781,17'd26782,17'd27515,17'd25707,17'd28723,17'd28717,17'd27637,17'd30126,17'd34137,17'd33651,17'd22501,17'd22680,17'd22677,17'd22331,17'd36426,17'd35865,17'd24087,17'd24742,17'd28850,17'd25565,17'd28725,17'd26782,17'd32016,17'd31352,17'd37908,17'd44827,17'd46553,17'd46436,17'd46554,17'd46555,17'd46435,17'd46556,17'd40216,17'd46557,17'd42595,17'd46558,17'd45870,17'd46559,17'd46560,17'd33308,17'd35570,17'd31352,17'd33963,17'd27514,17'd27882,17'd36701,17'd40833,17'd46561,17'd46218,17'd46562,17'd46563,17'd46564,17'd46565,17'd46566,17'd46567,17'd35592,17'd46568,17'd44947,17'd46569,17'd34278,17'd32008,17'd30579,17'd35865,17'd29827,17'd23387,17'd46570,17'd30428,17'd33948,17'd35708,17'd46571,17'd46572,17'd46573,17'd46574,17'd46575,17'd46576,17'd46577,17'd46578,17'd46579,17'd46580,17'd45897,17'd46581,17'd19821,17'd23786,17'd46464,17'd23459,17'd46582,17'd37027,17'd22765,17'd22420,17'd18498,17'd43581,17'd37286,17'd22943,17'd36028,17'd12622,17'd12468,17'd15728,17'd27935,17'd4686,17'd4836,17'd41612,17'd4832,17'd42772,17'd39313,17'd33839,17'd4190,17'd4359,17'd4357,17'd33533,17'd4997,17'd4995,17'd4683,17'd4683,17'd4525,17'd34157,17'd4016,17'd36165,17'd6206,17'd46229,17'd41758,17'd46583,17'd4178,17'd33198,17'd46466,17'd43049,17'd46584,17'd46585,17'd3678,17'd46586,17'd46587,17'd46588,17'd46589,17'd45064,17'd46236,17'd46590,17'd2880,17'd46591,17'd37953,17'd46592,17'd46593,17'd46594,17'd46595,17'd10071,17'd46596,17'd41003,17'd40716,17'd38458,17'd38334,17'd41481,17'd38203,17'd13420,17'd16492,17'd16492,17'd16492,17'd16492,17'd6418,17'd6418,17'd8507,17'd35769,17'd8186,17'd8186,17'd4713,17'd5630,17'd16382,17'd16256,17'd2394,17'd1950,17'd417,17'd42786,17'd950,17'd1110,17'd2117,17'd46597
},
'{
17'd46598,17'd46357,17'd30047,17'd5053,17'd46480,17'd4890,17'd4088,17'd15746,17'd15357,17'd15495,17'd2,17'd2,17'd17,17'd17,17'd3905,17'd653,17'd27,17'd4430,17'd289,17'd31,17'd982,17'd983,17'd46358,17'd3103,17'd2939,17'd2122,17'd1702,17'd1557,17'd19499,17'd19609,17'd992,17'd17553,17'd1285,17'd1561,17'd2797,17'd3447,17'd46481,17'd41910,17'd44743,17'd44853,17'd24516,17'd25800,17'd30954,17'd25801,17'd30057,17'd46025,17'd18884,17'd17317,17'd17206,17'd21185,17'd17572,17'd18656,17'd18655,17'd19006,17'd24347,17'd33550,17'd34359,17'd19622,17'd43337,17'd20886,17'd34358,17'd46599,17'd36189,17'd16884,17'd15647,17'd34677,17'd31576,17'd46600,17'd46601,17'd6134,17'd6300,17'd13471,17'd9703,17'd10694,17'd12534,17'd10430,17'd9302,17'd5254,17'd6627,17'd4924,17'd7089,17'd7254,17'd7915,17'd39647,17'd6482,17'd46491,17'd46492,17'd43204,17'd46493,17'd46602,17'd43075,17'd40124,17'd46495,17'd46603,17'd46604,17'd46497,17'd46498,17'd46605,17'd46606,17'd46607,17'd46608,17'd46609,17'd46376,17'd46610,17'd45304,17'd46611,17'd46612,17'd19780,17'd24545,17'd24368,17'd8886,17'd10175,17'd26875,17'd17841,17'd46613,17'd17717,17'd17717,17'd10171,17'd46614,17'd13368,17'd36348,17'd27985,17'd28110,17'd24537,17'd25927,17'd25927,17'd26149,17'd24031,17'd26149,17'd28231,17'd20608,17'd22992,17'd16325,17'd15185,17'd12582,17'd18559,17'd24030,17'd26370,17'd28343,17'd29923,17'd30369,17'd46615,17'd46616,17'd29640,17'd26493,17'd24031,17'd33084,17'd30230,17'd11668,17'd19280,17'd10024,17'd9885,17'd9479,17'd9480,17'd9620,17'd9480,17'd17011,17'd9619,17'd12116,17'd9885,17'd27003,17'd46051,17'd46617,17'd37987,17'd46506,17'd46507,17'd37858,17'd32448,17'd32603,17'd12717,17'd11805,17'd10735,17'd14518,17'd25530,17'd46618,17'd46619,17'd45817,17'd46620,17'd46621,17'd46622,17'd46623,17'd45822,17'd46055,17'd37992,17'd36084,17'd36224,17'd46512,17'd46513,17'd46391,17'd46624,17'd44425,17'd46282,17'd46625,17'd46626,17'd46627,17'd46628,17'd46629,17'd46414,17'd46414,17'd46630,17'd46631,17'd46632,17'd46633,17'd46634,17'd46635,17'd46634,17'd46636,17'd46637,17'd46638,17'd46639,17'd37493,17'd45471,17'd40033,17'd46313,17'd46640,17'd46640,17'd46313,17'd33766,17'd46641,17'd46642,17'd46643,17'd46644,17'd46645,17'd46646,17'd35274,17'd35835,17'd46647,17'd46648,17'd43534,17'd46539,17'd46649,17'd46650,17'd43412,17'd38262,17'd38645,17'd36244,17'd37366,17'd37095,17'd38007,17'd37763,17'd46541,17'd39412,17'd38391,17'd38391,17'd36813,17'd36669,17'd39412,17'd46651,17'd46315,17'd39416,17'd39567,17'd39415,17'd44922,17'd46652,17'd46653,17'd46654,17'd46655,17'd46656,17'd42879,17'd44100,17'd44354,17'd44224,17'd46657,17'd43833,17'd46658,17'd43701,17'd44938,17'd43834,17'd44823,17'd43548,17'd43548,17'd41864,17'd46659,17'd29244,17'd46549,17'd31856,17'd27512,17'd25030,17'd34467,17'd29528,17'd39588,17'd31496,17'd22164,17'd22165,17'd32344,17'd23218,17'd29975,17'd30879,17'd25030,17'd28717,17'd25567,17'd26064,17'd32016,17'd39437,17'd33308,17'd46552,17'd42882,17'd40520,17'd35291,17'd35150,17'd37248,17'd36264,17'd30279,17'd30279,17'd27642,17'd28979,17'd35023,17'd33963,17'd26782,17'd27514,17'd25833,17'd28720,17'd28717,17'd25180,17'd35159,17'd23384,17'd32352,17'd33158,17'd22680,17'd22680,17'd22331,17'd30425,17'd29099,17'd24249,17'd24744,17'd28369,17'd25833,17'd26782,17'd26781,17'd31353,17'd29379,17'd33791,17'd44700,17'd46660,17'd46661,17'd46662,17'd46663,17'd46664,17'd46665,17'd43546,17'd42296,17'd41995,17'd46666,17'd46667,17'd46668,17'd45266,17'd33476,17'd35570,17'd29245,17'd26782,17'd25949,17'd25177,17'd35999,17'd46669,17'd46670,17'd46218,17'd46671,17'd46672,17'd46564,17'd46673,17'd46674,17'd46567,17'd35592,17'd46675,17'd45761,17'd46569,17'd44591,17'd33158,17'd29974,17'd30579,17'd23387,17'd34124,17'd45040,17'd46676,17'd46677,17'd41422,17'd46678,17'd46679,17'd46680,17'd46681,17'd46682,17'd46683,17'd21091,17'd46684,17'd46685,17'd46580,17'd45897,17'd46686,17'd19469,17'd46687,17'd46688,17'd6383,17'd46689,17'd24802,17'd15340,17'd26585,17'd22942,17'd37940,17'd37286,17'd22943,17'd28059,17'd12622,17'd14050,17'd35609,17'd28185,17'd4686,17'd4836,17'd41458,17'd4357,17'd39165,17'd44258,17'd33839,17'd4190,17'd4359,17'd4515,17'd39468,17'd38442,17'd4995,17'd4683,17'd4683,17'd4525,17'd34157,17'd4831,17'd46013,17'd37147,17'd34151,17'd4351,17'd42465,17'd33527,17'd33198,17'd46466,17'd46690,17'd46691,17'd41151,17'd46692,17'd46693,17'd46694,17'd46588,17'd46695,17'd46696,17'd46697,17'd3194,17'd2880,17'd46591,17'd37953,17'd46592,17'd46476,17'd46698,17'd46595,17'd45656,17'd46477,17'd41003,17'd40716,17'd39790,17'd38859,17'd38334,17'd38203,17'd13420,17'd16492,17'd16492,17'd16492,17'd16492,17'd6418,17'd6418,17'd8507,17'd35769,17'd8186,17'd8186,17'd4882,17'd5630,17'd16382,17'd14586,17'd28428,17'd1950,17'd417,17'd417,17'd13573,17'd950,17'd1381,17'd46699
},
'{
17'd46598,17'd31905,17'd30047,17'd5053,17'd46700,17'd4735,17'd4088,17'd15746,17'd2594,17'd2595,17'd2,17'd2,17'd17,17'd17,17'd653,17'd652,17'd27,17'd652,17'd289,17'd31,17'd982,17'd983,17'd984,17'd13303,17'd2939,17'd1973,17'd1702,17'd1557,17'd19499,17'd19609,17'd826,17'd992,17'd35772,17'd1708,17'd13072,17'd3447,17'd46481,17'd42198,17'd46701,17'd28666,17'd24010,17'd25800,17'd46702,17'd25801,17'd30057,17'd28667,17'd12532,17'd17317,17'd19255,17'd19255,17'd17572,17'd17572,17'd18655,17'd20292,17'd13211,17'd34180,17'd9433,17'd43599,17'd29048,17'd16765,17'd34015,17'd46703,17'd19623,17'd36053,17'd46704,17'd46705,17'd46706,17'd46707,17'd46708,17'd14221,17'd6134,17'd9300,17'd9703,17'd9703,17'd12534,17'd12534,17'd9302,17'd4927,17'd4926,17'd4610,17'd6933,17'd7096,17'd6780,17'd46709,17'd46710,17'd46491,17'd46492,17'd43073,17'd46253,17'd46494,17'd43892,17'd40124,17'd46495,17'd46711,17'd46712,17'd46713,17'd46714,17'd46605,17'd46606,17'd46715,17'd46716,17'd46609,17'd46717,17'd46045,17'd46718,17'd46719,17'd46720,17'd8251,17'd23173,17'd31759,17'd8879,17'd9043,17'd9742,17'd16561,17'd46613,17'd37607,17'd46721,17'd46722,17'd28688,17'd28821,17'd36348,17'd30229,17'd25925,17'd24537,17'd25927,17'd25927,17'd26149,17'd27122,17'd26149,17'd28231,17'd20608,17'd19920,17'd15185,17'd15185,17'd12582,17'd17722,17'd24030,17'd26370,17'd29923,17'd30831,17'd29066,17'd30218,17'd30525,17'd27346,17'd29196,17'd24857,17'd26150,17'd44982,17'd18326,17'd11669,17'd26152,17'd10856,17'd10742,17'd10743,17'd9620,17'd9480,17'd17011,17'd9619,17'd17011,17'd10742,17'd27003,17'd46267,17'd46723,17'd39663,17'd46506,17'd46724,17'd46725,17'd31778,17'd43083,17'd12412,17'd21982,17'd29332,17'd15943,17'd15431,17'd46726,17'd46727,17'd39983,17'd46728,17'd46729,17'd46730,17'd46055,17'd46276,17'd46158,17'd36643,17'd46731,17'd36224,17'd46732,17'd46513,17'd46733,17'd46280,17'd46514,17'd46282,17'd46734,17'd46735,17'd46736,17'd46737,17'd46738,17'd46739,17'd46740,17'd46521,17'd46741,17'd46742,17'd46743,17'd35973,17'd46744,17'd45733,17'd46745,17'd43004,17'd34075,17'd42135,17'd42135,17'd36674,17'd36379,17'd42424,17'd42135,17'd42135,17'd34591,17'd34591,17'd40945,17'd33769,17'd46746,17'd46746,17'd46744,17'd46747,17'd35834,17'd36247,17'd36965,17'd39262,17'd39567,17'd39720,17'd38958,17'd39720,17'd39887,17'd39262,17'd39720,17'd44922,17'd37230,17'd37362,17'd37363,17'd37230,17'd37368,17'd37367,17'd36670,17'd38391,17'd36812,17'd37367,17'd46315,17'd39260,17'd37636,17'd46649,17'd39568,17'd45258,17'd43005,17'd46748,17'd38266,17'd46749,17'd46750,17'd46751,17'd43422,17'd44473,17'd44224,17'd44472,17'd45609,17'd46752,17'd43692,17'd44103,17'd46546,17'd43975,17'd42883,17'd46753,17'd46753,17'd42300,17'd43976,17'd25568,17'd33803,17'd33484,17'd28719,17'd24895,17'd30431,17'd31190,17'd36986,17'd31496,17'd22164,17'd22156,17'd30276,17'd23217,17'd29687,17'd32659,17'd25178,17'd33000,17'd28597,17'd25949,17'd36127,17'd36127,17'd41417,17'd46754,17'd39275,17'd33941,17'd34877,17'd35704,17'd35290,17'd36127,17'd27885,17'd30279,17'd31352,17'd26901,17'd35023,17'd26782,17'd27259,17'd27514,17'd26174,17'd28720,17'd25177,17'd25030,17'd23916,17'd23384,17'd29975,17'd32008,17'd32827,17'd22329,17'd22679,17'd23217,17'd23733,17'd32659,17'd24898,17'd28130,17'd26903,17'd35023,17'd26781,17'd31353,17'd27642,17'd33941,17'd43021,17'd46755,17'd46756,17'd46757,17'd46758,17'd46759,17'd46760,17'd39582,17'd42880,17'd41579,17'd46761,17'd46762,17'd46763,17'd46764,17'd33790,17'd31354,17'd29245,17'd27371,17'd28602,17'd28254,17'd23918,17'd45754,17'd46106,17'd46765,17'd46766,17'd46767,17'd46768,17'd46769,17'd46770,17'd46771,17'd46772,17'd46675,17'd46773,17'd46774,17'd45754,17'd36543,17'd23569,17'd23388,17'd23387,17'd23387,17'd46570,17'd34759,17'd22007,17'd35427,17'd46775,17'd46776,17'd46777,17'd46574,17'd46778,17'd33184,17'd25038,17'd46779,17'd40974,17'd46780,17'd46781,17'd46782,17'd20087,17'd29155,17'd11691,17'd25628,17'd46783,17'd37027,17'd23116,17'd22420,17'd16247,17'd22942,17'd36734,17'd19479,17'd27198,17'd24945,17'd12161,17'd15990,17'd5335,17'd4686,17'd4836,17'd41612,17'd4832,17'd4185,17'd39165,17'd4515,17'd4189,17'd4190,17'd4515,17'd33840,17'd30486,17'd5327,17'd5328,17'd4840,17'd5000,17'd33991,17'd4356,17'd46013,17'd37147,17'd34151,17'd4351,17'd42184,17'd33527,17'd46231,17'd46784,17'd46690,17'd46785,17'd40708,17'd46786,17'd46787,17'd3539,17'd37036,17'd46352,17'd46788,17'd46697,17'd46789,17'd46790,17'd44386,17'd37953,17'd46592,17'd45784,17'd4551,17'd7680,17'd41625,17'd46596,17'd18629,17'd40716,17'd11048,17'd38202,17'd38334,17'd38203,17'd38072,17'd44387,17'd43596,17'd16492,17'd16492,17'd6258,17'd6094,17'd8507,17'd35769,17'd8186,17'd8186,17'd5940,17'd5630,17'd16382,17'd15233,17'd2560,17'd2560,17'd417,17'd600,17'd1110,17'd41627,17'd972,17'd46791
},
'{
17'd46792,17'd31905,17'd5200,17'd5053,17'd46700,17'd4735,17'd4088,17'd15746,17'd2594,17'd2595,17'd2,17'd2,17'd17,17'd17,17'd653,17'd652,17'd27,17'd652,17'd289,17'd31,17'd982,17'd984,17'd811,17'd471,17'd2939,17'd2939,17'd1972,17'd1282,17'd46793,17'd46794,17'd826,17'd992,17'd35772,17'd46024,17'd2797,17'd2958,17'd46481,17'd42198,17'd46701,17'd44853,17'd24516,17'd25800,17'd46702,17'd25801,17'd30057,17'd28205,17'd17204,17'd17204,17'd19008,17'd17320,17'd16767,17'd17572,17'd18655,17'd20292,17'd13211,17'd23325,17'd27458,17'd12531,17'd28667,17'd16765,17'd34015,17'd38081,17'd46795,17'd20428,17'd31575,17'd46796,17'd46797,17'd46707,17'd15263,17'd46798,17'd46798,17'd13972,17'd13469,17'd10113,17'd9301,17'd12534,17'd9302,17'd4927,17'd4926,17'd6627,17'd5085,17'd7089,17'd41019,17'd46709,17'd46799,17'd46491,17'd46492,17'd43073,17'd46253,17'd46800,17'd43207,17'd40124,17'd46495,17'd46711,17'd46801,17'd46802,17'd46714,17'd46803,17'd46804,17'd46715,17'd46805,17'd46806,17'd46375,17'd46263,17'd46807,17'd46808,17'd35091,17'd17352,17'd13373,17'd11531,17'd8725,17'd9045,17'd26875,17'd16561,17'd46809,17'd46613,17'd27744,17'd46810,17'd42674,17'd28821,17'd36348,17'd27985,17'd28110,17'd24537,17'd24856,17'd28105,17'd32127,17'd27122,17'd26149,17'd28231,17'd20608,17'd16325,17'd15185,17'd19158,17'd12582,17'd18198,17'd24030,17'd26872,17'd28943,17'd29066,17'd29066,17'd30831,17'd30674,17'd30524,17'd32759,17'd27483,17'd26628,17'd46811,17'd36481,17'd21206,17'd10329,17'd16796,17'd9885,17'd10743,17'd9620,17'd9620,17'd10742,17'd9619,17'd9619,17'd10742,17'd27003,17'd46267,17'd31952,17'd33420,17'd46812,17'd46507,17'd46384,17'd31603,17'd29653,17'd15686,17'd21982,17'd29332,17'd20756,17'd15431,17'd46813,17'd46814,17'd46815,17'd46816,17'd46817,17'd46818,17'd46055,17'd46276,17'd46158,17'd36643,17'd46731,17'd46819,17'd46820,17'd43487,17'd46821,17'd46822,17'd44659,17'd46823,17'd46824,17'd46825,17'd46826,17'd46827,17'd46517,17'd46739,17'd46740,17'd46828,17'd45730,17'd46829,17'd46830,17'd41566,17'd43272,17'd43273,17'd43004,17'd38639,17'd34994,17'd34994,17'd36674,17'd42424,17'd33453,17'd35137,17'd33769,17'd37235,17'd33619,17'd35679,17'd33619,17'd46831,17'd43272,17'd43272,17'd45597,17'd45732,17'd35273,17'd36245,17'd38262,17'd38133,17'd38009,17'd38133,17'd38262,17'd39887,17'd43412,17'd39415,17'd38260,17'd46194,17'd37231,17'd37231,17'd37095,17'd37096,17'd37368,17'd37367,17'd36670,17'd38391,17'd39569,17'd37092,17'd37231,17'd46541,17'd46540,17'd43534,17'd44922,17'd46832,17'd45362,17'd39263,17'd46833,17'd46834,17'd46835,17'd40047,17'd45035,17'd44473,17'd44224,17'd46657,17'd43833,17'd45481,17'd41997,17'd44103,17'd45483,17'd42883,17'd43154,17'd43979,17'd42885,17'd42597,17'd43836,17'd27512,17'd28480,17'd33484,17'd25029,17'd24895,17'd32186,17'd38806,17'd34458,17'd31657,17'd37385,17'd22161,17'd22331,17'd37117,17'd23384,17'd28977,17'd25177,17'd33000,17'd28597,17'd25707,17'd36127,17'd46836,17'd46837,17'd46838,17'd41109,17'd38025,17'd37907,17'd35704,17'd35425,17'd31503,17'd32832,17'd27885,17'd31352,17'd26901,17'd35023,17'd27371,17'd27640,17'd27515,17'd26174,17'd28594,17'd25177,17'd25030,17'd24415,17'd23384,17'd23386,17'd23388,17'd23389,17'd36543,17'd36426,17'd30128,17'd24087,17'd28851,17'd27637,17'd28720,17'd28725,17'd33963,17'd28726,17'd39437,17'd31503,17'd33790,17'd44823,17'd46839,17'd46840,17'd46841,17'd46840,17'd46842,17'd46843,17'd46844,17'd46845,17'd46846,17'd46847,17'd45479,17'd46763,17'd46848,17'd36264,17'd31503,17'd28727,17'd27371,17'd26064,17'd24897,17'd29376,17'd40523,17'd46849,17'd46850,17'd46851,17'd46852,17'd46853,17'd46854,17'd46447,17'd46855,17'd46772,17'd46856,17'd41285,17'd39920,17'd44702,17'd36543,17'd32351,17'd30128,17'd23387,17'd34124,17'd46857,17'd46858,17'd31658,17'd46859,17'd46860,17'd46861,17'd46862,17'd46863,17'd46864,17'd25441,17'd46865,17'd46866,17'd46867,17'd46780,17'd46781,17'd46868,17'd20237,17'd28055,17'd46869,17'd31088,17'd46783,17'd37027,17'd15094,17'd17066,17'd17533,17'd17533,17'd38190,17'd18970,17'd16123,17'd24484,17'd13679,17'd29296,17'd5335,17'd4686,17'd4836,17'd33533,17'd42462,17'd41612,17'd33534,17'd34157,17'd4524,17'd4189,17'd34157,17'd33691,17'd30486,17'd5328,17'd4841,17'd4686,17'd4526,17'd33991,17'd4356,17'd46870,17'd46871,17'd46872,17'd4351,17'd42184,17'd33527,17'd46231,17'd46873,17'd46874,17'd40704,17'd46875,17'd46876,17'd46877,17'd37812,17'd46878,17'd37705,17'd46879,17'd46697,17'd46880,17'd45782,17'd44386,17'd46881,17'd46592,17'd42334,17'd46882,17'd46883,17'd45656,17'd46477,17'd18629,17'd40716,17'd39181,17'd38859,17'd38334,17'd38203,17'd38072,17'd44387,17'd43596,17'd16492,17'd16492,17'd6258,17'd6094,17'd8507,17'd35769,17'd8186,17'd8186,17'd5940,17'd5630,17'd16382,17'd14586,17'd28916,17'd33847,17'd417,17'd196,17'd13809,17'd601,17'd32250,17'd1966
},
'{
17'd4243,17'd4891,17'd5201,17'd5197,17'd5052,17'd5201,17'd3904,17'd15746,17'd2594,17'd466,17'd17,17'd17,17'd17,17'd17,17'd653,17'd652,17'd27,17'd652,17'd289,17'd31,17'd982,17'd983,17'd657,17'd471,17'd2939,17'd2939,17'd1972,17'd16966,17'd46884,17'd46793,17'd46885,17'd992,17'd35772,17'd46024,17'd46886,17'd36606,17'd46887,17'd32412,17'd17308,17'd44853,17'd24516,17'd46888,17'd46702,17'd24518,17'd45406,17'd28667,17'd12681,17'd17204,17'd19008,17'd17320,17'd46889,17'd20425,17'd18774,17'd28667,17'd13211,17'd17096,17'd24347,17'd13969,17'd16658,17'd12361,17'd13093,17'd34938,17'd46890,17'd20888,17'd46891,17'd46892,17'd46893,17'd46707,17'd15771,17'd46798,17'd23670,17'd13972,17'd13470,17'd15138,17'd9301,17'd9007,17'd4611,17'd4767,17'd4926,17'd6627,17'd4924,17'd8375,17'd7100,17'd46894,17'd46895,17'd46896,17'd46897,17'd43073,17'd46253,17'd46898,17'd46899,17'd46900,17'd46901,17'd46711,17'd46801,17'd46902,17'd46903,17'd46904,17'd46905,17'd46906,17'd46907,17'd46908,17'd46608,17'd46044,17'd46909,17'd46910,17'd46911,17'd18203,17'd22993,17'd11405,17'd12264,17'd9044,17'd10025,17'd16561,17'd27006,17'd46809,17'd16561,17'd10332,17'd42674,17'd28821,17'd36348,17'd24208,17'd25925,17'd24537,17'd24856,17'd24856,17'd24538,17'd27122,17'd26149,17'd28231,17'd20608,17'd16325,17'd19158,17'd19158,17'd18917,17'd18198,17'd23512,17'd26370,17'd28943,17'd29066,17'd29329,17'd29066,17'd46912,17'd30218,17'd30524,17'd27346,17'd25526,17'd26258,17'd36626,17'd11668,17'd19280,17'd16796,17'd9741,17'd9885,17'd10743,17'd9341,17'd10743,17'd17011,17'd9619,17'd10742,17'd16319,17'd20044,17'd27743,17'd33420,17'd46913,17'd46914,17'd46915,17'd31141,17'd30984,17'd15808,17'd29342,17'd41796,17'd15688,17'd29226,17'd46916,17'd46814,17'd46815,17'd46816,17'd46817,17'd46818,17'd46158,17'd46276,17'd46158,17'd36643,17'd46917,17'd46918,17'd46919,17'd46920,17'd46733,17'd46921,17'd46922,17'd46923,17'd45559,17'd46924,17'd35261,17'd46925,17'd46926,17'd46927,17'd45974,17'd40805,17'd46928,17'd33451,17'd46929,17'd46930,17'd36249,17'd33916,17'd46314,17'd46831,17'd42581,17'd42581,17'd43824,17'd34082,17'd44347,17'd36240,17'd46931,17'd42581,17'd34591,17'd34590,17'd46932,17'd46933,17'd35679,17'd44689,17'd37637,17'd36246,17'd41716,17'd38133,17'd38133,17'd40034,17'd46934,17'd40034,17'd36246,17'd35971,17'd36669,17'd37096,17'd37362,17'd37363,17'd37230,17'd37096,17'd37096,17'd37495,17'd37096,17'd37368,17'd39568,17'd37634,17'd37092,17'd46935,17'd46936,17'd46937,17'd46938,17'd46939,17'd37636,17'd46940,17'd46652,17'd46941,17'd46942,17'd46943,17'd46944,17'd46945,17'd46946,17'd44224,17'd46947,17'd44936,17'd46752,17'd46948,17'd43844,17'd44227,17'd43693,17'd43016,17'd43424,17'd44106,17'd43018,17'd43017,17'd38156,17'd27512,17'd25568,17'd25568,17'd25029,17'd28851,17'd29241,17'd29974,17'd36009,17'd46949,17'd37659,17'd22333,17'd22679,17'd36987,17'd23731,17'd25032,17'd28717,17'd31055,17'd28594,17'd29535,17'd36127,17'd35151,17'd46838,17'd46950,17'd40961,17'd38025,17'd46429,17'd46951,17'd35854,17'd27885,17'd28373,17'd30279,17'd30735,17'd26902,17'd26782,17'd27371,17'd27640,17'd27515,17'd25949,17'd28594,17'd25177,17'd25030,17'd24090,17'd30275,17'd23566,17'd23387,17'd29828,17'd29974,17'd32514,17'd29530,17'd30431,17'd24898,17'd25568,17'd27766,17'd26902,17'd46431,17'd28726,17'd39437,17'd31503,17'd34105,17'd46547,17'd46556,17'd46952,17'd46953,17'd46952,17'd46954,17'd46843,17'd44474,17'd41996,17'd46955,17'd46956,17'd45479,17'd46957,17'd45155,17'd38025,17'd31503,17'd28727,17'd27259,17'd28720,17'd24744,17'd23387,17'd46958,17'd46959,17'd46960,17'd46961,17'd46852,17'd46853,17'd46854,17'd46962,17'd46963,17'd46964,17'd46856,17'd46965,17'd40065,17'd45492,17'd36543,17'd23570,17'd46966,17'd23387,17'd23387,17'd46115,17'd23391,17'd31030,17'd46859,17'd21704,17'd46967,17'd46862,17'd46968,17'd46969,17'd46970,17'd46971,17'd46972,17'd46867,17'd44126,17'd46973,17'd46974,17'd20237,17'd28181,17'd46975,17'd31088,17'd46783,17'd46976,17'd27198,17'd16847,17'd46977,17'd46978,17'd38190,17'd19222,17'd14301,17'd35609,17'd35609,17'd35194,17'd5160,17'd4687,17'd5000,17'd39468,17'd42462,17'd41612,17'd41458,17'd33991,17'd4836,17'd4524,17'd34157,17'd46979,17'd4996,17'd4841,17'd4686,17'd32552,17'd4839,17'd4188,17'd4356,17'd46013,17'd35602,17'd46980,17'd46981,17'd46982,17'd46583,17'd46983,17'd46983,17'd41894,17'd46984,17'd46985,17'd46986,17'd46987,17'd46988,17'd46989,17'd37299,17'd46879,17'd46697,17'd46990,17'd2880,17'd40257,17'd37817,17'd46475,17'd46991,17'd7511,17'd5351,17'd41625,17'd41002,17'd18629,17'd40716,17'd11048,17'd39948,17'd38202,17'd38203,17'd38072,17'd44387,17'd44387,17'd16492,17'd16492,17'd16492,17'd6094,17'd6416,17'd8186,17'd5958,17'd5958,17'd5940,17'd5630,17'd16256,17'd15233,17'd33847,17'd33847,17'd944,17'd196,17'd13809,17'd46355,17'd1966,17'd971
},
'{
17'd4243,17'd4891,17'd5201,17'd5197,17'd5052,17'd5201,17'd3904,17'd14743,17'd2594,17'd466,17'd17,17'd17,17'd17,17'd17,17'd652,17'd652,17'd27,17'd652,17'd289,17'd31,17'd982,17'd984,17'd811,17'd471,17'd13303,17'd2939,17'd1972,17'd1971,17'd1134,17'd19609,17'd826,17'd992,17'd35772,17'd46024,17'd2798,17'd36606,17'd46992,17'd32412,17'd17308,17'd44853,17'd24516,17'd25910,17'd46702,17'd25801,17'd30057,17'd28205,17'd17204,17'd19754,17'd17320,17'd17448,17'd16034,17'd17207,17'd19007,17'd28667,17'd13211,17'd13093,17'd13094,17'd14471,17'd22630,17'd12361,17'd13093,17'd11626,17'd11914,17'd46993,17'd46994,17'd46995,17'd46996,17'd46997,17'd15140,17'd46998,17'd13844,17'd13844,17'd13470,17'd13470,17'd9301,17'd9007,17'd4611,17'd4767,17'd4926,17'd6627,17'd5250,17'd8541,17'd8691,17'd6779,17'd46999,17'd46896,17'd46897,17'd43073,17'd47000,17'd46800,17'd43207,17'd47001,17'd46495,17'd46711,17'd46801,17'd46902,17'd30210,17'd47002,17'd47003,17'd47004,17'd47005,17'd46805,17'd46716,17'd45928,17'd47006,17'd46910,17'd47007,17'd11968,17'd17240,17'd23343,17'd12723,17'd15297,17'd46380,17'd33725,17'd27006,17'd27006,17'd16561,17'd10332,17'd42674,17'd35799,17'd47008,17'd47009,17'd30076,17'd24537,17'd24856,17'd26371,17'd35513,17'd27122,17'd26149,17'd28231,17'd20608,17'd16442,17'd16326,17'd19158,17'd18917,17'd18198,17'd23515,17'd26370,17'd28943,17'd47010,17'd29329,17'd29329,17'd47011,17'd46912,17'd46912,17'd29778,17'd26493,17'd23170,17'd23169,17'd18326,17'd11400,17'd26152,17'd10024,17'd9741,17'd10743,17'd10857,17'd10743,17'd17011,17'd9619,17'd17011,17'd16319,17'd20044,17'd27864,17'd41346,17'd46913,17'd47012,17'd46915,17'd32940,17'd47013,17'd15808,17'd32590,17'd27002,17'd17839,17'd28578,17'd47014,17'd47015,17'd47016,17'd47017,17'd47018,17'd39986,17'd46158,17'd46160,17'd46158,17'd36643,17'd46917,17'd47019,17'd36364,17'd47020,17'd47021,17'd47022,17'd47023,17'd47024,17'd47025,17'd47026,17'd35261,17'd47027,17'd47028,17'd39411,17'd40805,17'd40501,17'd47029,17'd47030,17'd46531,17'd47031,17'd42865,17'd40502,17'd47032,17'd34732,17'd44578,17'd47033,17'd47033,17'd47034,17'd33452,17'd33452,17'd47035,17'd44465,17'd44465,17'd34075,17'd36388,17'd36522,17'd35835,17'd33620,17'd35273,17'd36965,17'd33620,17'd46934,17'd46934,17'd40034,17'd37370,17'd36246,17'd36384,17'd36669,17'd37096,17'd37230,17'd37231,17'd37095,17'd37095,17'd37095,17'd37230,17'd37095,17'd37096,17'd37366,17'd44922,17'd39412,17'd37362,17'd37762,17'd47036,17'd47037,17'd46938,17'd45361,17'd37364,17'd47038,17'd47039,17'd47040,17'd47041,17'd47042,17'd47043,17'd47044,17'd44588,17'd44224,17'd44472,17'd44828,17'd44592,17'd47045,17'd43559,17'd44935,17'd46547,17'd46425,17'd42599,17'd45749,17'd43156,17'd43155,17'd29825,17'd27512,17'd25568,17'd25178,17'd24897,17'd24742,17'd29099,17'd30277,17'd31343,17'd31657,17'd30427,17'd22680,17'd36426,17'd29686,17'd29534,17'd25030,17'd28717,17'd31055,17'd27766,17'd32006,17'd35707,17'd35567,17'd47046,17'd41416,17'd34275,17'd36264,17'd45748,17'd46951,17'd36541,17'd32832,17'd28373,17'd33952,17'd30735,17'd26902,17'd26782,17'd43290,17'd27883,17'd26903,17'd25949,17'd28594,17'd25177,17'd25030,17'd24090,17'd23732,17'd34137,17'd29376,17'd23923,17'd30579,17'd47047,17'd23733,17'd30126,17'd28254,17'd25709,17'd26174,17'd28486,17'd34767,17'd28979,17'd39437,17'd31354,17'd34104,17'd43834,17'd46661,17'd47048,17'd47049,17'd47050,17'd47051,17'd47052,17'd43545,17'd46846,17'd47053,17'd47054,17'd46762,17'd47055,17'd47056,17'd38025,17'd31503,17'd28979,17'd27515,17'd28600,17'd24416,17'd23388,17'd31348,17'd46330,17'd47057,17'd47058,17'd46767,17'd47059,17'd47060,17'd47061,17'd47062,17'd47063,17'd40687,17'd25183,17'd47064,17'd47065,17'd36543,17'd23570,17'd46442,17'd23387,17'd36152,17'd32030,17'd44944,17'd31192,17'd47066,17'd47067,17'd47068,17'd47069,17'd47070,17'd47071,17'd47072,17'd47073,17'd47074,17'd46867,17'd44006,17'd47075,17'd47076,17'd20524,17'd47077,17'd46975,17'd25225,17'd46783,17'd37027,17'd13925,17'd16847,17'd46977,17'd47078,17'd47079,17'd26585,17'd12760,17'd35609,17'd15990,17'd25084,17'd5160,17'd4687,17'd5000,17'd33691,17'd4358,17'd33533,17'd44009,17'd41891,17'd5000,17'd4999,17'd33991,17'd46979,17'd5153,17'd4841,17'd4686,17'd4687,17'd4683,17'd4991,17'd4356,17'd40547,17'd45394,17'd46980,17'd46981,17'd32871,17'd46583,17'd46873,17'd46231,17'd33688,17'd42036,17'd47080,17'd46986,17'd47081,17'd47082,17'd47083,17'd37568,17'd46879,17'd3365,17'd47084,17'd45066,17'd39480,17'd46881,17'd38855,17'd47085,17'd7511,17'd5351,17'd45656,17'd46136,17'd47086,17'd10790,17'd39181,17'd39483,17'd38202,17'd38203,17'd38203,17'd38581,17'd44387,17'd16492,17'd16492,17'd16492,17'd16492,17'd6258,17'd8186,17'd5958,17'd5958,17'd5940,17'd5630,17'd16382,17'd14586,17'd28428,17'd33847,17'd943,17'd417,17'd13573,17'd422,17'd1537,17'd1685
},
'{
17'd4892,17'd4891,17'd5201,17'd5645,17'd6263,17'd5202,17'd3904,17'd14743,17'd4247,17'd466,17'd17,17'd17,17'd289,17'd289,17'd652,17'd652,17'd980,17'd652,17'd289,17'd31,17'd982,17'd983,17'd984,17'd471,17'd13303,17'd2939,17'd1972,17'd1839,17'd47087,17'd46793,17'd16967,17'd17553,17'd35772,17'd46024,17'd2798,17'd36606,17'd46992,17'd32412,17'd17308,17'd16153,17'd47088,17'd25910,17'd46702,17'd24518,17'd45406,17'd18884,17'd11362,17'd11915,17'd17207,17'd16034,17'd46889,17'd20425,17'd18774,17'd29048,17'd13211,17'd13599,17'd14621,17'd14471,17'd22630,17'd13969,17'd12679,17'd24345,17'd11764,17'd47089,17'd47090,17'd47091,17'd47092,17'd47093,17'd15011,17'd15010,17'd13721,17'd13721,17'd13470,17'd13470,17'd12958,17'd9007,17'd4611,17'd4767,17'd4926,17'd6627,17'd5087,17'd8690,17'd8691,17'd6779,17'd47094,17'd40581,17'd6157,17'd6159,17'd47000,17'd46898,17'd46899,17'd46900,17'd46901,17'd46711,17'd46801,17'd47095,17'd47096,17'd8555,17'd47097,17'd47098,17'd47099,17'd47100,17'd47101,17'd47102,17'd47103,17'd47104,17'd47105,17'd17238,17'd13258,17'd8579,17'd19535,17'd8566,17'd13370,17'd10332,17'd27490,17'd27490,17'd17718,17'd13522,17'd22820,17'd11398,17'd23167,17'd24208,17'd26036,17'd24537,17'd27483,17'd26493,17'd35513,17'd27122,17'd35513,17'd47106,17'd20608,17'd16442,17'd16326,17'd13762,17'd12996,17'd18198,17'd23515,17'd29778,17'd29066,17'd47010,17'd29329,17'd29329,17'd47107,17'd30830,17'd30830,17'd30218,17'd29065,17'd24992,17'd23167,17'd23337,17'd12584,17'd10329,17'd10024,17'd9741,17'd10743,17'd10857,17'd9341,17'd17011,17'd25673,17'd16319,17'd10742,17'd9740,17'd29338,17'd41511,17'd46913,17'd31959,17'd46507,17'd47108,17'd47109,17'd47110,17'd10735,17'd10164,17'd12116,17'd15298,17'd47111,17'd47112,17'd47016,17'd47113,17'd47018,17'd46159,17'd47114,17'd46160,17'd46158,17'd36497,17'd47115,17'd47019,17'd47116,17'd37214,17'd47117,17'd47118,17'd47119,17'd47120,17'd47121,17'd47122,17'd47123,17'd44463,17'd41715,17'd47124,17'd38952,17'd47125,17'd47126,17'd47127,17'd47128,17'd38005,17'd47129,17'd47130,17'd35957,17'd34730,17'd34586,17'd34586,17'd34586,17'd35830,17'd47131,17'd36239,17'd33452,17'd42581,17'd35678,17'd36969,17'd37101,17'd35407,17'd33620,17'd33620,17'd35964,17'd47132,17'd34076,17'd38787,17'd37101,17'd33620,17'd36245,17'd36813,17'd37229,17'd46935,17'd37094,17'd37093,17'd37096,17'd37095,17'd37230,17'd37231,17'd37364,17'd38520,17'd37092,17'd37495,17'd38260,17'd39260,17'd47133,17'd47134,17'd46936,17'd43411,17'd47135,17'd47136,17'd37364,17'd47137,17'd44467,17'd47138,17'd47139,17'd47140,17'd47141,17'd47142,17'd43691,17'd44224,17'd44587,17'd38971,17'd46093,17'd41416,17'd43426,17'd42436,17'd43021,17'd42599,17'd43288,17'd33156,17'd44230,17'd43285,17'd39591,17'd25177,17'd25320,17'd25180,17'd24897,17'd34467,17'd23387,17'd22679,17'd31343,17'd37510,17'd22332,17'd39131,17'd39278,17'd29099,17'd29688,17'd25180,17'd28717,17'd28598,17'd25833,17'd32343,17'd41429,17'd36401,17'd47143,17'd43701,17'd34105,17'd35291,17'd38665,17'd39275,17'd32506,17'd28134,17'd28134,17'd33952,17'd31035,17'd26782,17'd26782,17'd33499,17'd33815,17'd26903,17'd28602,17'd27765,17'd25568,17'd24898,17'd24090,17'd24086,17'd34137,17'd29099,17'd35865,17'd29530,17'd47144,17'd29527,17'd34276,17'd25568,17'd25567,17'd25833,17'd31035,17'd47145,17'd28980,17'd31354,17'd35570,17'd37658,17'd45610,17'd46661,17'd47146,17'd47147,17'd47148,17'd47051,17'd40364,17'd42881,17'd46955,17'd43830,17'd47054,17'd46762,17'd47055,17'd47056,17'd33791,17'd39437,17'd26781,17'd27514,17'd28484,17'd23916,17'd23388,17'd31031,17'd47149,17'd47150,17'd47058,17'd47151,17'd47152,17'd47153,17'd47154,17'd47155,17'd47156,17'd47157,17'd24905,17'd47158,17'd47159,17'd36543,17'd23570,17'd31836,17'd23923,17'd29374,17'd31836,17'd32190,17'd21850,17'd47160,17'd47161,17'd47162,17'd47163,17'd47070,17'd47164,17'd47165,17'd47166,17'd40973,17'd47167,17'd47168,17'd47169,17'd22548,17'd47170,17'd22411,17'd47171,17'd47172,17'd46783,17'd46976,17'd16123,17'd16847,17'd46978,17'd47173,17'd26710,17'd19088,17'd13800,17'd15990,17'd15990,17'd6392,17'd5160,17'd4845,17'd5001,17'd4515,17'd4018,17'd33533,17'd33840,17'd41891,17'd5000,17'd4525,17'd4188,17'd33532,17'd47174,17'd4842,17'd5005,17'd4845,17'd4840,17'd38442,17'd4356,17'd46228,17'd35602,17'd34327,17'd46981,17'd47175,17'd46230,17'd46873,17'd46231,17'd41464,17'd41469,17'd47176,17'd47177,17'd47081,17'd47082,17'd47178,17'd37299,17'd46788,17'd47179,17'd35056,17'd22095,17'd47180,17'd37817,17'd47181,17'd4050,17'd5023,17'd5351,17'd10071,17'd45185,17'd47086,17'd10790,17'd11048,17'd39948,17'd38202,17'd38203,17'd38203,17'd38581,17'd44387,17'd16492,17'd16492,17'd16492,17'd6258,17'd8186,17'd8186,17'd5958,17'd5958,17'd5940,17'd5630,17'd16382,17'd15233,17'd33847,17'd2560,17'd943,17'd417,17'd194,17'd1381,17'd972,17'd971
},
'{
17'd4244,17'd4891,17'd5201,17'd4735,17'd4888,17'd4087,17'd3904,17'd47182,17'd4247,17'd466,17'd17,17'd17,17'd289,17'd653,17'd652,17'd28,17'd980,17'd652,17'd289,17'd31,17'd982,17'd983,17'd984,17'd471,17'd13303,17'd1968,17'd1972,17'd1971,17'd1134,17'd19609,17'd992,17'd17553,17'd35772,17'd1561,17'd2798,17'd36606,17'd46992,17'd20018,17'd17308,17'd16153,17'd47183,17'd47184,17'd24683,17'd25801,17'd45406,17'd18884,17'd17941,17'd16766,17'd16519,17'd15902,17'd16034,17'd20425,17'd18774,17'd16765,17'd13211,17'd13093,17'd13094,17'd13969,17'd13969,17'd14764,17'd12527,17'd12813,17'd11764,17'd22463,17'd22462,17'd47185,17'd47185,17'd47093,17'd47186,17'd15010,17'd22631,17'd13721,17'd13721,17'd13470,17'd12959,17'd9301,17'd4611,17'd4767,17'd4767,17'd4926,17'd6627,17'd5251,17'd8690,17'd7099,17'd47187,17'd40731,17'd47188,17'd6159,17'd46253,17'd46800,17'd43207,17'd47001,17'd46495,17'd46711,17'd47189,17'd33561,17'd47096,17'd47190,17'd47191,17'd47098,17'd47192,17'd47193,17'd47100,17'd47194,17'd47195,17'd47104,17'd47196,17'd47197,17'd17850,17'd10028,17'd17481,17'd8879,17'd10026,17'd27744,17'd27490,17'd27490,17'd17718,17'd13522,17'd22820,17'd43622,17'd29783,17'd46383,17'd30076,17'd24537,17'd27483,17'd26493,17'd35513,17'd27122,17'd35513,17'd32127,17'd20608,17'd18443,17'd18444,17'd16326,17'd18917,17'd18559,17'd23515,17'd26872,17'd29066,17'd47010,17'd30527,17'd30527,17'd47010,17'd47107,17'd30831,17'd29923,17'd29327,17'd24538,17'd24858,17'd17478,17'd11398,17'd11526,17'd16796,17'd9741,17'd10742,17'd10857,17'd9341,17'd17011,17'd9619,17'd16319,17'd27003,17'd10856,17'd28819,17'd23510,17'd35655,17'd31959,17'd46724,17'd47198,17'd33411,17'd47199,17'd10852,17'd10741,17'd11809,17'd24366,17'd47111,17'd47200,17'd35527,17'd47201,17'd47202,17'd47203,17'd31972,17'd46158,17'd47114,17'd36497,17'd47204,17'd47205,17'd47206,17'd47207,17'd35533,17'd46921,17'd47208,17'd47209,17'd47210,17'd46393,17'd47211,17'd47211,17'd46518,17'd47212,17'd34728,17'd47213,17'd47030,17'd47214,17'd47215,17'd47216,17'd47217,17'd47218,17'd34856,17'd47219,17'd34992,17'd34586,17'd47219,17'd47220,17'd47221,17'd33452,17'd43136,17'd44347,17'd34994,17'd35678,17'd33916,17'd33916,17'd40199,17'd42424,17'd47222,17'd47222,17'd33916,17'd38787,17'd35834,17'd38645,17'd39116,17'd37229,17'd38646,17'd37093,17'd37093,17'd37093,17'd37095,17'd37231,17'd37363,17'd37231,17'd38520,17'd37635,17'd36661,17'd37096,17'd46194,17'd47223,17'd47224,17'd47225,17'd38520,17'd41567,17'd47226,17'd47227,17'd37636,17'd47228,17'd47229,17'd47230,17'd47231,17'd47232,17'd47233,17'd47234,17'd39582,17'd46947,17'd45370,17'd45872,17'd43692,17'd44103,17'd42436,17'd43021,17'd46200,17'd44590,17'd43288,17'd33156,17'd44230,17'd46426,17'd28484,17'd25709,17'd25320,17'd25030,17'd24745,17'd23917,17'd30128,17'd23038,17'd35296,17'd30426,17'd22680,17'd32830,17'd38976,17'd23920,17'd28977,17'd25320,17'd31520,17'd27513,17'd25707,17'd33477,17'd41274,17'd40823,17'd47235,17'd43434,17'd34105,17'd35425,17'd40365,17'd38805,17'd39437,17'd27885,17'd28134,17'd30279,17'd28486,17'd27371,17'd26782,17'd33499,17'd33815,17'd27515,17'd28602,17'd27765,17'd25568,17'd24897,17'd24090,17'd23731,17'd34137,17'd23918,17'd31502,17'd23566,17'd47236,17'd34883,17'd30432,17'd31366,17'd27513,17'd27259,17'd29245,17'd44703,17'd29246,17'd32356,17'd35707,17'd43696,17'd46432,17'd46756,17'd47237,17'd47234,17'd47238,17'd47148,17'd46954,17'd43153,17'd46955,17'd47239,17'd46956,17'd45879,17'd47240,17'd47241,17'd36690,17'd31353,17'd26782,17'd25949,17'd28484,17'd23916,17'd23569,17'd31193,17'd47149,17'd47150,17'd47242,17'd47243,17'd47244,17'd47245,17'd47246,17'd47247,17'd47156,17'd47157,17'd47248,17'd47158,17'd47065,17'd36543,17'd23570,17'd34277,17'd30128,17'd23215,17'd32679,17'd23926,17'd21850,17'd35428,17'd47249,17'd47250,17'd21703,17'd46968,17'd47251,17'd47252,17'd47253,17'd47254,17'd47255,17'd43724,17'd47256,17'd47257,17'd21134,17'd22411,17'd46975,17'd47258,17'd46582,17'd37027,17'd12622,17'd16847,17'd38190,17'd47259,17'd47260,17'd26585,17'd14049,17'd15990,17'd44613,17'd6391,17'd5160,17'd4845,17'd5001,17'd34157,17'd4358,17'd39468,17'd33840,17'd33841,17'd5156,17'd5155,17'd38442,17'd33532,17'd5152,17'd5005,17'd5005,17'd5002,17'd4841,17'd38442,17'd4356,17'd46228,17'd45394,17'd34327,17'd46981,17'd47175,17'd46230,17'd46873,17'd47261,17'd44134,17'd47262,17'd47263,17'd47177,17'd47264,17'd47265,17'd46988,17'd47266,17'd3364,17'd47267,17'd35056,17'd21940,17'd47268,17'd46881,17'd2892,17'd47269,17'd5023,17'd5351,17'd10071,17'd45185,17'd47086,17'd10790,17'd39181,17'd39483,17'd38202,17'd38580,17'd38203,17'd38581,17'd44387,17'd37959,17'd16492,17'd16492,17'd6258,17'd8186,17'd8186,17'd5958,17'd4882,17'd5940,17'd5630,17'd16382,17'd35060,17'd34000,17'd1950,17'd942,17'd417,17'd415,17'd424,17'd972,17'd972
},
'{
17'd47270,17'd29756,17'd4087,17'd4426,17'd27097,17'd4892,17'd2784,17'd14188,17'd2594,17'd1127,17'd17,17'd17,17'd3905,17'd1128,17'd980,17'd1278,17'd652,17'd652,17'd289,17'd31,17'd2940,17'd45516,17'd46358,17'd13303,17'd2428,17'd2261,17'd2121,17'd1282,17'd19499,17'd19609,17'd992,17'd18150,17'd2610,17'd3439,17'd2797,17'd2801,17'd46887,17'd47271,17'd14329,17'd16153,17'd24516,17'd25257,17'd47272,17'd46359,17'd47273,17'd28667,17'd19006,17'd19007,17'd16519,17'd24348,17'd47274,17'd16986,17'd19006,17'd12361,17'd13211,17'd17096,17'd12530,17'd13840,17'd47275,17'd19890,17'd13092,17'd13093,17'd12531,17'd16410,17'd47186,17'd47276,17'd5407,17'd47277,17'd5407,17'd47278,17'd22631,17'd13843,17'd13721,17'd13470,17'd12959,17'd12958,17'd8538,17'd7750,17'd10430,17'd4927,17'd5252,17'd8689,17'd8692,17'd7259,17'd39647,17'd47279,17'd44155,17'd42503,17'd47000,17'd47280,17'd45668,17'd41334,17'd39202,17'd47281,17'd47282,17'd47283,17'd47284,17'd47190,17'd47285,17'd47286,17'd28333,17'd47287,17'd47005,17'd47288,17'd47195,17'd47289,17'd47290,17'd47291,17'd9350,17'd8580,17'd24713,17'd47292,17'd47293,17'd34042,17'd27006,17'd17479,17'd17847,17'd26369,17'd17966,17'd43622,17'd24540,17'd46383,17'd30076,17'd24537,17'd25527,17'd24857,17'd32127,17'd27122,17'd47294,17'd32127,17'd22992,17'd19158,17'd11964,17'd16326,17'd18917,17'd18198,17'd19407,17'd23511,17'd28460,17'd29067,17'd31764,17'd47295,17'd47296,17'd29329,17'd47010,17'd30831,17'd29923,17'd27004,17'd23170,17'd24858,17'd11397,17'd28352,17'd10330,17'd10856,17'd10742,17'd10743,17'd9340,17'd9341,17'd9741,17'd9740,17'd46267,17'd46267,17'd18916,17'd41194,17'd35243,17'd47012,17'd47297,17'd46915,17'd32940,17'd29492,17'd29342,17'd10023,17'd10174,17'd17347,17'd47298,17'd47299,17'd47300,17'd47301,17'd47302,17'd47303,17'd47304,17'd47305,17'd47114,17'd47306,17'd47019,17'd47307,17'd47308,17'd47309,17'd47310,17'd47311,17'd47312,17'd47313,17'd47314,17'd47315,17'd47316,17'd47317,17'd47318,17'd47319,17'd46396,17'd47320,17'd47321,17'd46928,17'd47322,17'd47323,17'd47324,17'd47130,17'd47219,17'd33920,17'd33920,17'd33915,17'd40502,17'd47033,17'd36249,17'd47221,17'd38644,17'd42581,17'd46931,17'd44465,17'd46931,17'd36378,17'd36378,17'd42581,17'd42135,17'd36969,17'd38787,17'd36247,17'd36384,17'd37368,17'd37096,17'd37230,17'd37230,17'd37230,17'd37096,17'd37096,17'd37096,17'd37096,17'd37095,17'd37095,17'd37495,17'd37366,17'd37093,17'd46935,17'd47325,17'd47325,17'd37494,17'd37362,17'd38262,17'd35972,17'd47326,17'd45976,17'd37366,17'd47327,17'd47328,17'd47329,17'd46943,17'd47330,17'd47331,17'd47332,17'd39582,17'd44472,17'd45264,17'd47333,17'd41416,17'd44935,17'd44700,17'd43021,17'd43548,17'd47334,17'd43979,17'd44106,17'd44359,17'd45036,17'd28130,17'd28597,17'd27512,17'd25032,17'd35159,17'd31502,17'd23218,17'd23038,17'd30427,17'd22333,17'd22330,17'd32830,17'd23387,17'd24249,17'd29533,17'd27512,17'd32669,17'd26174,17'd28724,17'd42301,17'd45747,17'd47235,17'd44361,17'd41108,17'd35707,17'd35853,17'd37904,17'd39741,17'd47335,17'd47336,17'd28370,17'd26277,17'd31035,17'd26782,17'd43290,17'd43290,17'd27640,17'd25833,17'd25566,17'd28369,17'd25178,17'd28718,17'd24743,17'd28722,17'd30879,17'd31033,17'd23731,17'd29378,17'd47337,17'd33802,17'd27882,17'd38671,17'd27639,17'd28853,17'd35011,17'd28726,17'd29246,17'd31354,17'd41731,17'd39436,17'd46660,17'd46759,17'd47146,17'd47338,17'd47339,17'd47340,17'd47341,17'd47342,17'd47343,17'd47344,17'd46847,17'd47345,17'd45872,17'd44700,17'd36264,17'd27642,17'd27259,17'd25708,17'd28369,17'd34467,17'd22501,17'd47346,17'd47347,17'd47348,17'd46209,17'd47349,17'd47350,17'd47351,17'd47352,17'd47353,17'd47354,17'd37269,17'd47355,17'd47356,17'd47357,17'd46442,17'd23217,17'd23218,17'd22502,17'd45874,17'd32190,17'd31834,17'd47358,17'd47359,17'd47360,17'd47361,17'd47362,17'd47363,17'd47364,17'd41127,17'd41438,17'd47365,17'd47366,17'd47367,17'd47368,17'd22050,17'd21134,17'd29156,17'd27304,17'd46126,17'd47369,17'd36443,17'd12622,17'd36028,17'd36030,17'd47370,17'd47259,17'd47371,17'd13678,17'd30179,17'd30332,17'd6220,17'd5335,17'd5002,17'd4529,17'd34157,17'd4833,17'd33839,17'd33840,17'd4999,17'd4683,17'd42910,17'd5145,17'd33532,17'd5152,17'd4842,17'd5004,17'd30637,17'd4841,17'd5144,17'd41455,17'd46013,17'd47372,17'd4825,17'd5601,17'd3827,17'd33688,17'd45511,17'd33529,17'd46232,17'd46875,17'd47373,17'd47374,17'd47375,17'd47177,17'd47376,17'd38063,17'd47377,17'd37038,17'd47378,17'd41310,17'd47379,17'd47380,17'd47381,17'd47382,17'd9661,17'd45656,17'd10071,17'd45185,17'd47086,17'd10790,17'd39032,17'd38458,17'd38202,17'd38860,17'd38860,17'd38581,17'd44387,17'd16492,17'd16492,17'd6258,17'd6258,17'd8186,17'd8186,17'd5958,17'd4882,17'd4882,17'd5940,17'd16256,17'd34000,17'd33847,17'd2560,17'd943,17'd195,17'd2920,17'd32250,17'd973,17'd270
},
'{
17'd30047,17'd5200,17'd4087,17'd4426,17'd27097,17'd25384,17'd2784,17'd14070,17'd1831,17'd1127,17'd17,17'd3905,17'd20404,17'd1128,17'd980,17'd980,17'd652,17'd29,17'd809,17'd31,17'd2940,17'd45516,17'd46358,17'd13303,17'd2428,17'd2261,17'd1971,17'd1837,17'd990,17'd19609,17'd992,17'd18150,17'd2610,17'd3439,17'd2797,17'd3447,17'd46887,17'd47271,17'd14329,17'd16153,17'd45188,17'd47383,17'd47384,17'd45519,17'd47273,17'd28667,17'd20148,17'd19007,17'd17320,17'd15524,17'd18414,17'd19007,17'd12681,17'd12362,17'd13211,17'd23154,17'd11913,17'd13969,17'd14891,17'd19890,17'd13598,17'd17096,17'd17317,17'd16164,17'd47186,17'd47385,17'd5407,17'd47277,17'd47276,17'd47386,17'd16032,17'd15007,17'd22631,17'd13721,17'd12959,17'd12959,17'd8538,17'd7750,17'd10430,17'd5255,17'd5252,17'd8689,17'd8692,17'd7259,17'd39647,17'd47279,17'd44155,17'd42800,17'd47000,17'd47387,17'd45668,17'd47388,17'd39061,17'd47281,17'd47282,17'd47389,17'd47284,17'd30362,17'd47390,17'd47391,17'd47392,17'd47287,17'd47393,17'd47394,17'd47395,17'd47396,17'd47397,17'd47398,17'd47399,17'd8580,17'd24713,17'd47400,17'd34383,17'd34042,17'd47401,17'd17479,17'd42674,17'd47402,17'd17966,17'd43622,17'd24540,17'd27860,17'd30076,17'd24856,17'd27347,17'd26493,17'd35513,17'd26871,17'd27622,17'd32127,17'd21361,17'd16326,17'd11964,17'd18444,17'd18917,17'd17722,17'd14807,17'd23855,17'd27857,17'd28686,17'd47403,17'd47404,17'd30527,17'd29329,17'd47010,17'd47010,17'd30831,17'd29778,17'd26756,17'd21362,17'd18327,17'd21206,17'd10330,17'd16796,17'd9885,17'd10743,17'd9620,17'd9620,17'd9741,17'd10856,17'd46267,17'd47405,17'd17012,17'd20044,17'd35243,17'd47012,17'd32141,17'd46914,17'd32449,17'd40746,17'd16198,17'd10023,17'd9194,17'd47406,17'd47407,17'd47408,17'd37618,17'd47301,17'd47016,17'd47409,17'd47203,17'd40147,17'd47410,17'd47306,17'd47019,17'd47411,17'd47412,17'd47413,17'd43488,17'd47414,17'd47415,17'd47209,17'd47416,17'd47417,17'd47418,17'd47419,17'd47420,17'd47421,17'd47418,17'd47422,17'd47423,17'd47424,17'd47425,17'd33616,17'd47324,17'd47130,17'd34992,17'd34856,17'd46313,17'd40033,17'd33618,17'd36099,17'd40502,17'd47033,17'd36249,17'd47035,17'd47035,17'd47035,17'd38644,17'd46931,17'd36378,17'd33916,17'd33769,17'd35407,17'd36246,17'd36385,17'd37634,17'd37366,17'd37096,17'd37096,17'd37495,17'd37366,17'd37495,17'd37495,17'd37096,17'd37096,17'd37495,17'd37495,17'd37366,17'd37495,17'd37093,17'd47426,17'd47427,17'd47428,17'd47325,17'd44922,17'd38263,17'd37634,17'd46935,17'd37093,17'd47429,17'd47430,17'd47431,17'd47432,17'd47433,17'd47434,17'd47435,17'd47436,17'd47148,17'd45480,17'd47437,17'd47045,17'd43700,17'd43693,17'd46200,17'd46200,17'd47334,17'd46753,17'd43018,17'd43156,17'd44359,17'd47438,17'd28130,17'd33000,17'd27512,17'd25032,17'd30431,17'd35865,17'd23389,17'd23038,17'd23573,17'd33311,17'd39131,17'd39278,17'd34137,17'd29688,17'd27637,17'd46549,17'd30734,17'd26174,17'd27260,17'd42298,17'd46658,17'd47439,17'd40217,17'd38974,17'd35152,17'd36125,17'd38973,17'd42890,17'd47335,17'd47440,17'd26276,17'd26652,17'd28727,17'd26782,17'd43290,17'd27371,17'd27640,17'd25833,17'd28723,17'd28369,17'd25178,17'd24417,17'd24743,17'd29100,17'd23917,17'd24415,17'd34467,17'd23563,17'd47441,17'd33318,17'd28598,17'd41115,17'd28009,17'd27027,17'd36542,17'd28486,17'd29379,17'd32356,17'd34275,17'd46094,17'd46755,17'd46842,17'd47237,17'd47442,17'd47443,17'd47341,17'd47444,17'd47445,17'd47343,17'd47446,17'd46666,17'd47345,17'd45872,17'd46200,17'd36127,17'd29379,17'd27259,17'd27766,17'd27882,17'd24252,17'd22501,17'd31347,17'd47447,17'd47448,17'd47449,17'd47450,17'd47350,17'd47351,17'd47451,17'd47452,17'd47453,17'd45625,17'd46219,17'd47454,17'd47455,17'd47456,17'd23217,17'd23218,17'd22327,17'd47457,17'd39441,17'd23394,17'd21850,17'd43557,17'd47360,17'd47458,17'd47459,17'd47460,17'd47461,17'd41127,17'd47462,17'd47463,17'd44723,17'd47464,17'd47465,17'd24458,17'd47466,17'd29156,17'd47467,17'd22588,17'd47468,17'd47469,17'd12622,17'd28059,17'd36444,17'd37429,17'd47259,17'd24803,17'd14049,17'd30179,17'd30332,17'd6219,17'd28185,17'd5002,17'd34656,17'd33992,17'd33991,17'd33691,17'd47470,17'd4999,17'd4683,17'd42910,17'd6067,17'd47471,17'd5152,17'd4842,17'd5004,17'd30637,17'd4686,17'd5144,17'd41612,17'd4828,17'd47372,17'd34496,17'd47472,17'd4179,17'd41464,17'd46690,17'd41760,17'd3675,17'd47473,17'd47474,17'd47374,17'd47375,17'd47475,17'd47476,17'd47477,17'd47478,17'd37038,17'd47479,17'd20706,17'd47480,17'd47481,17'd47482,17'd47483,17'd9661,17'd45656,17'd10071,17'd45185,17'd43462,17'd10790,17'd39181,17'd39483,17'd38859,17'd38860,17'd38860,17'd38581,17'd44387,17'd16492,17'd16492,17'd6258,17'd6258,17'd8186,17'd8186,17'd5958,17'd4882,17'd4882,17'd4882,17'd9123,17'd35060,17'd47484,17'd33847,17'd196,17'd778,17'd951,17'd1966,17'd1963,17'd269
},
'{
17'd5202,17'd5201,17'd4087,17'd4891,17'd27441,17'd25384,17'd2784,17'd27714,17'd2594,17'd1127,17'd17,17'd3905,17'd20404,17'd1128,17'd980,17'd980,17'd652,17'd652,17'd289,17'd30,17'd3256,17'd45516,17'd46358,17'd13303,17'd2428,17'd2261,17'd1971,17'd1282,17'd19499,17'd46885,17'd17079,17'd18150,17'd2610,17'd3439,17'd2797,17'd2801,17'd47485,17'd47486,17'd17088,17'd47487,17'd24516,17'd47488,17'd47489,17'd45519,17'd47273,17'd28667,17'd20148,17'd19007,17'd17320,17'd24348,17'd47490,17'd21649,17'd12532,17'd12362,17'd13211,17'd17096,17'd12361,17'd13840,17'd16286,17'd19890,17'd12954,17'd17096,17'd17317,17'd16289,17'd15139,17'd47491,17'd47385,17'd4603,17'd47492,17'd16031,17'd14625,17'd14475,17'd14100,17'd13468,17'd12959,17'd9575,17'd8538,17'd8538,17'd7750,17'd5255,17'd5253,17'd8689,17'd8692,17'd8070,17'd46709,17'd47279,17'd40733,17'd42800,17'd44864,17'd47280,17'd45668,17'd45669,17'd39202,17'd47281,17'd47282,17'd47389,17'd47493,17'd47494,17'd47495,17'd47496,17'd47497,17'd28091,17'd47192,17'd47498,17'd47499,17'd47500,17'd47501,17'd47502,17'd42809,17'd8251,17'd23343,17'd31759,17'd47503,17'd37470,17'd27006,17'd12585,17'd11526,17'd36482,17'd17966,17'd23166,17'd36348,17'd27985,17'd30076,17'd25927,17'd24537,17'd24030,17'd24992,17'd26372,17'd27122,17'd35513,17'd24706,17'd18327,17'd11964,17'd18444,17'd18917,17'd18197,17'd14807,17'd23855,17'd28104,17'd29645,17'd47295,17'd47403,17'd30527,17'd30527,17'd47296,17'd29329,17'd30071,17'd28343,17'd24859,17'd21363,17'd23513,17'd11808,17'd24996,17'd16796,17'd9885,17'd9885,17'd9742,17'd9742,17'd9885,17'd10856,17'd46267,17'd47405,17'd9472,17'd9611,17'd29795,17'd47504,17'd32141,17'd31957,17'd47505,17'd34709,17'd16198,17'd10741,17'd9348,17'd37604,17'd28840,17'd47506,17'd47507,17'd47300,17'd47508,17'd39519,17'd40893,17'd47509,17'd47510,17'd47511,17'd47205,17'd47512,17'd47412,17'd47513,17'd47514,17'd47515,17'd47516,17'd47517,17'd46515,17'd47518,17'd47519,17'd39411,17'd47213,17'd47520,17'd47521,17'd46412,17'd34073,17'd47029,17'd46928,17'd40661,17'd47522,17'd42865,17'd33765,17'd33765,17'd40033,17'd40033,17'd33618,17'd36099,17'd36099,17'd40502,17'd47033,17'd36249,17'd47221,17'd36523,17'd42581,17'd42135,17'd34994,17'd37235,17'd41716,17'd35972,17'd36669,17'd37634,17'd37367,17'd37367,17'd37367,17'd37634,17'd36669,17'd36670,17'd38391,17'd37634,17'd37366,17'd37366,17'd37366,17'd37366,17'd37495,17'd37096,17'd37094,17'd47426,17'd47134,17'd47427,17'd47428,17'd39262,17'd36965,17'd47523,17'd37362,17'd46315,17'd47524,17'd38960,17'd47525,17'd47526,17'd47527,17'd47528,17'd47529,17'd47530,17'd47531,17'd45157,17'd44592,17'd46658,17'd44103,17'd42741,17'd42886,17'd42886,17'd46753,17'd44934,17'd46095,17'd46095,17'd43978,17'd43978,17'd28130,17'd33484,17'd27637,17'd28368,17'd31033,17'd23923,17'd41273,17'd23038,17'd22856,17'd22500,17'd23740,17'd29828,17'd24087,17'd40964,17'd25029,17'd31520,17'd26062,17'd25833,17'd47334,17'd46658,17'd46948,17'd39129,17'd47532,17'd40958,17'd37658,17'd39274,17'd37904,17'd34275,17'd35152,17'd36127,17'd26276,17'd25697,17'd28979,17'd33963,17'd27371,17'd27259,17'd26903,17'd25833,17'd28723,17'd28369,17'd27637,17'd24744,17'd28601,17'd24090,17'd32659,17'd32659,17'd29688,17'd47533,17'd28367,17'd38282,17'd28594,17'd27639,17'd27883,17'd33163,17'd35426,17'd28727,17'd27642,17'd32506,17'd34451,17'd42436,17'd46839,17'd47050,17'd47443,17'd47534,17'd47444,17'd47535,17'd47536,17'd47537,17'd47344,17'd47538,17'd46847,17'd47539,17'd46752,17'd42886,17'd36127,17'd29379,17'd27640,17'd27766,17'd27882,17'd24743,17'd30277,17'd31347,17'd47540,17'd47541,17'd47542,17'd47543,17'd47544,17'd47545,17'd45993,17'd47452,17'd47453,17'd47546,17'd46219,17'd47547,17'd47455,17'd47456,17'd23216,17'd36986,17'd22326,17'd22325,17'd23926,17'd23394,17'd22013,17'd47548,17'd47360,17'd47069,17'd47549,17'd47550,17'd47551,17'd41127,17'd47552,17'd47553,17'd47554,17'd47555,17'd47556,17'd47557,17'd21605,17'd22411,17'd47467,17'd47558,17'd47468,17'd23633,17'd14301,17'd28059,17'd36444,17'd36310,17'd47259,17'd36028,17'd12160,17'd30179,17'd10514,17'd6219,17'd28185,17'd5329,17'd34656,17'd33991,17'd4833,17'd33839,17'd33840,17'd4999,17'd4683,17'd42910,17'd6067,17'd4997,17'd4995,17'd5005,17'd5004,17'd5004,17'd4686,17'd4838,17'd4016,17'd4828,17'd34654,17'd34154,17'd47559,17'd4179,17'd41302,17'd47560,17'd47561,17'd47562,17'd47563,17'd46986,17'd47375,17'd39619,17'd47564,17'd47476,17'd47565,17'd47478,17'd37163,17'd47566,17'd47567,17'd47568,17'd47569,17'd3556,17'd7023,17'd9661,17'd45656,17'd10071,17'd46354,17'd43462,17'd10790,17'd39482,17'd39483,17'd38859,17'd38860,17'd38860,17'd38072,17'd13420,17'd16492,17'd16492,17'd16492,17'd6258,17'd8186,17'd8186,17'd5958,17'd4882,17'd4882,17'd5940,17'd16256,17'd15233,17'd29440,17'd33847,17'd196,17'd600,17'd422,17'd205,17'd1963,17'd261
},
'{
17'd5201,17'd4735,17'd4087,17'd4891,17'd27590,17'd6420,17'd2784,17'd14070,17'd1831,17'd1127,17'd17,17'd3905,17'd1128,17'd1128,17'd27,17'd980,17'd652,17'd29,17'd809,17'd31,17'd2940,17'd45516,17'd46358,17'd13303,17'd2428,17'd2261,17'd1971,17'd1837,17'd989,17'd19609,17'd992,17'd18150,17'd2610,17'd34168,17'd2797,17'd3447,17'd46887,17'd47271,17'd14329,17'd16153,17'd45188,17'd47488,17'd47489,17'd47570,17'd47571,17'd28667,17'd20148,17'd27461,17'd17320,17'd15902,17'd22980,17'd21649,17'd12532,17'd12362,17'd13211,17'd23154,17'd11913,17'd13969,17'd14891,17'd19890,17'd13599,17'd29904,17'd23155,17'd16519,17'd15260,17'd47572,17'd47573,17'd47491,17'd47574,17'd16031,17'd16030,17'd14474,17'd14345,17'd14099,17'd13468,17'd9575,17'd8538,17'd8538,17'd7750,17'd5689,17'd5253,17'd5252,17'd6137,17'd7259,17'd39647,17'd47279,17'd40584,17'd44283,17'd47575,17'd47576,17'd47577,17'd45199,17'd39202,17'd47281,17'd47282,17'd47578,17'd47579,17'd47580,17'd47581,17'd47582,17'd47583,17'd47584,17'd47585,17'd47586,17'd47587,17'd47588,17'd47589,17'd47590,17'd25410,17'd8251,17'd8579,17'd24712,17'd47591,17'd47592,17'd27006,17'd31445,17'd34956,17'd17966,17'd37983,17'd23166,17'd36348,17'd29928,17'd30076,17'd24856,17'd24537,17'd24538,17'd26495,17'd26150,17'd26871,17'd47009,17'd14259,17'd18327,17'd13516,17'd13516,17'd12996,17'd18917,17'd16321,17'd12254,17'd28103,17'd29645,17'd31764,17'd47403,17'd47593,17'd47594,17'd47595,17'd30527,17'd35931,17'd28344,17'd27004,17'd22818,17'd22472,17'd11396,17'd28352,17'd26152,17'd10024,17'd9741,17'd9742,17'd9742,17'd9885,17'd9885,17'd9473,17'd27003,17'd18332,17'd47596,17'd34217,17'd47597,17'd47598,17'd47297,17'd47505,17'd34049,17'd21982,17'd10164,17'd9348,17'd8575,17'd47599,17'd47600,17'd47507,17'd47601,17'd47602,17'd47603,17'd47604,17'd36224,17'd47605,17'd47606,17'd47601,17'd47512,17'd47607,17'd47608,17'd47609,17'd47610,17'd47611,17'd47612,17'd47613,17'd47614,17'd42864,17'd47521,17'd46927,17'd47029,17'd39719,17'd43003,17'd47615,17'd33913,17'd47616,17'd47617,17'd40944,17'd45471,17'd33764,17'd47618,17'd47619,17'd33915,17'd33915,17'd40502,17'd47033,17'd45860,17'd36249,17'd47035,17'd38644,17'd42581,17'd34994,17'd33769,17'd35407,17'd36965,17'd36385,17'd38391,17'd38391,17'd38391,17'd36670,17'd36244,17'd36384,17'd36244,17'd36244,17'd36384,17'd36384,17'd36670,17'd36669,17'd37367,17'd37367,17'd37367,17'd37366,17'd37495,17'd37096,17'd37230,17'd37361,17'd47225,17'd46194,17'd44690,17'd39116,17'd37762,17'd37363,17'd47620,17'd47621,17'd47622,17'd47623,17'd47624,17'd47625,17'd47626,17'd40215,17'd46953,17'd47627,17'd47628,17'd44479,17'd43844,17'd42298,17'd43021,17'd46425,17'd46425,17'd44934,17'd44934,17'd47629,17'd47629,17'd37778,17'd37778,17'd27765,17'd28480,17'd27637,17'd28368,17'd23732,17'd29828,17'd41273,17'd22678,17'd22330,17'd22329,17'd32667,17'd23566,17'd38978,17'd38667,17'd28719,17'd28598,17'd27515,17'd35012,17'd45745,17'd47630,17'd44479,17'd46658,17'd47631,17'd43289,17'd41417,17'd47632,17'd36686,17'd34877,17'd35854,17'd32356,17'd47633,17'd26780,17'd28726,17'd35023,17'd27371,17'd26782,17'd27259,17'd25833,17'd28723,17'd27882,17'd25029,17'd24744,17'd34884,17'd24415,17'd29688,17'd30126,17'd34276,17'd47634,17'd28974,17'd44229,17'd26064,17'd26530,17'd27371,17'd30735,17'd39437,17'd29246,17'd30279,17'd36403,17'd34274,17'd43693,17'd47635,17'd47636,17'd47637,17'd47638,17'd47639,17'd47640,17'd47640,17'd45607,17'd47641,17'd47641,17'd46847,17'd45879,17'd44102,17'd42886,17'd39437,17'd29246,17'd27640,17'd27766,17'd25709,17'd24743,17'd23218,17'd31347,17'd47540,17'd47642,17'd47643,17'd47644,17'd47544,17'd47645,17'd47646,17'd47647,17'd46337,17'd47648,17'd47649,17'd47547,17'd47455,17'd31836,17'd23389,17'd32827,17'd22500,17'd22504,17'd23926,17'd46677,17'd21842,17'd47650,17'd47651,17'd47652,17'd47549,17'd47653,17'd47551,17'd41127,17'd47654,17'd47655,17'd47656,17'd47657,17'd47658,17'd24934,17'd21136,17'd22584,17'd10043,17'd47558,17'd47468,17'd23633,17'd14301,17'd28186,17'd41141,17'd38701,17'd47659,17'd16956,17'd11576,17'd30487,17'd10514,17'd6390,17'd28185,17'd5329,17'd34656,17'd41891,17'd33838,17'd42180,17'd47660,17'd4999,17'd4683,17'd4995,17'd4682,17'd30485,17'd5327,17'd4842,17'd5004,17'd5004,17'd4687,17'd5144,17'd41612,17'd4828,17'd34654,17'd34154,17'd47559,17'd47661,17'd44134,17'd33363,17'd47662,17'd40401,17'd40554,17'd47663,17'd47664,17'd47664,17'd47665,17'd47666,17'd46876,17'd47478,17'd37163,17'd47566,17'd47667,17'd47568,17'd47668,17'd47669,17'd7023,17'd9661,17'd45786,17'd45185,17'd18629,17'd18629,17'd41004,17'd39482,17'd39483,17'd38859,17'd38860,17'd38580,17'd38072,17'd13420,17'd43596,17'd16492,17'd16492,17'd6258,17'd8186,17'd8186,17'd5958,17'd4882,17'd4713,17'd4882,17'd9123,17'd14586,17'd34000,17'd33847,17'd417,17'd194,17'd423,17'd605,17'd410,17'd47670
},
'{
17'd4087,17'd4426,17'd3902,17'd3902,17'd27713,17'd6420,17'd2592,17'd27714,17'd2425,17'd1416,17'd3905,17'd3905,17'd980,17'd27,17'd27,17'd980,17'd652,17'd652,17'd289,17'd30,17'd3256,17'd45516,17'd46358,17'd13303,17'd2428,17'd2261,17'd1971,17'd1282,17'd46793,17'd46885,17'd17079,17'd18150,17'd2610,17'd34168,17'd2797,17'd3447,17'd46887,17'd47271,17'd14329,17'd47671,17'd24010,17'd47488,17'd47672,17'd46359,17'd47273,17'd20292,17'd20148,17'd17206,17'd17445,17'd16034,17'd47490,17'd21964,17'd12531,17'd12815,17'd13211,17'd17096,17'd12361,17'd12530,17'd15137,17'd19890,17'd13599,17'd17096,17'd17204,17'd17207,17'd14346,17'd15900,17'd47572,17'd47572,17'd47572,17'd47673,17'd16030,17'd14474,17'd14475,17'd14100,17'd13466,17'd12959,17'd9007,17'd8538,17'd7750,17'd5689,17'd5253,17'd5252,17'd6137,17'd7259,17'd39647,17'd40271,17'd42063,17'd44283,17'd47575,17'd47576,17'd47577,17'd45199,17'd47674,17'd47675,17'd47676,17'd47677,17'd47678,17'd47679,17'd47680,17'd47681,17'd47682,17'd47683,17'd47684,17'd47685,17'd45929,17'd44405,17'd47686,17'd47687,17'd47688,17'd17850,17'd19780,17'd11531,17'd36073,17'd34695,17'd27006,17'd11401,17'd11400,17'd17966,17'd36349,17'd23166,17'd29783,17'd29928,17'd28110,17'd24856,17'd24857,17'd24031,17'd26495,17'd36346,17'd26871,17'd47009,17'd14259,17'd18327,17'd13516,17'd13516,17'd12996,17'd15053,17'd17603,17'd19407,17'd27121,17'd28571,17'd39211,17'd31763,17'd47403,17'd47295,17'd47594,17'd47593,17'd30072,17'd28571,17'd28816,17'd23856,17'd21362,17'd17478,17'd28463,17'd22820,17'd9884,17'd10024,17'd9885,17'd9885,17'd9885,17'd9885,17'd27003,17'd19918,17'd19415,17'd47689,17'd32942,17'd47690,17'd47691,17'd32141,17'd30986,17'd30089,17'd11665,17'd17720,17'd8723,17'd23342,17'd47692,17'd47693,17'd35528,17'd47694,17'd47695,17'd47696,17'd47302,17'd38918,17'd36224,17'd31625,17'd47205,17'd47601,17'd47697,17'd47698,17'd47699,17'd47700,17'd47701,17'd47702,17'd39716,17'd42422,17'd47703,17'd47704,17'd47705,17'd47706,17'd47705,17'd47704,17'd47707,17'd47708,17'd47709,17'd47710,17'd34420,17'd46743,17'd47711,17'd47711,17'd47712,17'd33618,17'd36099,17'd45860,17'd47221,17'd36523,17'd38644,17'd44465,17'd42581,17'd33916,17'd33769,17'd35407,17'd41716,17'd38645,17'd35972,17'd36385,17'd38645,17'd35971,17'd35971,17'd36245,17'd36245,17'd35971,17'd36384,17'd36244,17'd36244,17'd36670,17'd38391,17'd36669,17'd37634,17'd37634,17'd37634,17'd37634,17'd46937,17'd37635,17'd37365,17'd47713,17'd47714,17'd47715,17'd47716,17'd47717,17'd46315,17'd47718,17'd47719,17'd47720,17'd47721,17'd47722,17'd47723,17'd47724,17'd47725,17'd47050,17'd46663,17'd47726,17'd46093,17'd44938,17'd44700,17'd44827,17'd40825,17'd42599,17'd44934,17'd43979,17'd47727,17'd47727,17'd37778,17'd33643,17'd25317,17'd27512,17'd25180,17'd29688,17'd23565,17'd37386,17'd23389,17'd32827,17'd22329,17'd41273,17'd37386,17'd23733,17'd34282,17'd28254,17'd46549,17'd28602,17'd25707,17'd43695,17'd46752,17'd47728,17'd44593,17'd47729,17'd47143,17'd45483,17'd44698,17'd47730,17'd42882,17'd36983,17'd35425,17'd40367,17'd31354,17'd28727,17'd26781,17'd35023,17'd27371,17'd28725,17'd26903,17'd26174,17'd28720,17'd27882,17'd28974,17'd28718,17'd34884,17'd24742,17'd28368,17'd32007,17'd30432,17'd47731,17'd25709,17'd28253,17'd26062,17'd27515,17'd26902,17'd35426,17'd31503,17'd37513,17'd27885,17'd36541,17'd44594,17'd45483,17'd46661,17'd47636,17'd47637,17'd47732,17'd47733,17'd47734,17'd47734,17'd47735,17'd47736,17'd47737,17'd47054,17'd45879,17'd39738,17'd46425,17'd37908,17'd29245,17'd27640,17'd28602,17'd25709,17'd24415,17'd23389,17'd31347,17'd22866,17'd47642,17'd47738,17'd47739,17'd47740,17'd47741,17'd47742,17'd47743,17'd47744,17'd47648,17'd47649,17'd47547,17'd47745,17'd34277,17'd46669,17'd44702,17'd22330,17'd22504,17'd32350,17'd33312,17'd47746,17'd47747,17'd47748,17'd47749,17'd47750,17'd47751,17'd47752,17'd47753,17'd47754,17'd47755,17'd47756,17'd47075,17'd46782,17'd47757,17'd21762,17'd24303,17'd27305,17'd24150,17'd47758,17'd24945,17'd12467,17'd16615,17'd36310,17'd38701,17'd47659,17'd28186,17'd10514,17'd30487,17'd28184,17'd6390,17'd27935,17'd5329,17'd34656,17'd33838,17'd4359,17'd42180,17'd47660,17'd41459,17'd4683,17'd4995,17'd4682,17'd38442,17'd4995,17'd4842,17'd5004,17'd5004,17'd4686,17'd4991,17'd4185,17'd4828,17'd34654,17'd47759,17'd47559,17'd47661,17'd47760,17'd42184,17'd47761,17'd47762,17'd40554,17'd47665,17'd47664,17'd39475,17'd47665,17'd46986,17'd47763,17'd46694,17'd37163,17'd47764,17'd34662,17'd47765,17'd47766,17'd3551,17'd7340,17'd5351,17'd10071,17'd45185,17'd18629,17'd10388,17'd47767,17'd39482,17'd40101,17'd38859,17'd38860,17'd38580,17'd44019,17'd13420,17'd43596,17'd43596,17'd16492,17'd6258,17'd8186,17'd9123,17'd4882,17'd4882,17'd4713,17'd5940,17'd16256,17'd15233,17'd33847,17'd33847,17'd1672,17'd194,17'd952,17'd971,17'd803,17'd47670
},
'{
17'd4087,17'd4426,17'd4244,17'd4892,17'd29897,17'd14743,17'd3250,17'd27714,17'd2425,17'd1416,17'd3905,17'd18,17'd980,17'd27,17'd27,17'd980,17'd652,17'd29,17'd809,17'd31,17'd2940,17'd45516,17'd3103,17'd13303,17'd2261,17'd2261,17'd1971,17'd1838,17'd21949,17'd19609,17'd992,17'd18150,17'd2610,17'd34168,17'd2797,17'd28197,17'd46481,17'd42198,17'd14329,17'd47768,17'd27104,17'd47488,17'd47672,17'd46359,17'd47571,17'd19006,17'd19893,17'd17206,17'd17445,17'd16034,17'd47490,17'd21649,17'd12531,17'd12815,17'd17096,17'd23154,17'd11764,17'd12361,17'd14764,17'd19890,17'd13599,17'd29904,17'd19893,17'd17445,17'd14893,17'd16166,17'd47769,17'd47769,17'd47769,17'd15900,17'd16030,17'd15641,17'd14473,17'd14100,17'd13466,17'd13468,17'd9704,17'd8538,17'd10430,17'd5255,17'd5253,17'd5252,17'd6137,17'd7259,17'd39647,17'd40271,17'd42063,17'd44283,17'd46898,17'd47770,17'd47771,17'd45199,17'd47674,17'd47675,17'd47676,17'd47772,17'd47773,17'd29911,17'd47774,17'd47775,17'd47776,17'd47777,17'd47778,17'd47099,17'd47779,17'd47780,17'd47781,17'd47687,17'd17851,17'd15056,17'd10028,17'd11967,17'd35096,17'd34695,17'd46809,17'd20045,17'd45208,17'd36349,17'd36349,17'd47782,17'd29783,17'd24539,17'd26149,17'd24537,17'd24857,17'd26871,17'd36479,17'd35800,17'd36346,17'd47009,17'd28112,17'd17478,17'd13516,17'd13645,17'd16204,17'd11806,17'd12719,17'd17348,17'd24991,17'd28818,17'd31587,17'd31761,17'd31763,17'd47403,17'd47783,17'd47784,17'd31764,17'd29645,17'd28943,17'd25672,17'd25926,17'd14259,17'd18326,17'd13647,17'd17847,17'd9884,17'd9885,17'd9885,17'd9741,17'd9885,17'd27003,17'd25529,17'd9343,17'd47785,17'd39830,17'd34838,17'd47691,17'd47598,17'd32296,17'd32610,17'd29341,17'd10606,17'd47786,17'd47787,17'd47788,17'd47789,17'd35383,17'd47694,17'd47790,17'd47791,17'd47603,17'd47303,17'd40893,17'd46918,17'd47205,17'd47792,17'd46814,17'd47793,17'd47794,17'd47795,17'd47796,17'd47797,17'd46515,17'd47798,17'd47799,17'd47704,17'd47705,17'd47706,17'd47800,17'd47705,17'd44217,17'd47801,17'd47802,17'd47803,17'd47804,17'd35685,17'd47805,17'd47806,17'd35408,17'd40033,17'd36099,17'd47221,17'd38644,17'd46931,17'd46931,17'd42581,17'd42135,17'd35678,17'd37101,17'd33620,17'd36965,17'd36246,17'd36965,17'd35273,17'd35407,17'd33620,17'd36247,17'd33620,17'd36247,17'd36965,17'd35971,17'd35972,17'd36385,17'd36384,17'd36670,17'd38391,17'd36669,17'd36669,17'd36669,17'd36669,17'd47807,17'd47808,17'd46936,17'd47809,17'd47810,17'd47811,17'd47812,17'd47813,17'd46541,17'd47814,17'd47815,17'd47816,17'd47817,17'd47818,17'd47819,17'd47638,17'd44474,17'd40364,17'd46556,17'd44356,17'd39129,17'd43426,17'd46200,17'd40825,17'd40959,17'd43287,17'd43695,17'd43979,17'd47438,17'd47727,17'd32996,17'd28721,17'd27882,17'd27512,17'd25030,17'd23916,17'd23566,17'd37386,17'd23218,17'd22329,17'd23218,17'd39278,17'd29827,17'd30431,17'd29533,17'd47820,17'd39444,17'd25708,17'd32995,17'd44104,17'd46947,17'd44224,17'd44102,17'd47821,17'd47821,17'd47822,17'd44828,17'd47823,17'd44234,17'd37907,17'd35425,17'd32831,17'd31503,17'd28979,17'd26781,17'd35023,17'd27371,17'd28725,17'd26903,17'd26174,17'd28594,17'd28717,17'd28485,17'd27763,17'd28718,17'd24895,17'd32668,17'd25179,17'd31034,17'd47824,17'd28720,17'd28252,17'd26530,17'd28725,17'd28486,17'd39437,17'd30279,17'd33952,17'd27885,17'd41731,17'd42889,17'd46660,17'd46756,17'd47237,17'd47444,17'd47825,17'd47826,17'd45607,17'd47827,17'd47828,17'd47736,17'd47737,17'd47054,17'd45987,17'd39738,17'd46425,17'd35426,17'd29245,17'd27883,17'd28723,17'd25438,17'd24090,17'd23389,17'd31347,17'd22866,17'd47829,17'd47541,17'd47738,17'd47830,17'd47831,17'd45991,17'd47832,17'd46114,17'd45997,17'd47833,17'd47547,17'd47745,17'd32679,17'd32015,17'd45754,17'd22330,17'd22504,17'd32350,17'd47834,17'd47835,17'd47836,17'd47837,17'd47838,17'd47839,17'd47840,17'd47752,17'd47841,17'd47842,17'd47843,17'd47844,17'd47845,17'd47846,17'd19337,17'd47847,17'd47848,17'd23458,17'd24150,17'd47758,17'd24945,17'd12467,17'd16615,17'd38701,17'd38701,17'd47370,17'd15727,17'd10641,17'd30487,17'd28184,17'd6554,17'd27935,17'd5329,17'd4529,17'd33841,17'd33838,17'd42180,17'd47660,17'd41459,17'd4683,17'd4995,17'd4682,17'd30486,17'd5327,17'd4842,17'd30637,17'd5004,17'd4687,17'd38442,17'd41455,17'd4828,17'd34654,17'd47759,17'd47849,17'd5601,17'd4179,17'd5473,17'd41146,17'd34497,17'd47850,17'd47851,17'd47852,17'd47852,17'd40254,17'd47853,17'd47474,17'd46694,17'd37038,17'd47854,17'd47855,17'd47856,17'd47857,17'd47858,17'd47859,17'd5351,17'd10071,17'd45185,17'd18629,17'd10388,17'd47767,17'd39482,17'd39483,17'd38859,17'd38860,17'd38580,17'd44019,17'd12913,17'd43596,17'd43596,17'd16492,17'd6258,17'd8186,17'd9123,17'd4882,17'd4882,17'd4713,17'd4882,17'd9123,17'd14586,17'd28428,17'd2560,17'd1671,17'd415,17'd952,17'd1963,17'd271,17'd47670
},
'{
17'd3902,17'd3902,17'd4428,17'd4428,17'd15358,17'd2935,17'd2781,17'd10535,17'd2425,17'd1416,17'd18,17'd18,17'd980,17'd27,17'd27,17'd27,17'd652,17'd652,17'd289,17'd30,17'd291,17'd2259,17'd1130,17'd656,17'd13303,17'd2261,17'd1971,17'd1282,17'd19499,17'd47860,17'd1139,17'd35772,17'd1707,17'd34168,17'd2797,17'd28197,17'd47861,17'd47862,17'd19509,17'd47768,17'd27104,17'd47488,17'd47272,17'd46359,17'd47571,17'd19006,17'd19893,17'd17206,17'd18657,17'd16034,17'd47490,17'd21649,17'd12532,17'd12815,17'd17096,17'd17096,17'd13969,17'd12530,17'd15137,17'd14890,17'd13599,17'd17096,17'd17204,17'd47863,17'd32739,17'd15767,17'd15900,17'd15900,17'd47864,17'd47864,17'd47865,17'd47866,17'd47867,17'd47868,17'd47869,17'd47870,17'd9007,17'd8538,17'd10430,17'd7750,17'd5255,17'd5252,17'd6137,17'd7259,17'd39647,17'd40271,17'd47871,17'd47872,17'd46898,17'd47576,17'd47577,17'd45199,17'd47873,17'd47874,17'd47875,17'd47876,17'd47877,17'd29768,17'd47878,17'd47879,17'd47880,17'd47778,17'd47778,17'd47585,17'd47881,17'd45679,17'd47882,17'd47290,17'd34694,17'd12265,17'd8580,17'd11811,17'd47883,17'd34541,17'd46809,17'd19919,17'd12423,17'd34205,17'd36349,17'd47884,17'd36348,17'd24539,17'd24208,17'd26149,17'd24538,17'd26495,17'd35800,17'd47885,17'd47886,17'd34832,17'd24363,17'd17478,17'd13645,17'd20451,17'd13362,17'd11806,17'd11958,17'd17348,17'd23511,17'd28460,17'd30072,17'd31761,17'd31761,17'd47887,17'd47888,17'd47403,17'd47295,17'd34551,17'd28461,17'd26872,17'd24705,17'd24995,17'd21985,17'd13521,17'd22820,17'd9884,17'd9885,17'd9885,17'd17011,17'd10742,17'd10742,17'd27856,17'd47889,17'd47890,17'd47891,17'd39515,17'd47892,17'd32297,17'd47893,17'd32775,17'd29341,17'd25928,17'd47786,17'd43763,17'd47894,17'd47895,17'd37212,17'd47896,17'd47897,17'd47898,17'd47603,17'd47409,17'd35660,17'd35661,17'd47307,17'd47792,17'd47899,17'd47900,17'd47901,17'd47902,17'd47903,17'd47613,17'd47904,17'd47905,17'd47906,17'd43003,17'd47907,17'd47908,17'd34073,17'd47909,17'd47910,17'd38952,17'd47802,17'd35126,17'd36238,17'd38638,17'd47911,17'd38387,17'd42865,17'd42865,17'd47912,17'd40502,17'd47221,17'd36523,17'd38644,17'd38644,17'd42581,17'd36378,17'd36969,17'd34076,17'd35834,17'd35274,17'd34076,17'd37235,17'd33769,17'd37101,17'd37235,17'd35274,17'd35834,17'd41716,17'd36965,17'd36246,17'd36245,17'd35971,17'd36384,17'd36244,17'd36244,17'd36244,17'd36670,17'd38391,17'd47913,17'd47914,17'd47713,17'd47915,17'd47916,17'd47917,17'd47717,17'd47918,17'd39412,17'd45146,17'd47919,17'd47920,17'd47921,17'd47922,17'd47923,17'd47924,17'd44931,17'd40216,17'd47925,17'd47926,17'd41416,17'd44935,17'd46200,17'd40959,17'd43287,17'd47927,17'd46095,17'd46095,17'd43978,17'd47438,17'd32996,17'd28721,17'd28717,17'd25178,17'd24745,17'd30879,17'd23386,17'd23215,17'd23218,17'd30277,17'd23216,17'd38976,17'd23918,17'd34621,17'd24898,17'd47928,17'd30734,17'd35012,17'd44699,17'd39738,17'd47929,17'd47930,17'd42146,17'd47931,17'd47931,17'd43973,17'd42878,17'd41994,17'd43692,17'd40824,17'd35990,17'd40367,17'd31352,17'd28979,17'd26781,17'd33963,17'd26782,17'd28853,17'd26903,17'd27766,17'd25567,17'd27512,17'd28485,17'd38407,17'd24745,17'd25031,17'd31034,17'd27511,17'd25317,17'd39283,17'd25707,17'd28978,17'd27883,17'd27027,17'd30735,17'd31354,17'd33319,17'd33001,17'd32832,17'd41429,17'd44235,17'd47932,17'd47933,17'd47934,17'd47536,17'd47935,17'd47827,17'd46321,17'd46321,17'd47936,17'd43281,17'd47937,17'd47828,17'd47938,17'd44226,17'd41270,17'd35426,17'd28727,17'd27883,17'd28723,17'd25177,17'd23731,17'd41273,17'd31347,17'd47939,17'd47829,17'd47448,17'd47541,17'd47940,17'd47941,17'd47942,17'd47943,17'd45761,17'd47944,17'd47753,17'd45378,17'd34453,17'd32015,17'd45754,17'd34278,17'd22331,17'd22500,17'd23393,17'd31192,17'd21840,17'd47945,17'd47946,17'd47947,17'd47948,17'd47949,17'd47950,17'd40834,17'd47951,17'd47952,17'd47953,17'd47954,17'd47955,17'd47956,17'd47957,17'd25081,17'd7660,17'd5916,17'd24483,17'd24945,17'd12467,17'd12906,17'd38701,17'd36171,17'd24803,17'd16615,17'd28184,17'd30487,17'd30487,17'd6554,17'd27935,17'd5329,17'd4529,17'd4189,17'd4359,17'd42180,17'd47660,17'd5155,17'd4841,17'd4683,17'd4682,17'd38442,17'd4683,17'd4842,17'd5004,17'd25627,17'd4687,17'd4991,17'd4185,17'd40848,17'd47958,17'd34495,17'd47959,17'd47960,17'd47661,17'd4824,17'd47959,17'd47961,17'd47962,17'd3841,17'd40089,17'd40089,17'd40254,17'd47963,17'd47373,17'd46694,17'd47964,17'd45781,17'd47965,17'd47966,17'd47967,17'd47858,17'd46882,17'd9789,17'd10071,17'd46354,17'd18629,17'd10388,17'd47767,17'd39482,17'd39483,17'd38859,17'd38860,17'd38580,17'd44019,17'd12913,17'd13176,17'd13176,17'd16492,17'd6258,17'd7365,17'd5776,17'd4882,17'd4882,17'd4713,17'd5940,17'd16256,17'd15233,17'd29440,17'd2560,17'd941,17'd2763,17'd952,17'd1963,17'd261,17'd802
},
'{
17'd4244,17'd3902,17'd4428,17'd4428,17'd3428,17'd2935,17'd2781,17'd10535,17'd2257,17'd1416,17'd18,17'd18,17'd980,17'd27,17'd27,17'd27,17'd652,17'd29,17'd809,17'd31,17'd982,17'd32,17'd656,17'd656,17'd13303,17'd1968,17'd47968,17'd1838,17'd1134,17'd46793,17'd16967,17'd35772,17'd1707,17'd35620,17'd13072,17'd28197,17'd47969,17'd44619,17'd47970,17'd28666,17'd27104,17'd47488,17'd47272,17'd46359,17'd47571,17'd19006,17'd19893,17'd17206,17'd18657,17'd16034,17'd47274,17'd21649,17'd12532,17'd12815,17'd17096,17'd34015,17'd11764,17'd12361,17'd14764,17'd14890,17'd13599,17'd29904,17'd19893,17'd17690,17'd15008,17'd15767,17'd15900,17'd16166,17'd47865,17'd47865,17'd47971,17'd47972,17'd47973,17'd47974,17'd47868,17'd47975,17'd9704,17'd7582,17'd10430,17'd7750,17'd5255,17'd5252,17'd6137,17'd7259,17'd39647,17'd40271,17'd47871,17'd47872,17'd46898,17'd47576,17'd47577,17'd45199,17'd47873,17'd47976,17'd47977,17'd47876,17'd47978,17'd47979,17'd47980,17'd47981,17'd47982,17'd47983,17'd47984,17'd47985,17'd46374,17'd47986,17'd47987,17'd47988,17'd47989,17'd10860,17'd17483,17'd24213,17'd47883,17'd34541,17'd46809,17'd20045,17'd47990,17'd34205,17'd47991,17'd47884,17'd47992,17'd47993,17'd47009,17'd28110,17'd26149,17'd26495,17'd35800,17'd37200,17'd47994,17'd34832,17'd24363,17'd17478,17'd19533,17'd14522,17'd12262,17'd12861,17'd12113,17'd16321,17'd12255,17'd28103,17'd28686,17'd31439,17'd31762,17'd31762,17'd47888,17'd47403,17'd47295,17'd34551,17'd31768,17'd28104,17'd23856,17'd24362,17'd23513,17'd28463,17'd11526,17'd19278,17'd10169,17'd9885,17'd17011,17'd10742,17'd10743,17'd27856,17'd47889,17'd47995,17'd47996,17'd47997,17'd30091,17'd47998,17'd47999,17'd48000,17'd11665,17'd45549,17'd48001,17'd48002,17'd48003,17'd48004,17'd47698,17'd48005,17'd48006,17'd48007,17'd48008,17'd40449,17'd46386,17'd48009,17'd48010,17'd48010,17'd48011,17'd48012,17'd48013,17'd42084,17'd48014,17'd48015,17'd48016,17'd48017,17'd48018,17'd46826,17'd48019,17'd48020,17'd46414,17'd47909,17'd48021,17'd48022,17'd38775,17'd38777,17'd46929,17'd48023,17'd48024,17'd48024,17'd42865,17'd36238,17'd36238,17'd46313,17'd33618,17'd40502,17'd47033,17'd36249,17'd47035,17'd36523,17'd42581,17'd34994,17'd36969,17'd35678,17'd33916,17'd34994,17'd33769,17'd33769,17'd37101,17'd35274,17'd36247,17'd36965,17'd36246,17'd41716,17'd36965,17'd38645,17'd36385,17'd36385,17'd35972,17'd35971,17'd35972,17'd38958,17'd48025,17'd48026,17'd47808,17'd46938,17'd48027,17'd48028,17'd47813,17'd37365,17'd46418,17'd39263,17'd48029,17'd48030,17'd48031,17'd48032,17'd48033,17'd48034,17'd44472,17'd47628,17'd46204,17'd48035,17'd41863,17'd43289,17'd43980,17'd40959,17'd43288,17'd33155,17'd43837,17'd46095,17'd37778,17'd47438,17'd37778,17'd43022,17'd25568,17'd29976,17'd24416,17'd30275,17'd29686,17'd23215,17'd30277,17'd22501,17'd38976,17'd30278,17'd24086,17'd33793,17'd48036,17'd31856,17'd25708,17'd46095,17'd48037,17'd44472,17'd48038,17'd47930,17'd44932,17'd47728,17'd48039,17'd44821,17'd48040,17'd48041,17'd46752,17'd43700,17'd48042,17'd40367,17'd29246,17'd28979,17'd26901,17'd33963,17'd26902,17'd28853,17'd27515,17'd28602,17'd28597,17'd28719,17'd28485,17'd38407,17'd25180,17'd32353,17'd39591,17'd27765,17'd28594,17'd48043,17'd27258,17'd27027,17'd43290,17'd28486,17'd31352,17'd32356,17'd32354,17'd33001,17'd32356,17'd34877,17'd44227,17'd48044,17'd48045,17'd47443,17'd48046,17'd48047,17'd48048,17'd48049,17'd48049,17'd47538,17'd43281,17'd47937,17'd47828,17'd47938,17'd47726,17'd43019,17'd32016,17'd28727,17'd33815,17'd28720,17'd25177,17'd30879,17'd41273,17'd31347,17'd47939,17'd48050,17'd47448,17'd47448,17'd48051,17'd48052,17'd48053,17'd48054,17'd44837,17'd40834,17'd43856,17'd45378,17'd47159,17'd32015,17'd40529,17'd44489,17'd44702,17'd22500,17'd32503,17'd31346,17'd48055,17'd48056,17'd48057,17'd48058,17'd32499,17'd48059,17'd47950,17'd44837,17'd48060,17'd48061,17'd48062,17'd48063,17'd48064,17'd19820,17'd48065,17'd25221,17'd48066,17'd5916,17'd24483,17'd14301,17'd11710,17'd12906,17'd36171,17'd36171,17'd24803,17'd16615,17'd28184,17'd30179,17'd30487,17'd31717,17'd27935,17'd5002,17'd4689,17'd33841,17'd33838,17'd42180,17'd46979,17'd5155,17'd4841,17'd5328,17'd4995,17'd30486,17'd5328,17'd4842,17'd5004,17'd25627,17'd4845,17'd5144,17'd41455,17'd4829,17'd47958,17'd48067,17'd47959,17'd5474,17'd47960,17'd47960,17'd48068,17'd4826,17'd48069,17'd48070,17'd48071,17'd40089,17'd40404,17'd47853,17'd46876,17'd47478,17'd48072,17'd44739,17'd47965,17'd48073,17'd48074,17'd47269,17'd8480,17'd9789,17'd46477,17'd18629,17'd10388,17'd10388,17'd47767,17'd39482,17'd39483,17'd38859,17'd38860,17'd38580,17'd44019,17'd12913,17'd13176,17'd13176,17'd16492,17'd6258,17'd7365,17'd5776,17'd4882,17'd4882,17'd4713,17'd4882,17'd9123,17'd14586,17'd34000,17'd1672,17'd421,17'd602,17'd192,17'd1963,17'd47670,17'd802
},
'{
17'd4244,17'd4244,17'd4088,17'd4245,17'd34512,17'd3252,17'd1689,17'd2594,17'd22965,17'd17,17'd18,17'd18,17'd980,17'd27,17'd27,17'd27,17'd19,17'd18,17'd289,17'd30,17'd291,17'd2259,17'd32,17'd656,17'd2260,17'd13303,17'd22615,17'd1282,17'd19499,17'd19499,17'd1138,17'd35772,17'd1707,17'd35620,17'd36605,17'd48075,17'd44389,17'd25654,17'd24970,17'd29046,17'd18288,17'd48076,17'd47272,17'd48077,17'd47571,17'd19006,17'd17689,17'd17206,17'd17207,17'd16169,17'd47863,17'd19754,17'd12531,17'd12362,17'd23325,17'd17096,17'd12361,17'd12530,17'd15137,17'd19890,17'd12954,17'd23325,17'd17204,17'd47863,17'd14767,17'd16029,17'd15767,17'd16166,17'd48078,17'd48079,17'd48080,17'd33857,17'd47973,17'd48081,17'd47868,17'd47975,17'd9704,17'd8538,17'd10430,17'd7750,17'd6626,17'd6305,17'd6138,17'd7422,17'd6782,17'd6484,17'd41782,17'd48082,17'd46898,17'd48083,17'd47577,17'd45669,17'd40278,17'd48084,17'd48085,17'd48086,17'd48087,17'd48088,17'd48089,17'd48090,17'd48091,17'd48092,17'd48093,17'd47778,17'd48094,17'd46145,17'd48095,17'd48096,17'd48097,17'd7788,17'd17850,17'd8248,17'd34699,17'd22645,17'd46613,17'd12585,17'd11525,17'd13368,17'd47782,17'd47884,17'd36626,17'd24993,17'd24208,17'd28231,17'd24208,17'd26496,17'd35800,17'd48098,17'd48099,17'd48100,17'd28947,17'd14264,17'd11397,17'd48101,17'd15810,17'd12861,17'd12111,17'd16321,17'd19407,17'd27121,17'd28461,17'd30676,17'd31762,17'd31762,17'd47887,17'd31763,17'd39211,17'd31587,17'd29067,17'd28345,17'd26370,17'd24992,17'd24858,17'd12583,17'd11525,17'd10330,17'd9884,17'd9885,17'd10742,17'd17011,17'd9479,17'd27856,17'd9336,17'd48102,17'd48103,17'd39665,17'd48104,17'd32298,17'd30091,17'd48105,17'd10853,17'd15943,17'd8568,17'd48106,17'd48107,17'd48108,17'd48109,17'd48110,17'd48111,17'd48112,17'd48113,17'd48114,17'd48114,17'd48115,17'd48116,17'd46619,17'd48117,17'd48118,17'd48119,17'd48120,17'd48121,17'd48122,17'd48123,17'd48124,17'd48125,17'd46523,17'd48126,17'd48127,17'd48128,17'd48129,17'd41255,17'd41255,17'd48130,17'd48131,17'd38005,17'd33616,17'd48132,17'd48133,17'd33766,17'd34074,17'd33766,17'd45471,17'd46313,17'd40033,17'd47912,17'd33618,17'd36099,17'd36249,17'd36523,17'd44465,17'd42581,17'd42581,17'd42581,17'd42135,17'd35678,17'd36969,17'd33769,17'd37101,17'd35407,17'd41716,17'd36246,17'd36965,17'd36965,17'd36245,17'd35972,17'd36385,17'd35971,17'd36245,17'd35972,17'd36669,17'd48134,17'd47808,17'd46937,17'd48135,17'd48136,17'd37761,17'd48137,17'd48138,17'd46652,17'd48139,17'd46942,17'd48140,17'd48141,17'd48142,17'd48143,17'd48144,17'd45370,17'd44226,17'd48145,17'd45745,17'd44227,17'd43298,17'd45484,17'd42598,17'd43288,17'd47927,17'd47727,17'd47629,17'd33157,17'd43286,17'd33157,17'd42749,17'd25178,17'd25031,17'd24090,17'd34137,17'd23387,17'd23215,17'd30277,17'd23217,17'd36987,17'd29242,17'd30733,17'd25180,17'd47820,17'd28721,17'd32995,17'd43018,17'd48146,17'd48147,17'd48148,17'd43972,17'd44100,17'd42594,17'd43283,17'd46946,17'd48149,17'd46438,17'd44821,17'd47439,17'd37907,17'd31503,17'd29246,17'd28726,17'd26781,17'd26781,17'd26902,17'd28724,17'd25833,17'd28720,17'd28717,17'd25029,17'd28595,17'd24897,17'd29976,17'd29244,17'd29970,17'd28594,17'd25833,17'd33815,17'd35011,17'd26781,17'd28486,17'd30735,17'd27642,17'd32832,17'd32192,17'd33319,17'd39743,17'd41109,17'd45482,17'd48150,17'd48151,17'd47534,17'd47935,17'd48152,17'd48049,17'd48153,17'd48153,17'd47736,17'd48154,17'd47737,17'd48155,17'd48156,17'd48157,17'd43019,17'd37908,17'd26901,17'd26530,17'd28594,17'd29244,17'd28722,17'd41273,17'd38041,17'd47939,17'd47829,17'd48158,17'd48159,17'd46968,17'd45766,17'd35320,17'd44708,17'd38685,17'd40971,17'd34139,17'd48160,17'd45492,17'd44702,17'd44489,17'd44489,17'd30428,17'd22856,17'd32666,17'd48161,17'd48162,17'd48163,17'd21702,17'd48164,17'd32498,17'd46677,17'd48165,17'd45271,17'd48166,17'd48167,17'd48168,17'd48169,17'd48170,17'd48171,17'd48172,17'd26583,17'd6383,17'd5332,17'd48173,17'd29297,17'd12760,17'd12761,17'd38701,17'd38316,17'd36028,17'd14423,17'd30179,17'd30179,17'd28058,17'd27935,17'd5160,17'd5329,17'd4840,17'd5144,17'd34157,17'd34157,17'd38442,17'd42910,17'd4841,17'd4840,17'd4682,17'd5144,17'd4840,17'd5002,17'd5004,17'd25627,17'd4687,17'd4991,17'd4016,17'd4829,17'd35889,17'd48174,17'd48175,17'd47559,17'd4983,17'd48176,17'd48177,17'd48178,17'd48179,17'd48180,17'd48181,17'd48071,17'd47851,17'd47963,17'd46786,17'd47478,17'd48182,17'd48183,17'd48184,17'd2883,17'd48185,17'd4050,17'd48186,17'd5626,17'd41002,17'd18629,17'd10388,17'd10388,17'd47767,17'd39482,17'd39483,17'd39033,17'd38580,17'd38580,17'd38580,17'd44019,17'd13176,17'd48187,17'd6094,17'd6258,17'd7365,17'd5776,17'd5958,17'd4882,17'd4713,17'd5940,17'd14178,17'd2098,17'd15233,17'd2394,17'd415,17'd203,17'd1409,17'd272,17'd262,17'd2115
},
'{
17'd4244,17'd4244,17'd4088,17'd4245,17'd34512,17'd2422,17'd1967,17'd2594,17'd22965,17'd17,17'd18,17'd18,17'd980,17'd27,17'd27,17'd27,17'd18,17'd16,17'd809,17'd31,17'd982,17'd32,17'd33,17'd656,17'd2939,17'd13303,17'd22615,17'd1838,17'd1134,17'd19499,17'd1138,17'd35772,17'd1707,17'd35620,17'd36605,17'd23661,17'd43597,17'd48188,17'd19886,17'd29046,17'd18288,17'd48076,17'd47272,17'd48077,17'd47571,17'd19006,17'd17689,17'd17318,17'd46889,17'd16169,17'd47863,17'd19754,17'd12531,17'd12218,17'd12813,17'd23154,17'd11913,17'd12530,17'd14890,17'd13210,17'd12954,17'd23325,17'd17204,17'd47863,17'd32739,17'd33548,17'd16029,17'd15767,17'd48079,17'd48189,17'd48080,17'd34178,17'd47971,17'd47973,17'd47974,17'd48190,17'd9704,17'd9007,17'd10430,17'd5409,17'd6626,17'd11089,17'd6138,17'd7422,17'd6782,17'd6484,17'd48191,17'd48082,17'd47575,17'd48083,17'd45668,17'd48192,17'd48193,17'd48084,17'd48085,17'd7930,17'd48087,17'd48088,17'd48194,17'd48195,17'd48196,17'd48093,17'd27471,17'd48197,17'd48198,17'd47881,17'd48199,17'd48200,17'd47398,17'd17851,17'd12120,17'd8419,17'd30217,17'd29334,17'd17601,17'd37735,17'd20046,17'd13368,17'd47782,17'd47884,17'd36626,17'd48201,17'd27985,17'd28231,17'd24208,17'd27985,17'd33572,17'd48202,17'd48203,17'd46050,17'd45684,17'd29783,17'd21985,17'd48204,17'd10989,17'd12861,17'd11961,17'd16321,17'd19407,17'd23511,17'd28818,17'd31440,17'd30834,17'd31762,17'd31761,17'd31761,17'd39211,17'd39211,17'd31587,17'd28461,17'd28816,17'd24030,17'd21363,17'd18327,17'd28463,17'd11526,17'd9884,17'd9741,17'd10742,17'd17011,17'd9479,17'd16554,17'd9469,17'd48205,17'd48206,17'd48207,17'd48208,17'd48209,17'd48210,17'd39515,17'd20910,17'd15181,17'd47786,17'd48211,17'd48212,17'd48213,17'd48214,17'd48215,17'd48216,17'd48217,17'd48218,17'd44411,17'd44411,17'd48219,17'd48220,17'd48221,17'd48222,17'd48117,17'd48223,17'd48224,17'd48225,17'd48226,17'd48227,17'd48228,17'd48229,17'd48230,17'd48231,17'd48232,17'd48233,17'd48234,17'd46518,17'd48235,17'd48236,17'd48237,17'd47128,17'd48238,17'd48239,17'd48240,17'd48241,17'd48242,17'd40198,17'd33766,17'd36238,17'd42865,17'd46313,17'd47912,17'd33915,17'd47033,17'd47221,17'd36523,17'd44465,17'd44465,17'd38644,17'd46931,17'd46931,17'd33916,17'd34994,17'd33769,17'd34076,17'd33620,17'd36247,17'd35834,17'd35273,17'd36246,17'd36245,17'd36246,17'd36246,17'd38645,17'd36384,17'd39416,17'd48243,17'd47913,17'd47810,17'd46537,17'd48244,17'd47809,17'd48245,17'd48246,17'd48247,17'd48248,17'd48249,17'd48250,17'd48251,17'd48252,17'd48253,17'd48254,17'd43973,17'd48255,17'd48256,17'd44228,17'd43021,17'd44827,17'd40218,17'd41111,17'd42437,17'd43838,17'd47438,17'd47727,17'd43550,17'd44359,17'd33157,17'd29825,17'd25178,17'd24895,17'd23731,17'd34137,17'd23388,17'd32351,17'd22501,17'd23216,17'd48257,17'd31033,17'd34276,17'd28974,17'd33484,17'd37778,17'd45749,17'd48258,17'd47924,17'd48259,17'd39431,17'd43689,17'd44099,17'd48041,17'd39580,17'd39735,17'd41265,17'd42295,17'd44100,17'd45481,17'd40961,17'd31503,17'd28980,17'd28726,17'd26781,17'd26902,17'd28853,17'd28724,17'd25708,17'd28594,17'd28717,17'd25029,17'd34283,17'd24898,17'd25178,17'd27511,17'd28723,17'd28481,17'd27259,17'd35723,17'd31352,17'd28726,17'd28727,17'd31352,17'd30279,17'd28373,17'd33654,17'd32354,17'd36541,17'd40958,17'd48035,17'd46760,17'd48260,17'd47534,17'd47935,17'd48261,17'd46199,17'd48262,17'd48262,17'd43281,17'd48263,17'd48264,17'd47343,17'd48265,17'd48266,17'd41111,17'd35426,17'd26781,17'd26530,17'd28594,17'd25320,17'd30275,17'd32827,17'd38041,17'd47939,17'd48267,17'd48268,17'd48052,17'd48269,17'd48270,17'd35456,17'd48271,17'd40065,17'd34139,17'd48272,17'd48160,17'd23391,17'd44591,17'd48273,17'd43854,17'd34619,17'd22332,17'd32666,17'd48274,17'd42441,17'd48275,17'd48276,17'd48277,17'd23041,17'd48278,17'd48279,17'd34640,17'd48280,17'd48281,17'd48282,17'd48283,17'd48284,17'd22733,17'd48285,17'd26584,17'd5914,17'd5332,17'd48173,17'd14301,17'd29161,17'd16615,17'd36171,17'd38191,17'd28059,17'd12906,17'd10514,17'd30179,17'd28058,17'd6554,17'd30638,17'd5329,17'd4840,17'd5144,17'd34157,17'd4998,17'd30486,17'd42910,17'd4841,17'd4841,17'd4995,17'd5153,17'd4841,17'd5002,17'd5004,17'd25627,17'd4687,17'd4997,17'd41612,17'd4829,17'd35889,17'd48174,17'd4352,17'd47849,17'd48176,17'd48068,17'd47759,17'd47372,17'd39776,17'd39471,17'd48286,17'd3837,17'd47851,17'd47853,17'd48287,17'd46694,17'd48182,17'd48288,17'd48289,17'd48290,17'd3551,17'd48291,17'd5024,17'd5493,17'd41002,17'd18629,17'd10388,17'd10388,17'd47767,17'd39482,17'd39483,17'd39033,17'd38580,17'd38580,17'd38580,17'd13420,17'd14060,17'd14060,17'd6258,17'd6258,17'd7365,17'd5776,17'd5958,17'd4882,17'd4713,17'd4882,17'd3073,17'd2098,17'd15233,17'd15233,17'd1529,17'd1408,17'd26595,17'd271,17'd408,17'd2115
},
'{
17'd4892,17'd4892,17'd4245,17'd4245,17'd3251,17'd2422,17'd1967,17'd2594,17'd22965,17'd17,17'd652,17'd980,17'd980,17'd27,17'd27,17'd27,17'd18,17'd18,17'd289,17'd30,17'd1129,17'd982,17'd32,17'd656,17'd2939,17'd13303,17'd2121,17'd16966,17'd1559,17'd19499,17'd1138,17'd35772,17'd2786,17'd31732,17'd48292,17'd28549,17'd48293,17'd48294,17'd48295,17'd17674,17'd14880,17'd48296,17'd47272,17'd48077,17'd47273,17'd19006,17'd18774,17'd17206,17'd18657,17'd48297,17'd29049,17'd19893,17'd12361,17'd14764,17'd12813,17'd13093,17'd12530,17'd12218,17'd14890,17'd21184,17'd13598,17'd17096,17'd17204,17'd18657,17'd24012,17'd15008,17'd33548,17'd16029,17'd48080,17'd48080,17'd48298,17'd34178,17'd47972,17'd48299,17'd48300,17'd48301,17'd9704,17'd9007,17'd9159,17'd6468,17'd6626,17'd11089,17'd6138,17'd8692,17'd48302,17'd48303,17'd48304,17'd48305,17'd47872,17'd48306,17'd45668,17'd42354,17'd40124,17'd48307,17'd48308,17'd48309,17'd8708,17'd47978,17'd48310,17'd48311,17'd48196,17'd48312,17'd48313,17'd47984,17'd48314,17'd46374,17'd46503,17'd48315,17'd46808,17'd42808,17'd48316,17'd8252,17'd9483,17'd8878,17'd14674,17'd11135,17'd12423,17'd13368,17'd47782,17'd47884,17'd36626,17'd24706,17'd30229,17'd24208,17'd28111,17'd29928,17'd33572,17'd48317,17'd48318,17'd48319,17'd35801,17'd24540,17'd24029,17'd48204,17'd11129,17'd11962,17'd11806,17'd11960,17'd14807,17'd20452,17'd26629,17'd31768,17'd31941,17'd32283,17'd30834,17'd31761,17'd31763,17'd39211,17'd31587,17'd29067,17'd28943,17'd25672,17'd24992,17'd23167,17'd37196,17'd28352,17'd10330,17'd9740,17'd16319,17'd10742,17'd9479,17'd16554,17'd9470,17'd48320,17'd48321,17'd48322,17'd48323,17'd48324,17'd48325,17'd41934,17'd16555,17'd15181,17'd48326,17'd48327,17'd13654,17'd48328,17'd48329,17'd48330,17'd47607,17'd48111,17'd47791,17'd41513,17'd48331,17'd41513,17'd48332,17'd47897,17'd48222,17'd48333,17'd48334,17'd48335,17'd48336,17'd48337,17'd48338,17'd48339,17'd48340,17'd48341,17'd48342,17'd48232,17'd48127,17'd48343,17'd48344,17'd48235,17'd38774,17'd48345,17'd38778,17'd47127,17'd33451,17'd48239,17'd48239,17'd41852,17'd48241,17'd40198,17'd34074,17'd33766,17'd36238,17'd42865,17'd46313,17'd33915,17'd40502,17'd36249,17'd36523,17'd36523,17'd47035,17'd36523,17'd36523,17'd46931,17'd36378,17'd33916,17'd36969,17'd37235,17'd35274,17'd34076,17'd35407,17'd35273,17'd36247,17'd33620,17'd35273,17'd36246,17'd36385,17'd38391,17'd47807,17'd45736,17'd48346,17'd48347,17'd47809,17'd37635,17'd47038,17'd48348,17'd48349,17'd48350,17'd48351,17'd48352,17'd48353,17'd47638,17'd47436,17'd46840,17'd48157,17'd44822,17'd45873,17'd43154,17'd43019,17'd42301,17'd42301,17'd33310,17'd44231,17'd43695,17'd37778,17'd44359,17'd43836,17'd43835,17'd43550,17'd39591,17'd25180,17'd24252,17'd24086,17'd23566,17'd32191,17'd32008,17'd32351,17'd37117,17'd29687,17'd29688,17'd25031,17'd34284,17'd43835,17'd43018,17'd44589,17'd46202,17'd47445,17'd48354,17'd48265,17'd48355,17'd45879,17'd45987,17'd48356,17'd41265,17'd48357,17'd48358,17'd43689,17'd44102,17'd33308,17'd31353,17'd38537,17'd28726,17'd33963,17'd26782,17'd28725,17'd25707,17'd25566,17'd28369,17'd27637,17'd24897,17'd24744,17'd24898,17'd25178,17'd27882,17'd27766,17'd26530,17'd26901,17'd28726,17'd27642,17'd38537,17'd29379,17'd31503,17'd28134,17'd32355,17'd33321,17'd28134,17'd41731,17'd43433,17'd47822,17'd46759,17'd48260,17'd47534,17'd48047,17'd48359,17'd48360,17'd48361,17'd48362,17'd48363,17'd48263,17'd48264,17'd47936,17'd48364,17'd47932,17'd40826,17'd32016,17'd33963,17'd28482,17'd28594,17'd25179,17'd30275,17'd22679,17'd38041,17'd48365,17'd48366,17'd48277,17'd45766,17'd22511,17'd32498,17'd33480,17'd48367,17'd48368,17'd47356,17'd48272,17'd48369,17'd30276,17'd22332,17'd44368,17'd48367,17'd22325,17'd22674,17'd48370,17'd21850,17'd41728,17'd41866,17'd46116,17'd22337,17'd23222,17'd33945,17'd48371,17'd45887,17'd48372,17'd48373,17'd48374,17'd47846,17'd25069,17'd23092,17'd29737,17'd7823,17'd6384,17'd5332,17'd48173,17'd24484,17'd11854,17'd16615,17'd40394,17'd48375,17'd12761,17'd14301,17'd29296,17'd29296,17'd6391,17'd28185,17'd25627,17'd5002,17'd4683,17'd5144,17'd33367,17'd4188,17'd38442,17'd42910,17'd4841,17'd4841,17'd4995,17'd5153,17'd4841,17'd5002,17'd5004,17'd25627,17'd4687,17'd4188,17'd4831,17'd4829,17'd36165,17'd37147,17'd4825,17'd47959,17'd48376,17'd48177,17'd4510,17'd4668,17'd48377,17'd39471,17'd48286,17'd48378,17'd48379,17'd48380,17'd48287,17'd48381,17'd48382,17'd48288,17'd48383,17'd48074,17'd48384,17'd46698,17'd5772,17'd48385,17'd41002,17'd39789,17'd10388,17'd10388,17'd47767,17'd39181,17'd39483,17'd39033,17'd38580,17'd38580,17'd38072,17'd13420,17'd16492,17'd16492,17'd6258,17'd8186,17'd5776,17'd5776,17'd5958,17'd4882,17'd4713,17'd5940,17'd14178,17'd2098,17'd15233,17'd15233,17'd2589,17'd1272,17'd24165,17'd1407,17'd969,17'd965
},
'{
17'd4428,17'd4892,17'd4733,17'd4246,17'd14188,17'd2422,17'd1967,17'd4247,17'd22965,17'd3905,17'd980,17'd980,17'd980,17'd27,17'd286,17'd27,17'd18,17'd18,17'd289,17'd30,17'd1129,17'd292,17'd33,17'd656,17'd2939,17'd13303,17'd2121,17'd2121,17'd1282,17'd19499,17'd1138,17'd35772,17'd2786,17'd31732,17'd48292,17'd27829,17'd37449,17'd5531,17'd48386,17'd17674,17'd18879,17'd30203,17'd30204,17'd46359,17'd47273,17'd19128,17'd19007,17'd21185,17'd17445,17'd17690,17'd19385,17'd19893,17'd12361,17'd14764,17'd13093,17'd13093,17'd13840,17'd12218,17'd12955,17'd13209,17'd13598,17'd13093,17'd11362,17'd29049,17'd24192,17'd15008,17'd31918,17'd31918,17'd48298,17'd48080,17'd48298,17'd34357,17'd48387,17'd48299,17'd48300,17'd48301,17'd9704,17'd9007,17'd9159,17'd6468,17'd6626,17'd11089,17'd6138,17'd8692,17'd48302,17'd48303,17'd48304,17'd48305,17'd47872,17'd48388,17'd48389,17'd48390,17'd47388,17'd48307,17'd48308,17'd48391,17'd48392,17'd48087,17'd48393,17'd28931,17'd48394,17'd48395,17'd48396,17'd48397,17'd47778,17'd48398,17'd46045,17'd48399,17'd48400,17'd48401,17'd48402,17'd18203,17'd8248,17'd8725,17'd24361,17'd14383,17'd20312,17'd28821,17'd47782,17'd47884,17'd48203,17'd48201,17'd27985,17'd24208,17'd28111,17'd29928,17'd47008,17'd47884,17'd37983,17'd31292,17'd24540,17'd24540,17'd24029,17'd48204,17'd20451,17'd11807,17'd11806,17'd13761,17'd12580,17'd19407,17'd23511,17'd28462,17'd31765,17'd31287,17'd31941,17'd30834,17'd31763,17'd31763,17'd31439,17'd31440,17'd30071,17'd28816,17'd24538,17'd21363,17'd22817,17'd13521,17'd19280,17'd9883,17'd9740,17'd27003,17'd10742,17'd17011,17'd9470,17'd48205,17'd21983,17'd9342,17'd48403,17'd48404,17'd48405,17'd32776,17'd27743,17'd48406,17'd48407,17'd48408,17'd8109,17'd48409,17'd48410,17'd48411,17'd48412,17'd48216,17'd48413,17'd48414,17'd48415,17'd48416,17'd48218,17'd48112,17'd48417,17'd48418,17'd48419,17'd48420,17'd48421,17'd48422,17'd48423,17'd48424,17'd48425,17'd48426,17'd48427,17'd43135,17'd48428,17'd48429,17'd48430,17'd48431,17'd45974,17'd48432,17'd48433,17'd48434,17'd46928,17'd33451,17'd48239,17'd41852,17'd48241,17'd48242,17'd33617,17'd40198,17'd34074,17'd48435,17'd45471,17'd40033,17'd33618,17'd40502,17'd36249,17'd36249,17'd45860,17'd45860,17'd47221,17'd36523,17'd46931,17'd36378,17'd35678,17'd38787,17'd33769,17'd38787,17'd33769,17'd35274,17'd35274,17'd35274,17'd33620,17'd35273,17'd38645,17'd36384,17'd45736,17'd48436,17'd48135,17'd45361,17'd37636,17'd47038,17'd48437,17'd48438,17'd38011,17'd48439,17'd48440,17'd48441,17'd48442,17'd47339,17'd48443,17'd46759,17'd48444,17'd45482,17'd44823,17'd41270,17'd43020,17'd33310,17'd33310,17'd44231,17'd43837,17'd47629,17'd43550,17'd33157,17'd43977,17'd43694,17'd44229,17'd29101,17'd25030,17'd24415,17'd23732,17'd23386,17'd32191,17'd32008,17'd23217,17'd36987,17'd30275,17'd34621,17'd24898,17'd27637,17'd42597,17'd42299,17'd48445,17'd46555,17'd46956,17'd48446,17'd48447,17'd48147,17'd47938,17'd48448,17'd41579,17'd48449,17'd48450,17'd42295,17'd43283,17'd44356,17'd32184,17'd31352,17'd28726,17'd28726,17'd26782,17'd28725,17'd28724,17'd26174,17'd28594,17'd25709,17'd28254,17'd24897,17'd24744,17'd24898,17'd25178,17'd25567,17'd25833,17'd43290,17'd29245,17'd37513,17'd31503,17'd28980,17'd27642,17'd27885,17'd32017,17'd32507,17'd33321,17'd32832,17'd34877,17'd44234,17'd48266,17'd46759,17'd48260,17'd47638,17'd48451,17'd45478,17'd48262,17'd48361,17'd45261,17'd48263,17'd48263,17'd48264,17'd47936,17'd46104,17'd46660,17'd33942,17'd30735,17'd33963,17'd28482,17'd27638,17'd29976,17'd30275,17'd39131,17'd38041,17'd48365,17'd47750,17'd48452,17'd48453,17'd22510,17'd23041,17'd31834,17'd44944,17'd34483,17'd47454,17'd48272,17'd48454,17'd22681,17'd22677,17'd35037,17'd48455,17'd22504,17'd23574,17'd35153,17'd21849,17'd33646,17'd34879,17'd48456,17'd48457,17'd35153,17'd33945,17'd23743,17'd48458,17'd48459,17'd48460,17'd48461,17'd48462,17'd19685,17'd48463,17'd24303,17'd7824,17'd6384,17'd6389,17'd25226,17'd12760,17'd29161,17'd16615,17'd40246,17'd48375,17'd16615,17'd12467,17'd29296,17'd29296,17'd6391,17'd31717,17'd31553,17'd5002,17'd4683,17'd5144,17'd33367,17'd4997,17'd30486,17'd42910,17'd4841,17'd4841,17'd4995,17'd5153,17'd4841,17'd5002,17'd5004,17'd25627,17'd4687,17'd4997,17'd4356,17'd4829,17'd5475,17'd35602,17'd48177,17'd48068,17'd48464,17'd4666,17'd4826,17'd48465,17'd48466,17'd42033,17'd4194,17'd48467,17'd39614,17'd48380,17'd46876,17'd48381,17'd48468,17'd48469,17'd48470,17'd48471,17'd3053,17'd46698,17'd4863,17'd48385,17'd41002,17'd39947,17'd10388,17'd10388,17'd39482,17'd39181,17'd38859,17'd39033,17'd38580,17'd44019,17'd38072,17'd13420,17'd16492,17'd16492,17'd6095,17'd7365,17'd5776,17'd5776,17'd4882,17'd4882,17'd4713,17'd4882,17'd5940,17'd14178,17'd15233,17'd413,17'd598,17'd1272,17'd1963,17'd268,17'd2255,17'd965
},
'{
17'd6420,17'd6420,17'd2935,17'd2935,17'd14188,17'd1688,17'd17187,17'd2257,17'd22965,17'd3905,17'd980,17'd980,17'd980,17'd27,17'd7061,17'd27,17'd18,17'd18,17'd289,17'd30,17'd1129,17'd982,17'd32,17'd656,17'd294,17'd13303,17'd2121,17'd1839,17'd1559,17'd1559,17'd1424,17'd2268,17'd3598,17'd2609,17'd32254,17'd27829,17'd48472,17'd42649,17'd48386,17'd17433,17'd18402,17'd24516,17'd30204,17'd48473,17'd47273,17'd19382,17'd18655,17'd17206,17'd18657,17'd18657,17'd20149,17'd19893,17'd12361,17'd14764,17'd13093,17'd13093,17'd12530,17'd13094,17'd13093,17'd13209,17'd13462,17'd13599,17'd12681,17'd20425,17'd24192,17'd15008,17'd31918,17'd31918,17'd32260,17'd32260,17'd34178,17'd34357,17'd33857,17'd47866,17'd48474,17'd13842,17'd9704,17'd12534,17'd9006,17'd8369,17'd6468,17'd6626,17'd6139,17'd8692,17'd6938,17'd46999,17'd40732,17'd42507,17'd44283,17'd48388,17'd48389,17'd43207,17'd46900,17'd48475,17'd48308,17'd48391,17'd48476,17'd30821,17'd48477,17'd48478,17'd48479,17'd28332,17'd48480,17'd48481,17'd48397,17'd48482,17'd46145,17'd48483,17'd48484,17'd47590,17'd48485,17'd14136,17'd8249,17'd8572,17'd17480,17'd14383,17'd20312,17'd28821,17'd37339,17'd48486,17'd48203,17'd24858,17'd24362,17'd28111,17'd28111,17'd28109,17'd36348,17'd47884,17'd48487,17'd12584,17'd48488,17'd24540,17'd11397,17'd48204,17'd14522,17'd11520,17'd12861,17'd13761,17'd12580,17'd17348,17'd12255,17'd28229,17'd30972,17'd30973,17'd34957,17'd33567,17'd32437,17'd31763,17'd31773,17'd30221,17'd29067,17'd28943,17'd27483,17'd23170,17'd23169,17'd22816,17'd28352,17'd10326,17'd10023,17'd10856,17'd9885,17'd17011,17'd27003,17'd48489,17'd17840,17'd9347,17'd9474,17'd48490,17'd48491,17'd40602,17'd26374,17'd29068,17'd48492,17'd10340,17'd48493,17'd48494,17'd48495,17'd48496,17'd48497,17'd48498,17'd48111,17'd48414,17'd48416,17'd48499,17'd48331,17'd48112,17'd48417,17'd48500,17'd48117,17'd48501,17'd48502,17'd48503,17'd48504,17'd48505,17'd48506,17'd48507,17'd48508,17'd48509,17'd43408,17'd47318,17'd48510,17'd48510,17'd46927,17'd47029,17'd45859,17'd45859,17'd45859,17'd48511,17'd33451,17'd41852,17'd33914,17'd40661,17'd40661,17'd48242,17'd40198,17'd34074,17'd36238,17'd46313,17'd40033,17'd33618,17'd40502,17'd36099,17'd33618,17'd33618,17'd47033,17'd47221,17'd38644,17'd36378,17'd35678,17'd34994,17'd34994,17'd33916,17'd36969,17'd37101,17'd33769,17'd37235,17'd35274,17'd33620,17'd35971,17'd36244,17'd48512,17'd48513,17'd48514,17'd36513,17'd48134,17'd48515,17'd48516,17'd48517,17'd48518,17'd48519,17'd48520,17'd48521,17'd48522,17'd48523,17'd48524,17'd46661,17'd48525,17'd43975,17'd43016,17'd42599,17'd44231,17'd33792,17'd31351,17'd35012,17'd28366,17'd47727,17'd44229,17'd43694,17'd43977,17'd43694,17'd43836,17'd31034,17'd24745,17'd23917,17'd23565,17'd29374,17'd32008,17'd32008,17'd38976,17'd29826,17'd32186,17'd30126,17'd34283,17'd44105,17'd48526,17'd48526,17'd46102,17'd47051,17'd48527,17'd47446,17'd48528,17'd48529,17'd48265,17'd47537,17'd48155,17'd48530,17'd40508,17'd48531,17'd41413,17'd44938,17'd32185,17'd31352,17'd28726,17'd26781,17'd26782,17'd28725,17'd27515,17'd28602,17'd25567,17'd25568,17'd24898,17'd24744,17'd24744,17'd24897,17'd25568,17'd28130,17'd28724,17'd26781,17'd29977,17'd33319,17'd26276,17'd25555,17'd26276,17'd28133,17'd30587,17'd29380,17'd33321,17'd28258,17'd38975,17'd44357,17'd48532,17'd48533,17'd48260,17'd47638,17'd48152,17'd48534,17'd48535,17'd48362,17'd45261,17'd48536,17'd48154,17'd47737,17'd47936,17'd48537,17'd46553,17'd33942,17'd30735,17'd35023,17'd26530,17'd27638,17'd25180,17'd23565,17'd30129,17'd36984,17'd32499,17'd22867,17'd48538,17'd48539,17'd21695,17'd23222,17'd22681,17'd44702,17'd44489,17'd43717,17'd48540,17'd34279,17'd22333,17'd32344,17'd35037,17'd48455,17'd48541,17'd48542,17'd30880,17'd22011,17'd32828,17'd48543,17'd48544,17'd23041,17'd22683,17'd46099,17'd47840,17'd48545,17'd48546,17'd41880,17'd48547,17'd22372,17'd25758,17'd21919,17'd24641,17'd7824,17'd6384,17'd6218,17'd25226,17'd12760,17'd29161,17'd16615,17'd35893,17'd48375,17'd12906,17'd12760,17'd29296,17'd25361,17'd6391,17'd30638,17'd5004,17'd5005,17'd4683,17'd5144,17'd33367,17'd4188,17'd5144,17'd42910,17'd4841,17'd4841,17'd4995,17'd5153,17'd4841,17'd5002,17'd5004,17'd25627,17'd5157,17'd33838,17'd4831,17'd4829,17'd5475,17'd35602,17'd34495,17'd34327,17'd48548,17'd48549,17'd48178,17'd48550,17'd42631,17'd42033,17'd4195,17'd48286,17'd48070,17'd48551,17'd46876,17'd48552,17'd48553,17'd48554,17'd48555,17'd47669,17'd48556,17'd48557,17'd7849,17'd48558,17'd41315,17'd39947,17'd48559,17'd10388,17'd39482,17'd39181,17'd38859,17'd39033,17'd38580,17'd44019,17'd13420,17'd13420,17'd16492,17'd6095,17'd7365,17'd7365,17'd9123,17'd16382,17'd5940,17'd5940,17'd4423,17'd6415,17'd2393,17'd14178,17'd1383,17'd413,17'd423,17'd1685,17'd803,17'd268,17'd2255,17'd2420
},
'{
17'd6420,17'd6420,17'd2935,17'd2935,17'd14070,17'd1688,17'd17187,17'd2257,17'd1416,17'd3905,17'd980,17'd980,17'd27,17'd286,17'd7061,17'd286,17'd18,17'd3905,17'd289,17'd30,17'd1129,17'd292,17'd33,17'd656,17'd294,17'd471,17'd2261,17'd2121,17'd1557,17'd1559,17'd1424,17'd2268,17'd3598,17'd2435,17'd32254,17'd31106,17'd3609,17'd48560,17'd48561,17'd46701,17'd16273,17'd45188,17'd48562,17'd25801,17'd45190,17'd19892,17'd27461,17'd21185,17'd17320,17'd17445,17'd19008,17'd23155,17'd12361,17'd14764,17'd13093,17'd13093,17'd12530,17'd12955,17'd13209,17'd13209,17'd13462,17'd13599,17'd12532,17'd20425,17'd16411,17'd14893,17'd31918,17'd31918,17'd32260,17'd32260,17'd34357,17'd48563,17'd33857,17'd47866,17'd14625,17'd13842,17'd9704,17'd10430,17'd12219,17'd6468,17'd6626,17'd6305,17'd6138,17'd6137,17'd7259,17'd46999,17'd40732,17'd48564,17'd43607,17'd44864,17'd48565,17'd45668,17'd45669,17'd48475,17'd48308,17'd48566,17'd48086,17'd48567,17'd29054,17'd28805,17'd48568,17'd48569,17'd48480,17'd48480,17'd48395,17'd48570,17'd48571,17'd48572,17'd43759,17'd48573,17'd42520,17'd48574,17'd8251,17'd11404,17'd15684,17'd19531,17'd20312,17'd28821,17'd37339,17'd48575,17'd48202,17'd33572,17'd29928,17'd30229,17'd28111,17'd29928,17'd33572,17'd48486,17'd47402,17'd11525,17'd48319,17'd48576,17'd12583,17'd29789,17'd14522,17'd11807,17'd11961,17'd13882,17'd12110,17'd17348,17'd24032,17'd28103,17'd31587,17'd30973,17'd34957,17'd33719,17'd31762,17'd32437,17'd36490,17'd34704,17'd31587,17'd30370,17'd32759,17'd24031,17'd33084,17'd30532,17'd13521,17'd19282,17'd10165,17'd17719,17'd9741,17'd9740,17'd9611,17'd48577,17'd21984,17'd8873,17'd23165,17'd9618,17'd48578,17'd40603,17'd17720,17'd48579,17'd48580,17'd8580,17'd48581,17'd48582,17'd48583,17'd48584,17'd48585,17'd48586,17'd48587,17'd48218,17'd48588,17'd48589,17'd48590,17'd48591,17'd48592,17'd48417,17'd48593,17'd48594,17'd48119,17'd48595,17'd48596,17'd48597,17'd48598,17'd48599,17'd48600,17'd48601,17'd47705,17'd48602,17'd47319,17'd46522,17'd40501,17'd47425,17'd47425,17'd48603,17'd47030,17'd48511,17'd46928,17'd38518,17'd48239,17'd48239,17'd41852,17'd40661,17'd48242,17'd33617,17'd47522,17'd48435,17'd45471,17'd46313,17'd33618,17'd33618,17'd47912,17'd33618,17'd45860,17'd36249,17'd47221,17'd36523,17'd44465,17'd46931,17'd42581,17'd42581,17'd35678,17'd35678,17'd33916,17'd36969,17'd33769,17'd35834,17'd36385,17'd35972,17'd46644,17'd46645,17'd48604,17'd37635,17'd48605,17'd48606,17'd48607,17'd41571,17'd48608,17'd48250,17'd46545,17'd48609,17'd48610,17'd46840,17'd48611,17'd46839,17'd48035,17'd42883,17'd42886,17'd43019,17'd33478,17'd28252,17'd25833,17'd25565,17'd28253,17'd43978,17'd43022,17'd43836,17'd29825,17'd43836,17'd43977,17'd29244,17'd24742,17'd23917,17'd29242,17'd29374,17'd29974,17'd23215,17'd37117,17'd29099,17'd34883,17'd24416,17'd29976,17'd48612,17'd48145,17'd48613,17'd48614,17'd44355,17'd48615,17'd47343,17'd46761,17'd48616,17'd43542,17'd45607,17'd48617,17'd48618,17'd48619,17'd42877,17'd47931,17'd42436,17'd35011,17'd31352,17'd26901,17'd26782,17'd28725,17'd26903,17'd25949,17'd30606,17'd28597,17'd27512,17'd24898,17'd24745,17'd24417,17'd24897,17'd25177,17'd28720,17'd31827,17'd28979,17'd32354,17'd28134,17'd27761,17'd26780,17'd26276,17'd28133,17'd29380,17'd31196,17'd32017,17'd39743,17'd38805,17'd43701,17'd48532,17'd48620,17'd48144,17'd47638,17'd48621,17'd46199,17'd48535,17'd48361,17'd48622,17'd48536,17'd48154,17'd47737,17'd47936,17'd46762,17'd48623,17'd33477,17'd31035,17'd35023,17'd26530,17'd27638,17'd25030,17'd23565,17'd30129,17'd48624,17'd48625,17'd48626,17'd48627,17'd22338,17'd22004,17'd22861,17'd30276,17'd32015,17'd48628,17'd43717,17'd48540,17'd33945,17'd22160,17'd30427,17'd35037,17'd48455,17'd48629,17'd23039,17'd21848,17'd21695,17'd48630,17'd48631,17'd46849,17'd32829,17'd22160,17'd35292,17'd45373,17'd46336,17'd48632,17'd44127,17'd48547,17'd25209,17'd19468,17'd22734,17'd25624,17'd23799,17'd5481,17'd6218,17'd14048,17'd11854,17'd11710,17'd16615,17'd35759,17'd35478,17'd13046,17'd14049,17'd44613,17'd25361,17'd6220,17'd31891,17'd32553,17'd5005,17'd4683,17'd5144,17'd4188,17'd4997,17'd4996,17'd4995,17'd4841,17'd4841,17'd4995,17'd42910,17'd4841,17'd5002,17'd5004,17'd25627,17'd5157,17'd41891,17'd4356,17'd4670,17'd5475,17'd36438,17'd44381,17'd35188,17'd33530,17'd36302,17'd47372,17'd48633,17'd4185,17'd4356,17'd4195,17'd48634,17'd48635,17'd48551,17'd47476,17'd37812,17'd48636,17'd48637,17'd3373,17'd3556,17'd48638,17'd48639,17'd7849,17'd5493,17'd41315,17'd41315,17'd41003,17'd10388,17'd39482,17'd39790,17'd38859,17'd39033,17'd38580,17'd44019,17'd13420,17'd13176,17'd16492,17'd6095,17'd7365,17'd7365,17'd9123,17'd16382,17'd5940,17'd5630,17'd4423,17'd4423,17'd5940,17'd2393,17'd1383,17'd2589,17'd1408,17'd411,17'd970,17'd2778,17'd211,17'd2420
},
'{
17'd6420,17'd6420,17'd2935,17'd2935,17'd14070,17'd1688,17'd17187,17'd22965,17'd4089,17'd18,17'd27,17'd27,17'd27,17'd286,17'd7385,17'd7061,17'd652,17'd3905,17'd289,17'd30,17'd1129,17'd982,17'd32,17'd656,17'd294,17'd2939,17'd2121,17'd1702,17'd1283,17'd1559,17'd1841,17'd2268,17'd4583,17'd4095,17'd3440,17'd2798,17'd3609,17'd48560,17'd20139,17'd48640,17'd28666,17'd24010,17'd25910,17'd25911,17'd29763,17'd19892,17'd27461,17'd21185,17'd17320,17'd18657,17'd19383,17'd23155,17'd12362,17'd14764,17'd13599,17'd13093,17'd12218,17'd12955,17'd13209,17'd13462,17'd13597,17'd13092,17'd11764,17'd19383,17'd15902,17'd14892,17'd24194,17'd24194,17'd32260,17'd32260,17'd48641,17'd48642,17'd48387,17'd47866,17'd14473,17'd13468,17'd13972,17'd9159,17'd12219,17'd12220,17'd6141,17'd6140,17'd6139,17'd6137,17'd7259,17'd46489,17'd40425,17'd48643,17'd48644,17'd43204,17'd48565,17'd45531,17'd44284,17'd48475,17'd48308,17'd47875,17'd48645,17'd48476,17'd48646,17'd29462,17'd48647,17'd48648,17'd48649,17'd48480,17'd48650,17'd48651,17'd48652,17'd48653,17'd44032,17'd48654,17'd48655,17'd48656,17'd14527,17'd9349,17'd9041,17'd11809,17'd11401,17'd48657,17'd29927,17'd48486,17'd48203,17'd23167,17'd24995,17'd30229,17'd28111,17'd27860,17'd45684,17'd35799,17'd28688,17'd29335,17'd36072,17'd14382,17'd18327,17'd22816,17'd31137,17'd13762,17'd11961,17'd13761,17'd12110,17'd12580,17'd19407,17'd28107,17'd30373,17'd31941,17'd33719,17'd48658,17'd32438,17'd32438,17'd48659,17'd48660,17'd31439,17'd29330,17'd29923,17'd26371,17'd24539,17'd24994,17'd38499,17'd11669,17'd19532,17'd10166,17'd9883,17'd9740,17'd46267,17'd19918,17'd24039,17'd9044,17'd19415,17'd28569,17'd9737,17'd40603,17'd10741,17'd15681,17'd48661,17'd32121,17'd48662,17'd48663,17'd48664,17'd48665,17'd48666,17'd48667,17'd48668,17'd48669,17'd48591,17'd48670,17'd48671,17'd48670,17'd48500,17'd48500,17'd48593,17'd48672,17'd46814,17'd48330,17'd48673,17'd48674,17'd48675,17'd48676,17'd48677,17'd48678,17'd48679,17'd48680,17'd48681,17'd35125,17'd48682,17'd48683,17'd48684,17'd46532,17'd45730,17'd48685,17'd47030,17'd48511,17'd38518,17'd33451,17'd48239,17'd33914,17'd40661,17'd40661,17'd48241,17'd47522,17'd33766,17'd36238,17'd46313,17'd46313,17'd40033,17'd33618,17'd40502,17'd36099,17'd36099,17'd40502,17'd47033,17'd45860,17'd36249,17'd36249,17'd47035,17'd38644,17'd44465,17'd33916,17'd36969,17'd35407,17'd36246,17'd38787,17'd48686,17'd47715,17'd48687,17'd48688,17'd46541,17'd48689,17'd48690,17'd48691,17'd48692,17'd48031,17'd45478,17'd46762,17'd43832,17'd46843,17'd48693,17'd48694,17'd46546,17'd43154,17'd42886,17'd42599,17'd32995,17'd25833,17'd27766,17'd25708,17'd25566,17'd33157,17'd38156,17'd38156,17'd39443,17'd43157,17'd43553,17'd29976,17'd24743,17'd28722,17'd29826,17'd23388,17'd29974,17'd23217,17'd32191,17'd31029,17'd34883,17'd24895,17'd48695,17'd48696,17'd48697,17'd48698,17'd46435,17'd44099,17'd48699,17'd48700,17'd47054,17'd48701,17'd46439,17'd48702,17'd48703,17'd48704,17'd42293,17'd42592,17'd48705,17'd39741,17'd30735,17'd29245,17'd27027,17'd28725,17'd28725,17'd27514,17'd28481,17'd28598,17'd28717,17'd25178,17'd25030,17'd24895,17'd24742,17'd24745,17'd25438,17'd32658,17'd32343,17'd29245,17'd28373,17'd32017,17'd27884,17'd26523,17'd27761,17'd28257,17'd31196,17'd31196,17'd32355,17'd35854,17'd40824,17'd43701,17'd48532,17'd48620,17'd48706,17'd47732,17'd48707,17'd46199,17'd48535,17'd48361,17'd48622,17'd48708,17'd48154,17'd47641,17'd48709,17'd45479,17'd48710,17'd27372,17'd26901,17'd35304,17'd28482,17'd25567,17'd24895,17'd34137,17'd23740,17'd31829,17'd32499,17'd48626,17'd22337,17'd22338,17'd22004,17'd48711,17'd30276,17'd32015,17'd48628,17'd43854,17'd48712,17'd23394,17'd22159,17'd37510,17'd44368,17'd48455,17'd48713,17'd48714,17'd48715,17'd48716,17'd35295,17'd48717,17'd45882,17'd33480,17'd22682,17'd22683,17'd38173,17'd48718,17'd48719,17'd48720,17'd47368,17'd48721,17'd19468,17'd48722,17'd48723,17'd23975,17'd5611,17'd5615,17'd14048,17'd14049,17'd11710,17'd16615,17'd48375,17'd35478,17'd12905,17'd11853,17'd44613,17'd25361,17'd6220,17'd30333,17'd30637,17'd5005,17'd4683,17'd5144,17'd4188,17'd4991,17'd5144,17'd4995,17'd5328,17'd4841,17'd4995,17'd42910,17'd4841,17'd5002,17'd5004,17'd25627,17'd5157,17'd33838,17'd45393,17'd4670,17'd5475,17'd45284,17'd35190,17'd36882,17'd5140,17'd4353,17'd48465,17'd48377,17'd41455,17'd4017,17'd48724,17'd48725,17'd48378,17'd48551,17'd48726,17'd48727,17'd48728,17'd48729,17'd48730,17'd48731,17'd48732,17'd48733,17'd7849,17'd4056,17'd41315,17'd41315,17'd41159,17'd39180,17'd10906,17'd39790,17'd38859,17'd39033,17'd38580,17'd44019,17'd44387,17'd16492,17'd6095,17'd6095,17'd7365,17'd5776,17'd16256,17'd16382,17'd5940,17'd5630,17'd4423,17'd4423,17'd5940,17'd2393,17'd413,17'd598,17'd204,17'd1685,17'd206,17'd257,17'd965,17'd182
},
'{
17'd6420,17'd6420,17'd2935,17'd2935,17'd14070,17'd1688,17'd17187,17'd22965,17'd4089,17'd18,17'd27,17'd27,17'd27,17'd286,17'd7555,17'd285,17'd980,17'd3905,17'd289,17'd30,17'd1129,17'd982,17'd32,17'd656,17'd294,17'd2939,17'd1972,17'd1972,17'd1557,17'd1559,17'd1841,17'd2268,17'd2786,17'd3917,17'd3268,17'd2798,17'd2625,17'd48560,17'd42198,17'd14757,17'd18526,17'd24341,17'd48734,17'd25911,17'd29763,17'd19128,17'd27461,17'd21650,17'd17320,17'd17207,17'd18656,17'd17317,17'd12362,17'd14764,17'd12954,17'd13599,17'd12955,17'd13093,17'd13209,17'd13462,17'd13597,17'd35352,17'd11764,17'd46245,17'd16034,17'd14768,17'd15008,17'd24194,17'd16029,17'd32260,17'd48641,17'd48735,17'd48298,17'd31743,17'd14475,17'd13721,17'd9300,17'd8537,17'd12219,17'd44629,17'd6140,17'd6305,17'd6138,17'd8692,17'd7259,17'd46489,17'd40425,17'd48736,17'd48644,17'd43204,17'd45079,17'd45531,17'd44284,17'd48475,17'd7113,17'd48737,17'd48391,17'd48738,17'd29910,17'd48393,17'd48739,17'd48740,17'd48741,17'd48742,17'd28332,17'd48743,17'd46374,17'd45678,17'd48744,17'd47104,17'd48745,17'd34694,17'd17730,17'd17126,17'd15297,17'd17232,17'd37735,17'd20046,17'd48657,17'd48486,17'd36626,17'd33572,17'd24539,17'd24362,17'd28111,17'd27985,17'd48201,17'd35799,17'd17842,17'd42674,17'd43622,17'd45207,17'd12583,17'd22816,17'd48746,17'd13762,17'd11960,17'd13761,17'd12109,17'd12580,17'd17348,17'd23681,17'd28572,17'd30972,17'd32283,17'd48658,17'd48747,17'd32438,17'd48659,17'd48660,17'd30834,17'd31440,17'd30831,17'd29327,17'd24031,17'd25143,17'd37196,17'd21206,17'd28352,17'd24996,17'd11134,17'd17719,17'd20044,17'd27003,17'd9192,17'd19033,17'd24039,17'd24037,17'd25675,17'd10023,17'd48748,17'd25530,17'd48749,17'd48750,17'd10610,17'd22481,17'd48751,17'd48752,17'd48753,17'd48754,17'd47412,17'd48006,17'd48755,17'd48670,17'd48756,17'd48757,17'd48758,17'd48759,17'd48222,17'd44774,17'd48117,17'd48760,17'd48761,17'd48762,17'd48763,17'd48764,17'd48765,17'd48766,17'd48767,17'd48679,17'd48768,17'd48769,17'd48770,17'd48771,17'd48772,17'd48773,17'd48774,17'd48511,17'd45859,17'd48511,17'd38518,17'd33451,17'd41852,17'd33914,17'd33914,17'd48775,17'd47031,17'd47522,17'd33766,17'd48435,17'd36238,17'd36238,17'd36238,17'd42865,17'd42865,17'd40033,17'd33915,17'd40502,17'd47033,17'd33915,17'd40033,17'd42865,17'd40033,17'd36099,17'd47035,17'd42135,17'd34994,17'd35274,17'd35274,17'd33618,17'd45731,17'd45733,17'd48688,17'd48776,17'd48777,17'd48778,17'd48779,17'd48780,17'd46544,17'd47330,17'd48781,17'd45744,17'd44697,17'd48782,17'd31648,17'd48783,17'd44823,17'd42599,17'd40825,17'd43288,17'd25707,17'd27766,17'd26064,17'd28723,17'd25435,17'd32996,17'd42749,17'd43977,17'd29101,17'd38282,17'd38406,17'd25032,17'd24415,17'd23564,17'd29830,17'd30579,17'd29974,17'd37117,17'd29530,17'd33801,17'd23916,17'd32007,17'd48784,17'd48145,17'd46327,17'd48785,17'd46758,17'd43831,17'd48786,17'd48700,17'd48787,17'd48701,17'd43420,17'd48787,17'd48788,17'd48789,17'd40814,17'd40512,17'd40822,17'd36690,17'd28727,17'd29245,17'd30586,17'd28725,17'd26903,17'd25949,17'd27638,17'd33000,17'd28717,17'd25178,17'd25180,17'd25032,17'd24417,17'd24897,17'd25709,17'd25565,17'd36542,17'd27642,17'd32355,17'd32355,17'd27884,17'd26652,17'd28370,17'd28372,17'd29106,17'd29106,17'd32505,17'd41429,17'd42740,17'd44822,17'd48790,17'd48791,17'd48706,17'd47444,17'd48792,17'd48360,17'd48362,17'd48361,17'd48264,17'd48793,17'd48154,17'd47737,17'd48709,17'd45479,17'd44228,17'd27146,17'd26781,17'd33499,17'd28482,17'd25567,17'd24898,17'd34137,17'd41419,17'd48794,17'd32347,17'd47939,17'd22337,17'd35156,17'd41865,17'd22162,17'd22331,17'd32015,17'd33645,17'd43854,17'd34905,17'd39745,17'd22161,17'd32660,17'd33944,17'd39441,17'd22334,17'd48795,17'd22009,17'd48796,17'd23044,17'd48797,17'd44716,17'd39441,17'd22860,17'd32666,17'd48798,17'd48799,17'd48800,17'd48801,17'd47368,17'd48802,17'd20237,17'd47957,17'd27079,17'd23975,17'd4844,17'd6219,17'd14049,17'd11853,17'd11710,17'd12906,17'd36735,17'd41142,17'd11710,17'd11576,17'd44613,17'd25361,17'd5919,17'd30333,17'd30180,17'd5005,17'd4683,17'd5144,17'd4997,17'd38442,17'd5145,17'd4995,17'd5328,17'd4841,17'd5327,17'd5152,17'd4841,17'd5329,17'd5004,17'd25627,17'd5157,17'd41891,17'd4017,17'd42630,17'd4828,17'd35748,17'd35190,17'd35190,17'd36301,17'd33990,17'd4827,17'd42628,17'd33208,17'd4186,17'd48803,17'd48724,17'd39315,17'd48804,17'd48805,17'd48727,17'd48806,17'd48807,17'd48808,17'd48731,17'd48809,17'd48810,17'd7849,17'd40411,17'd48811,17'd48812,17'd41159,17'd41160,17'd10906,17'd39790,17'd38859,17'd39033,17'd38580,17'd44019,17'd44387,17'd16492,17'd6095,17'd6095,17'd7365,17'd5776,17'd9123,17'd5940,17'd5940,17'd5630,17'd4713,17'd4713,17'd5940,17'd2393,17'd14178,17'd598,17'd1537,17'd1111,17'd207,17'd1242,17'd1682,17'd182
},
'{
17'd4892,17'd6420,17'd2935,17'd2422,17'd10535,17'd1688,17'd1415,17'd17,17'd4089,17'd3905,17'd27,17'd27,17'd26,17'd285,17'd1832,17'd285,17'd27,17'd652,17'd289,17'd290,17'd291,17'd982,17'd32,17'd33,17'd2260,17'd13303,17'd22615,17'd1702,17'd1558,17'd1559,17'd1841,17'd2434,17'd3917,17'd33851,17'd3268,17'd48813,17'd48814,17'd5395,17'd48815,17'd44620,17'd48816,17'd14758,17'd48817,17'd48818,17'd29763,17'd19128,17'd19007,17'd21185,17'd17320,17'd17207,17'd17205,17'd17317,17'd12361,17'd14621,17'd13599,17'd13210,17'd13599,17'd13209,17'd14469,17'd14469,17'd12678,17'd35352,17'd13969,17'd19620,17'd48297,17'd14219,17'd17811,17'd32101,17'd15384,17'd48387,17'd48819,17'd48820,17'd48821,17'd47866,17'd14347,17'd16880,17'd15517,17'd10694,17'd8369,17'd6468,17'd6467,17'd10695,17'd6304,17'd8073,17'd7259,17'd39647,17'd48822,17'd40120,17'd48823,17'd43607,17'd48824,17'd48825,17'd44760,17'd48826,17'd48827,17'd7113,17'd48828,17'd48829,17'd48830,17'd48831,17'd48832,17'd48833,17'd48834,17'd48835,17'd48836,17'd48837,17'd48838,17'd47881,17'd48839,17'd48840,17'd48841,17'd48842,17'd46378,17'd48843,17'd20176,17'd12117,17'd11276,17'd19919,17'd34205,17'd39069,17'd36626,17'd47008,17'd47886,17'd26372,17'd26496,17'd27985,17'd24706,17'd18327,17'd17966,17'd48844,17'd12423,17'd48845,17'd13254,17'd22816,17'd48746,17'd11964,17'd13761,17'd12109,17'd12418,17'd13517,17'd48846,17'd26755,17'd26758,17'd28825,17'd31588,17'd32592,17'd48847,17'd48847,17'd38498,17'd33568,17'd34381,17'd31439,17'd31764,17'd47107,17'd27483,17'd21363,17'd11396,17'd10854,17'd11669,17'd28352,17'd19532,17'd10023,17'd46267,17'd16319,17'd15180,17'd9044,17'd38496,17'd48848,17'd15048,17'd11670,17'd27236,17'd10023,17'd48849,17'd47406,17'd7786,17'd17852,17'd48850,17'd48851,17'd48852,17'd48853,17'd48854,17'd48855,17'd45816,17'd48856,17'd48499,17'd48857,17'd48858,17'd48859,17'd48860,17'd48333,17'd48861,17'd48862,17'd48863,17'd48864,17'd48865,17'd48866,17'd48867,17'd48868,17'd48869,17'd48870,17'd48871,17'd48872,17'd48873,17'd46630,17'd48874,17'd48875,17'd48876,17'd48877,17'd33763,17'd33763,17'd46520,17'd48878,17'd48879,17'd48880,17'd48774,17'd48774,17'd33616,17'd47031,17'd39115,17'd48881,17'd35263,17'd35263,17'd35397,17'd45596,17'd36238,17'd36238,17'd35542,17'd35542,17'd46640,17'd33766,17'd33766,17'd48882,17'd48883,17'd34421,17'd48884,17'd34591,17'd48885,17'd46744,17'd48886,17'd46830,17'd48887,17'd43411,17'd37367,17'd45029,17'd48247,17'd48888,17'd48889,17'd48890,17'd48891,17'd48892,17'd48893,17'd47930,17'd48894,17'd46556,17'd48157,17'd48525,17'd42883,17'd43019,17'd40826,17'd33310,17'd33642,17'd28602,17'd28600,17'd28600,17'd29970,17'd43550,17'd25435,17'd27765,17'd25317,17'd41730,17'd32668,17'd32659,17'd23731,17'd28976,17'd29374,17'd30579,17'd29374,17'd29531,17'd29241,17'd30424,17'd34883,17'd48895,17'd48526,17'd48896,17'd48897,17'd48898,17'd47237,17'd48899,17'd48900,17'd47936,17'd46847,17'd48901,17'd46105,17'd48902,17'd48903,17'd48904,17'd47828,17'd48905,17'd43298,17'd27642,17'd29246,17'd28980,17'd27027,17'd28853,17'd26903,17'd30734,17'd28369,17'd28719,17'd27512,17'd25320,17'd30432,17'd25180,17'd24897,17'd28974,17'd32669,17'd28978,17'd30577,17'd26276,17'd28257,17'd28371,17'd28133,17'd26897,17'd28372,17'd28857,17'd33166,17'd29249,17'd28258,17'd37114,17'd43700,17'd48444,17'd48906,17'd48907,17'd47933,17'd48908,17'd46321,17'd48360,17'd48361,17'd48264,17'd48362,17'd48793,17'd48363,17'd48909,17'd48910,17'd42296,17'd44104,17'd27027,17'd27027,17'd27515,17'd26064,17'd27882,17'd25032,17'd29242,17'd35158,17'd34455,17'd32499,17'd35855,17'd22511,17'd23044,17'd45876,17'd32350,17'd44591,17'd44702,17'd40523,17'd46958,17'd30728,17'd32503,17'd48911,17'd22158,17'd32344,17'd22333,17'd30728,17'd32829,17'd21695,17'd32347,17'd22510,17'd48912,17'd23393,17'd32190,17'd48913,17'd48914,17'd48915,17'd48916,17'd48917,17'd48918,17'd48919,17'd48920,17'd48921,17'd24299,17'd27080,17'd5326,17'd5331,17'd8303,17'd30332,17'd10642,17'd11710,17'd13046,17'd30488,17'd30488,17'd11577,17'd10514,17'd44613,17'd6392,17'd28185,17'd5004,17'd5004,17'd5005,17'd4526,17'd4999,17'd33992,17'd41891,17'd5145,17'd4683,17'd4686,17'd4686,17'd28536,17'd31552,17'd4842,17'd25627,17'd5004,17'd25627,17'd5157,17'd41891,17'd33533,17'd42772,17'd4828,17'd43455,17'd35602,17'd37147,17'd35748,17'd35889,17'd46013,17'd42772,17'd33208,17'd5477,17'd4366,17'd48922,17'd39316,17'd48923,17'd48924,17'd36448,17'd48925,17'd48926,17'd48927,17'd48731,17'd3865,17'd45785,17'd7849,17'd4056,17'd40411,17'd3709,17'd41160,17'd4554,17'd10906,17'd38458,17'd38334,17'd41481,17'd38072,17'd38072,17'd37959,17'd37959,17'd6095,17'd6095,17'd7365,17'd9123,17'd3073,17'd3073,17'd5940,17'd4729,17'd5630,17'd5776,17'd16382,17'd12496,17'd2393,17'd11337,17'd1111,17'd803,17'd262,17'd801,17'd1682,17'd592
},
'{
17'd4892,17'd4428,17'd2593,17'd2784,17'd3252,17'd1688,17'd17187,17'd17,17'd4089,17'd3905,17'd27,17'd27,17'd26,17'd285,17'd1832,17'd285,17'd980,17'd652,17'd289,17'd30,17'd1129,17'd982,17'd32,17'd33,17'd2260,17'd13303,17'd2121,17'd1972,17'd1701,17'd1559,17'd1841,17'd2434,17'd3917,17'd33851,17'd3268,17'd48813,17'd48814,17'd5395,17'd48928,17'd44620,17'd48929,17'd18163,17'd47088,17'd48818,17'd29763,17'd19128,17'd19007,17'd36756,17'd27833,17'd19008,17'd18774,17'd11629,17'd11913,17'd12218,17'd13093,17'd13210,17'd32570,17'd13463,17'd16284,17'd14469,17'd15516,17'd35352,17'd12361,17'd48930,17'd47863,17'd14219,17'd17811,17'd14893,17'd14474,17'd48387,17'd48931,17'd48932,17'd48821,17'd47972,17'd14347,17'd15766,17'd15517,17'd10694,17'd6468,17'd6468,17'd6467,17'd10695,17'd6304,17'd8073,17'd6938,17'd47187,17'd48303,17'd40583,17'd42063,17'd48305,17'd48824,17'd48825,17'd44760,17'd48933,17'd48934,17'd48935,17'd48936,17'd48829,17'd48937,17'd48938,17'd48939,17'd48940,17'd48941,17'd48835,17'd48942,17'd9326,17'd47778,17'd46374,17'd48943,17'd48944,17'd43901,17'd47398,17'd48945,17'd8098,17'd8727,17'd8874,17'd14383,17'd19919,17'd34205,17'd18326,17'd36626,17'd47008,17'd47886,17'd36346,17'd26495,17'd29928,17'd21361,17'd18327,17'd29790,17'd47402,17'd11525,17'd24364,17'd13254,17'd11668,17'd29789,17'd18444,17'd11960,17'd12109,17'd12418,17'd14003,17'd34558,17'd13515,17'd16685,17'd27858,17'd31129,17'd31287,17'd33088,17'd48946,17'd48947,17'd38498,17'd48660,17'd34704,17'd31763,17'd36777,17'd29778,17'd23170,17'd17478,17'd11808,17'd28463,17'd11669,17'd28352,17'd10165,17'd9740,17'd9619,17'd15187,17'd8720,17'd17237,17'd16441,17'd15566,17'd11670,17'd27739,17'd10023,17'd48849,17'd48948,17'd19780,17'd25154,17'd48949,17'd48950,17'd48951,17'd48952,17'd48953,17'd48954,17'd48011,17'd48955,17'd48757,17'd48956,17'd48957,17'd48958,17'd48959,17'd48759,17'd48861,17'd48960,17'd48961,17'd48962,17'd48963,17'd48964,17'd48965,17'd48966,17'd48967,17'd48968,17'd48969,17'd48970,17'd48971,17'd40032,17'd33913,17'd42134,17'd48972,17'd43961,17'd38780,17'd48973,17'd46398,17'd38771,17'd48974,17'd38771,17'd48975,17'd48603,17'd33616,17'd33616,17'd48241,17'd48976,17'd44464,17'd48977,17'd46632,17'd46632,17'd48242,17'd48242,17'd47031,17'd46929,17'd46929,17'd46929,17'd47522,17'd34420,17'd33767,17'd48978,17'd35399,17'd34733,17'd48979,17'd45731,17'd48980,17'd46536,17'd46746,17'd43534,17'd42868,17'd44924,17'd48981,17'd48982,17'd48983,17'd48984,17'd48985,17'd46945,17'd41861,17'd44355,17'd48782,17'd48986,17'd48444,17'd45610,17'd46425,17'd41111,17'd40826,17'd43551,17'd25565,17'd28594,17'd28130,17'd29970,17'd28484,17'd44229,17'd28600,17'd27765,17'd28369,17'd29103,17'd38808,17'd30431,17'd23732,17'd23386,17'd23923,17'd23387,17'd48257,17'd23385,17'd32186,17'd29534,17'd48987,17'd48988,17'd48896,17'd46553,17'd47932,17'd46756,17'd48522,17'd40669,17'd48788,17'd47446,17'd46558,17'd43542,17'd43420,17'd48989,17'd48788,17'd47736,17'd47054,17'd48990,17'd39740,17'd33952,17'd37513,17'd28980,17'd27027,17'd28724,17'd26174,17'd28599,17'd29244,17'd24897,17'd27637,17'd25177,17'd29244,17'd29976,17'd24897,17'd27764,17'd38671,17'd27027,17'd27368,17'd27884,17'd28371,17'd28372,17'd29247,17'd28855,17'd28857,17'd29690,17'd48991,17'd29249,17'd32831,17'd41274,17'd43844,17'd48157,17'd48992,17'd48533,17'd48045,17'd48993,17'd48049,17'd48361,17'd45261,17'd48622,17'd48362,17'd48994,17'd48995,17'd43541,17'd47053,17'd43422,17'd42883,17'd27027,17'd27258,17'd27514,17'd28594,17'd27882,17'd24898,17'd29242,17'd35158,17'd34455,17'd32499,17'd35855,17'd22511,17'd35156,17'd48996,17'd23926,17'd32190,17'd23391,17'd23926,17'd46958,17'd23393,17'd36289,17'd48911,17'd36289,17'd32344,17'd22333,17'd30728,17'd45755,17'd48717,17'd48631,17'd48457,17'd31344,17'd34107,17'd44591,17'd48913,17'd44939,17'd48997,17'd48998,17'd48999,17'd48918,17'd49000,17'd48920,17'd22915,17'd24301,17'd10043,17'd5326,17'd5158,17'd8303,17'd10514,17'd10642,17'd11710,17'd13046,17'd49001,17'd49001,17'd11577,17'd30487,17'd35475,17'd6221,17'd5335,17'd5004,17'd5002,17'd5005,17'd4684,17'd41459,17'd41891,17'd41891,17'd5145,17'd4683,17'd4841,17'd4841,17'd28536,17'd31401,17'd30180,17'd25627,17'd5004,17'd25627,17'd4848,17'd34657,17'd39468,17'd4185,17'd40848,17'd5475,17'd45394,17'd45284,17'd36165,17'd46228,17'd43046,17'd4185,17'd5604,17'd4990,17'd4362,17'd4021,17'd39169,17'd49002,17'd49003,17'd49004,17'd49005,17'd49006,17'd49007,17'd3558,17'd48733,17'd8786,17'd7849,17'd5493,17'd40411,17'd3709,17'd41160,17'd18383,17'd11048,17'd38458,17'd38334,17'd41481,17'd38072,17'd38072,17'd37959,17'd37959,17'd6095,17'd6095,17'd7365,17'd9123,17'd3073,17'd2097,17'd4882,17'd4729,17'd49008,17'd49009,17'd16382,17'd12496,17'd2409,17'd604,17'd1111,17'd641,17'd1097,17'd610,17'd212,17'd40102
},
'{
17'd4243,17'd25384,17'd2935,17'd2422,17'd1831,17'd1127,17'd16,17'd16,17'd4089,17'd18,17'd27,17'd27,17'd26,17'd285,17'd1832,17'd285,17'd980,17'd652,17'd289,17'd468,17'd290,17'd291,17'd2259,17'd32,17'd2262,17'd13303,17'd2121,17'd1702,17'd1558,17'd1283,17'd1704,17'd2434,17'd3917,17'd3603,17'd30949,17'd49010,17'd49011,17'd21337,17'd49012,17'd24970,17'd49013,17'd14609,17'd27216,17'd48818,17'd29763,17'd19128,17'd19007,17'd27461,17'd19255,17'd19008,17'd18774,17'd12531,17'd12530,17'd14890,17'd13599,17'd13599,17'd32570,17'd13463,17'd14469,17'd14469,17'd11625,17'd35352,17'd12362,17'd32102,17'd47863,17'd15902,17'd17208,17'd17691,17'd14768,17'd47866,17'd48931,17'd48932,17'd48821,17'd47866,17'd49014,17'd10565,17'd9574,17'd10428,17'd8369,17'd6468,17'd7417,17'd6466,17'd9008,17'd8074,17'd39646,17'd47187,17'd49015,17'd40583,17'd48736,17'd49016,17'd43608,17'd49017,17'd44633,17'd48933,17'd48475,17'd49018,17'd49019,17'd31933,17'd49020,17'd49021,17'd49022,17'd49023,17'd49024,17'd49025,17'd49026,17'd27226,17'd47984,17'd48398,17'd49027,17'd49028,17'd49029,17'd49030,17'd43218,17'd49031,17'd8408,17'd8720,17'd16549,17'd12585,17'd11525,17'd36072,17'd44772,17'd36348,17'd33084,17'd24993,17'd29928,17'd29928,17'd24363,17'd17478,17'd22991,17'd48487,17'd11525,17'd33714,17'd13254,17'd11808,17'd48101,17'd18082,17'd11958,17'd12109,17'd12859,17'd12418,17'd13515,17'd13515,17'd18564,17'd25528,17'd31285,17'd32283,17'd49032,17'd49033,17'd48947,17'd38498,17'd48660,17'd34381,17'd30834,17'd30072,17'd29923,17'd24538,17'd23167,17'd11397,17'd11668,17'd21206,17'd28352,17'd19532,17'd10023,17'd25673,17'd10742,17'd8874,17'd9348,17'd8720,17'd18556,17'd12585,17'd10165,17'd10023,17'd15681,17'd49034,17'd49035,17'd48003,17'd49036,17'd49037,17'd49038,17'd48665,17'd49039,17'd49040,17'd49041,17'd49042,17'd49043,17'd49044,17'd49045,17'd49046,17'd49047,17'd49048,17'd49049,17'd44534,17'd49050,17'd49051,17'd49052,17'd49053,17'd49054,17'd49055,17'd49056,17'd49057,17'd49058,17'd49059,17'd49060,17'd47708,17'd35125,17'd49061,17'd49062,17'd49063,17'd49064,17'd49065,17'd48877,17'd47030,17'd34419,17'd41092,17'd41092,17'd34419,17'd33914,17'd41852,17'd41852,17'd46829,17'd46742,17'd48132,17'd40661,17'd33914,17'd49066,17'd46415,17'd33451,17'd48239,17'd49067,17'd47323,17'd40198,17'd33766,17'd36238,17'd34730,17'd47032,17'd44465,17'd38519,17'd48132,17'd49068,17'd49069,17'd48512,17'd49070,17'd49071,17'd49072,17'd38266,17'd49073,17'd49074,17'd49075,17'd49076,17'd49077,17'd49078,17'd49079,17'd46556,17'd48897,17'd46546,17'd42741,17'd43019,17'd43288,17'd42437,17'd32995,17'd28602,17'd27638,17'd27765,17'd25317,17'd28484,17'd42749,17'd28484,17'd25317,17'd29103,17'd29976,17'd30733,17'd24087,17'd34137,17'd23386,17'd29530,17'd23388,17'd29975,17'd23918,17'd33652,17'd34883,17'd49080,17'd49081,17'd48897,17'd46553,17'd48986,17'd47051,17'd43015,17'd42144,17'd48704,17'd49082,17'd48701,17'd45262,17'd46847,17'd49083,17'd49084,17'd47538,17'd46666,17'd49085,17'd32184,17'd29379,17'd37513,17'd28980,17'd27027,17'd26903,17'd26064,17'd33000,17'd27637,17'd28595,17'd27637,17'd29244,17'd30432,17'd29976,17'd28974,17'd28480,17'd27767,17'd33163,17'd49086,17'd28256,17'd29537,17'd29380,17'd28257,17'd29104,17'd29536,17'd29979,17'd48991,17'd29249,17'd39438,17'd39275,17'd43974,17'd44226,17'd49087,17'd49088,17'd48151,17'd47445,17'd49089,17'd49090,17'd48622,17'd48622,17'd49091,17'd49092,17'd49093,17'd43541,17'd48910,17'd45035,17'd43016,17'd26902,17'd28853,17'd27514,17'd28594,17'd25438,17'd24745,17'd28976,17'd35158,17'd31347,17'd32347,17'd35855,17'd22511,17'd33798,17'd38172,17'd39441,17'd40523,17'd48913,17'd23926,17'd32503,17'd32503,17'd32661,17'd49094,17'd22158,17'd22674,17'd22333,17'd33480,17'd46670,17'd49095,17'd48631,17'd32498,17'd49096,17'd40523,17'd44591,17'd39281,17'd44121,17'd49097,17'd49098,17'd49099,17'd48720,17'd49100,17'd49101,17'd49102,17'd22082,17'd27305,17'd5479,17'd5158,17'd8303,17'd10514,17'd10642,17'd11710,17'd12905,17'd49001,17'd11709,17'd13678,17'd30487,17'd25361,17'd26828,17'd5160,17'd5004,17'd5005,17'd4686,17'd5156,17'd41459,17'd41891,17'd33841,17'd5145,17'd4839,17'd4840,17'd4841,17'd28536,17'd31552,17'd30180,17'd25627,17'd5004,17'd5329,17'd34921,17'd5154,17'd33691,17'd41612,17'd4829,17'd5475,17'd35748,17'd35748,17'd4669,17'd4828,17'd5476,17'd4831,17'd33041,17'd5754,17'd4190,17'd4673,17'd49103,17'd49104,17'd49105,17'd49106,17'd49005,17'd3371,17'd49107,17'd49108,17'd48733,17'd4863,17'd7849,17'd4056,17'd48812,17'd39179,17'd4554,17'd4865,17'd5026,17'd38458,17'd38334,17'd41481,17'd38072,17'd13420,17'd37959,17'd37959,17'd6095,17'd7365,17'd5776,17'd9123,17'd5940,17'd5940,17'd4713,17'd4729,17'd49008,17'd49009,17'd12496,17'd12026,17'd2409,17'd192,17'd1396,17'd271,17'd408,17'd460,17'd639,17'd40102
},
'{
17'd4243,17'd4892,17'd2593,17'd2422,17'd1831,17'd1127,17'd16,17'd17,17'd4089,17'd18,17'd27,17'd27,17'd26,17'd285,17'd1832,17'd285,17'd980,17'd652,17'd289,17'd30,17'd1129,17'd982,17'd292,17'd33,17'd2260,17'd2939,17'd2121,17'd1972,17'd1701,17'd1283,17'd1704,17'd2268,17'd3917,17'd33851,17'd3268,17'd48813,17'd48814,17'd5672,17'd49109,17'd49110,17'd49111,17'd18648,17'd47088,17'd48818,17'd29763,17'd19128,17'd19007,17'd27461,17'd19255,17'd19008,17'd17689,17'd10815,17'd12956,17'd12065,17'd13093,17'd13599,17'd13463,17'd13598,17'd14469,17'd14469,17'd11625,17'd35352,17'd12362,17'd32102,17'd18657,17'd15524,17'd17208,17'd17811,17'd14346,17'd47866,17'd48931,17'd48932,17'd48821,17'd48299,17'd49014,17'd15766,17'd15517,17'd9159,17'd6468,17'd6468,17'd7417,17'd7085,17'd6304,17'd8073,17'd49112,17'd47187,17'd49015,17'd40426,17'd48736,17'd42507,17'd43608,17'd49017,17'd44633,17'd49113,17'd49114,17'd38356,17'd49115,17'd49116,17'd49117,17'd48830,17'd48310,17'd49118,17'd49119,17'd49120,17'd49121,17'd49122,17'd48397,17'd49123,17'd46145,17'd49124,17'd49125,17'd49126,17'd49127,17'd49128,17'd19535,17'd9621,17'd17232,17'd17479,17'd20046,17'd31292,17'd23337,17'd14382,17'd24858,17'd26258,17'd24539,17'd24539,17'd24363,17'd14382,17'd23166,17'd48487,17'd13647,17'd16687,17'd11523,17'd25280,17'd29789,17'd30980,17'd13883,17'd12109,17'd12859,17'd12859,17'd14003,17'd13515,17'd12108,17'd23511,17'd31768,17'd30834,17'd33875,17'd49033,17'd48947,17'd49129,17'd48660,17'd34835,17'd30973,17'd31439,17'd30071,17'd27004,17'd21363,17'd18327,17'd11398,17'd11399,17'd11669,17'd19532,17'd10741,17'd9739,17'd9741,17'd9344,17'd8873,17'd9044,17'd26875,17'd37735,17'd11670,17'd9883,17'd26759,17'd47298,17'd47599,17'd49130,17'd49131,17'd49132,17'd49133,17'd49134,17'd49135,17'd49136,17'd49137,17'd49138,17'd48117,17'd49139,17'd49047,17'd49140,17'd49045,17'd49140,17'd49141,17'd44036,17'd49142,17'd39217,17'd49143,17'd49144,17'd49145,17'd49146,17'd49147,17'd49148,17'd49149,17'd49150,17'd49151,17'd37089,17'd42580,17'd47319,17'd49152,17'd49153,17'd49154,17'd49155,17'd49156,17'd38779,17'd48345,17'd47802,17'd49157,17'd49158,17'd47616,17'd38771,17'd46534,17'd46534,17'd38770,17'd38770,17'd46928,17'd46928,17'd47616,17'd49159,17'd48511,17'd38518,17'd48775,17'd47322,17'd48242,17'd40198,17'd33766,17'd46313,17'd45860,17'd38644,17'd45596,17'd49160,17'd49161,17'd49162,17'd33621,17'd49163,17'd48247,17'd49164,17'd49165,17'd49166,17'd49167,17'd49168,17'd49169,17'd49170,17'd49078,17'd43546,17'd46201,17'd45745,17'd42436,17'd41271,17'd43288,17'd42437,17'd42147,17'd28253,17'd28723,17'd28130,17'd25567,17'd28717,17'd29970,17'd42749,17'd39591,17'd31034,17'd29976,17'd30126,17'd35159,17'd24086,17'd29242,17'd29827,17'd29530,17'd29374,17'd23386,17'd29528,17'd34883,17'd34106,17'd49171,17'd48785,17'd48897,17'd46327,17'd47635,17'd39582,17'd49172,17'd42144,17'd49173,17'd49082,17'd49174,17'd47735,17'd47446,17'd49175,17'd48994,17'd47936,17'd49176,17'd49177,17'd33942,17'd29379,17'd37513,17'd28979,17'd28853,17'd26174,17'd28598,17'd25709,17'd24898,17'd34622,17'd28254,17'd29244,17'd25178,17'd27637,17'd28485,17'd28717,17'd26062,17'd30735,17'd49178,17'd49179,17'd36848,17'd31196,17'd28372,17'd29380,17'd36848,17'd36132,17'd48991,17'd29249,17'd45613,17'd39584,17'd43692,17'd39903,17'd49180,17'd49181,17'd47637,17'd45607,17'd48262,17'd49182,17'd49183,17'd45261,17'd48264,17'd49092,17'd49184,17'd48622,17'd46955,17'd45035,17'd43154,17'd26902,17'd28853,17'd27514,17'd28720,17'd25438,17'd24744,17'd28976,17'd35158,17'd31347,17'd32347,17'd33161,17'd22338,17'd33796,17'd49094,17'd39281,17'd40523,17'd39441,17'd30728,17'd32503,17'd36427,17'd31031,17'd49094,17'd32503,17'd22506,17'd22333,17'd32666,17'd49185,17'd48631,17'd49186,17'd31660,17'd22008,17'd32190,17'd44591,17'd35157,17'd38420,17'd46450,17'd49187,17'd49188,17'd43863,17'd49189,17'd24628,17'd26705,17'd25622,17'd27305,17'd5479,17'd5612,17'd8303,17'd28184,17'd10642,17'd29161,17'd11710,17'd49001,17'd11709,17'd30332,17'd28058,17'd35194,17'd26949,17'd25627,17'd5004,17'd5005,17'd4842,17'd4684,17'd41459,17'd41891,17'd33841,17'd6067,17'd4995,17'd4841,17'd4841,17'd28536,17'd31716,17'd30180,17'd25627,17'd5004,17'd5329,17'd34921,17'd5154,17'd33691,17'd41612,17'd4829,17'd4669,17'd36165,17'd5475,17'd40848,17'd5476,17'd4185,17'd4017,17'd5477,17'd4359,17'd4517,17'd49190,17'd39019,17'd49191,17'd49192,17'd49193,17'd21154,17'd49194,17'd49195,17'd49108,17'd48639,17'd4863,17'd7849,17'd4056,17'd49196,17'd41159,17'd39180,17'd10906,17'd11048,17'd11867,17'd38334,17'd41481,17'd38072,17'd13420,17'd37959,17'd37959,17'd6095,17'd7365,17'd5776,17'd5776,17'd5940,17'd5940,17'd4713,17'd4729,17'd49008,17'd49009,17'd12496,17'd12026,17'd6868,17'd192,17'd1396,17'd207,17'd40563,17'd403,17'd592,17'd591
},
'{
17'd4243,17'd25384,17'd2935,17'd2422,17'd1831,17'd1127,17'd16,17'd17,17'd4089,17'd18,17'd27,17'd27,17'd285,17'd285,17'd285,17'd285,17'd980,17'd652,17'd289,17'd468,17'd3433,17'd3254,17'd982,17'd32,17'd2262,17'd2939,17'd2121,17'd1702,17'd1558,17'd1558,17'd1704,17'd2268,17'd1978,17'd33851,17'd3268,17'd49010,17'd49011,17'd21337,17'd49012,17'd49110,17'd49197,17'd47768,17'd27600,17'd49198,17'd45190,17'd19382,17'd17689,17'd19007,17'd19255,17'd18656,17'd17941,17'd11913,17'd12218,17'd12955,17'd13599,17'd13599,17'd13463,17'd13462,17'd14763,17'd14763,17'd11762,17'd35352,17'd12218,17'd32261,17'd20425,17'd24348,17'd17575,17'd17811,17'd14346,17'd15641,17'd49199,17'd48820,17'd49200,17'd48299,17'd14220,17'd10429,17'd9702,17'd9574,17'd8369,17'd6468,17'd6141,17'd7085,17'd49201,17'd8847,17'd7423,17'd49202,17'd49203,17'd40425,17'd48736,17'd42507,17'd42938,17'd48824,17'd46899,17'd49113,17'd49204,17'd49205,17'd49206,17'd49207,17'd49208,17'd29767,17'd49209,17'd49210,17'd49211,17'd48941,17'd49212,17'd49213,17'd48313,17'd49214,17'd49215,17'd49216,17'd44032,17'd49217,17'd49127,17'd49218,17'd8245,17'd8881,17'd10173,17'd17718,17'd19919,17'd16687,17'd25280,17'd11396,17'd23167,17'd24706,17'd24993,17'd29488,17'd14259,17'd14382,17'd35799,17'd49219,17'd36349,17'd28821,17'd11523,17'd11523,17'd22816,17'd49220,17'd11806,17'd12110,17'd12256,17'd12859,17'd14003,17'd13515,17'd14003,17'd49221,17'd28572,17'd29785,17'd33875,17'd34545,17'd49222,17'd48947,17'd33568,17'd34203,17'd31128,17'd31765,17'd31940,17'd28816,17'd24992,17'd16442,17'd11397,17'd11398,17'd11669,17'd11400,17'd10326,17'd11134,17'd9884,17'd11809,17'd10174,17'd15682,17'd10172,17'd27490,17'd11135,17'd11671,17'd16070,17'd28578,17'd33238,17'd49223,17'd49224,17'd49225,17'd49226,17'd49227,17'd48964,17'd47789,17'd49228,17'd49229,17'd49230,17'd45816,17'd49049,17'd49231,17'd49232,17'd49233,17'd49234,17'd42521,17'd49235,17'd49236,17'd49237,17'd49238,17'd49239,17'd49240,17'd49241,17'd49242,17'd49243,17'd49244,17'd49245,17'd49246,17'd49247,17'd49248,17'd49249,17'd49250,17'd47420,17'd49251,17'd46529,17'd49252,17'd49253,17'd49254,17'd49255,17'd49256,17'd49257,17'd47321,17'd49258,17'd49259,17'd48771,17'd48682,17'd48973,17'd38775,17'd33763,17'd33763,17'd34419,17'd49260,17'd48239,17'd41852,17'd33616,17'd47323,17'd46640,17'd35542,17'd49261,17'd33765,17'd46828,17'd35396,17'd49262,17'd49263,17'd37638,17'd49264,17'd49265,17'd49266,17'd49267,17'd49268,17'd49269,17'd49270,17'd49271,17'd49272,17'd47930,17'd40364,17'd48613,17'd43975,17'd44827,17'd41111,17'd33155,17'd43695,17'd49273,17'd28721,17'd28600,17'd27765,17'd33000,17'd31856,17'd42749,17'd43977,17'd41730,17'd32353,17'd30126,17'd23916,17'd30431,17'd23732,17'd29242,17'd23566,17'd23387,17'd29374,17'd31502,17'd29527,17'd34883,17'd49080,17'd49274,17'd49275,17'd46437,17'd46433,17'd40364,17'd44588,17'd49276,17'd42144,17'd49277,17'd49278,17'd48700,17'd49279,17'd49280,17'd49281,17'd48994,17'd48446,17'd49282,17'd49283,17'd36542,17'd29379,17'd37513,17'd28979,17'd28725,17'd28602,17'd28597,17'd25178,17'd24744,17'd23562,17'd25030,17'd25320,17'd28254,17'd25029,17'd28485,17'd28597,17'd27514,17'd31352,17'd49284,17'd49285,17'd36848,17'd31196,17'd28857,17'd28728,17'd49286,17'd36132,17'd48991,17'd29249,17'd35990,17'd40366,17'd44362,17'd44937,17'd49180,17'd48144,17'd49287,17'd48049,17'd45261,17'd49288,17'd49289,17'd49090,17'd43281,17'd49092,17'd49184,17'd48264,17'd41267,17'd49078,17'd41418,17'd27027,17'd28853,17'd27514,17'd28720,17'd27511,17'd24744,17'd28976,17'd35158,17'd48624,17'd34110,17'd32663,17'd22510,17'd23041,17'd36427,17'd48913,17'd40523,17'd23926,17'd23393,17'd32666,17'd49094,17'd38172,17'd33649,17'd22683,17'd49290,17'd22160,17'd32013,17'd48797,17'd48625,17'd32011,17'd21848,17'd46099,17'd30276,17'd48913,17'd39745,17'd49291,17'd49292,17'd49293,17'd38176,17'd43035,17'd46010,17'd24630,17'd21450,17'd22083,17'd7989,17'd5609,17'd5158,17'd8154,17'd28184,17'd10642,17'd29161,17'd29161,17'd49294,17'd11431,17'd10514,17'd6555,17'd6392,17'd5335,17'd5004,17'd5004,17'd5005,17'd4686,17'd5156,17'd41459,17'd41891,17'd33841,17'd6067,17'd4682,17'd4840,17'd4841,17'd28536,17'd31716,17'd30637,17'd25627,17'd5002,17'd5329,17'd5157,17'd33841,17'd33691,17'd41612,17'd42630,17'd4669,17'd4669,17'd35332,17'd4670,17'd42630,17'd4831,17'd4357,17'd4358,17'd4189,17'd49295,17'd4030,17'd49296,17'd49297,17'd49298,17'd49299,17'd49300,17'd49301,17'd49302,17'd48638,17'd41905,17'd42043,17'd3869,17'd3870,17'd49196,17'd41159,17'd10388,17'd39032,17'd38458,17'd11867,17'd38334,17'd38580,17'd38072,17'd13420,17'd37959,17'd37959,17'd6095,17'd7365,17'd5940,17'd5940,17'd4882,17'd4882,17'd4713,17'd4729,17'd8185,17'd5630,17'd5630,17'd8185,17'd11062,17'd411,17'd259,17'd257,17'd2115,17'd17551,17'd40102,17'd40102
},
'{
17'd4243,17'd4892,17'd2593,17'd2422,17'd1831,17'd1127,17'd16,17'd17,17'd4089,17'd18,17'd286,17'd286,17'd285,17'd285,17'd285,17'd286,17'd652,17'd652,17'd289,17'd289,17'd3595,17'd3254,17'd982,17'd32,17'd2262,17'd2939,17'd2121,17'd1972,17'd1701,17'd1558,17'd2267,17'd1706,17'd1978,17'd31732,17'd3603,17'd48813,17'd48814,17'd5672,17'd49109,17'd49110,17'd49197,17'd47768,17'd27600,17'd49198,17'd45406,17'd19382,17'd17689,17'd19007,17'd19255,17'd18656,17'd17941,17'd12680,17'd12218,17'd12955,17'd13599,17'd13599,17'd13598,17'd13597,17'd14763,17'd14763,17'd11762,17'd35352,17'd12218,17'd32261,17'd17572,17'd15899,17'd17692,17'd16987,17'd14219,17'd15641,17'd49303,17'd48820,17'd49200,17'd48299,17'd14220,17'd15898,17'd13471,17'd9574,17'd8369,17'd6468,17'd6141,17'd7085,17'd49201,17'd8847,17'd7423,17'd49202,17'd46895,17'd40425,17'd48736,17'd42507,17'd42938,17'd48824,17'd48825,17'd49304,17'd39969,17'd49305,17'd49306,17'd49307,17'd49308,17'd49309,17'd29054,17'd49310,17'd49311,17'd49312,17'd49313,17'd49212,17'd49314,17'd49315,17'd47685,17'd49316,17'd49317,17'd49318,17'd49319,17'd49320,17'd14135,17'd10027,17'd26153,17'd16561,17'd10331,17'd14134,17'd17236,17'd11396,17'd23513,17'd24858,17'd24993,17'd24993,17'd24706,17'd14382,17'd36072,17'd49321,17'd36349,17'd13368,17'd25280,17'd11523,17'd22816,17'd49322,17'd13883,17'd12109,17'd12859,17'd12859,17'd14003,17'd13515,17'd14003,17'd21504,17'd37206,17'd29482,17'd33568,17'd34545,17'd49033,17'd49222,17'd33720,17'd34203,17'd31127,17'd30973,17'd37065,17'd29066,17'd26493,17'd21363,17'd17478,17'd11274,17'd21206,17'd11525,17'd19282,17'd10326,17'd10329,17'd12116,17'd9345,17'd9190,17'd49323,17'd17606,17'd27490,17'd14928,17'd16070,17'd32916,17'd49324,17'd49325,17'd49326,17'd49327,17'd49328,17'd49329,17'd49330,17'd48753,17'd49331,17'd30556,17'd49332,17'd49333,17'd44410,17'd49231,17'd49232,17'd49334,17'd49335,17'd49336,17'd49337,17'd49338,17'd49339,17'd49340,17'd49341,17'd49342,17'd49343,17'd49344,17'd49345,17'd49346,17'd49347,17'd49348,17'd49349,17'd49350,17'd49351,17'd49352,17'd49353,17'd40347,17'd33615,17'd49354,17'd49355,17'd49356,17'd49357,17'd49358,17'd49359,17'd49360,17'd49361,17'd49362,17'd49363,17'd47908,17'd48130,17'd48432,17'd46530,17'd48973,17'd41092,17'd47616,17'd33451,17'd48239,17'd47322,17'd47323,17'd49364,17'd33764,17'd49365,17'd47425,17'd46740,17'd48024,17'd49366,17'd49367,17'd49368,17'd49369,17'd49370,17'd49371,17'd48351,17'd49372,17'd49373,17'd49374,17'd47234,17'd49375,17'd43691,17'd46756,17'd48526,17'd42886,17'd45878,17'd43551,17'd35012,17'd43837,17'd47438,17'd42749,17'd28369,17'd28717,17'd31520,17'd31366,17'd42749,17'd29825,17'd33483,17'd34276,17'd24249,17'd31033,17'd32186,17'd23918,17'd29376,17'd29376,17'd29686,17'd23386,17'd29241,17'd29375,17'd48987,17'd49376,17'd49377,17'd49377,17'd49378,17'd46665,17'd39582,17'd43284,17'd49379,17'd40669,17'd49380,17'd48446,17'd48155,17'd47538,17'd48536,17'd49381,17'd49382,17'd49383,17'd49384,17'd49385,17'd37908,17'd29379,17'd29246,17'd28979,17'd27515,17'd28594,17'd25709,17'd24898,17'd24743,17'd23562,17'd25030,17'd25320,17'd25029,17'd33951,17'd33951,17'd28594,17'd27259,17'd27642,17'd49179,17'd49285,17'd29831,17'd29106,17'd29536,17'd29536,17'd49286,17'd36132,17'd49386,17'd29249,17'd40677,17'd45612,17'd44362,17'd45157,17'd49387,17'd48151,17'd49388,17'd47937,17'd49183,17'd49389,17'd49390,17'd49182,17'd48263,17'd49391,17'd48708,17'd47737,17'd49392,17'd44225,17'd41270,17'd26902,17'd28853,17'd26530,17'd28723,17'd27511,17'd24417,17'd28976,17'd35158,17'd48624,17'd48796,17'd35295,17'd32498,17'd31345,17'd32503,17'd32190,17'd40523,17'd32350,17'd45986,17'd48911,17'd31193,17'd48624,17'd33649,17'd45986,17'd22334,17'd35292,17'd31344,17'd48544,17'd48625,17'd35156,17'd30880,17'd22334,17'd30276,17'd48913,17'd36717,17'd45756,17'd49393,17'd49394,17'd49395,17'd49396,17'd49397,17'd19687,17'd21606,17'd49398,17'd7989,17'd5610,17'd5331,17'd8154,17'd28184,17'd11037,17'd11577,17'd11577,17'd33209,17'd11181,17'd28184,17'd37031,17'd26828,17'd25627,17'd30637,17'd25627,17'd5005,17'd4686,17'd5156,17'd5154,17'd41891,17'd33841,17'd6067,17'd4995,17'd5328,17'd4841,17'd28536,17'd28536,17'd30637,17'd25627,17'd5002,17'd5329,17'd5157,17'd41891,17'd33691,17'd41612,17'd4830,17'd40848,17'd40848,17'd4670,17'd4830,17'd4016,17'd4017,17'd4515,17'd33991,17'd49295,17'd49399,17'd4199,17'd49400,17'd49401,17'd49402,17'd49403,17'd49404,17'd49405,17'd49406,17'd49407,17'd41905,17'd6081,17'd3869,17'd4394,17'd40099,17'd41159,17'd10388,17'd45186,17'd39181,17'd38859,17'd38860,17'd44019,17'd38072,17'd13420,17'd37959,17'd37959,17'd6095,17'd4869,17'd5630,17'd5940,17'd4882,17'd4882,17'd4713,17'd4729,17'd8185,17'd5630,17'd5630,17'd5372,17'd192,17'd1111,17'd260,17'd1242,17'd211,17'd1095,17'd591,17'd592
},
'{
17'd4243,17'd25384,17'd2935,17'd2422,17'd1831,17'd1127,17'd16,17'd3905,17'd2938,17'd652,17'd286,17'd286,17'd285,17'd467,17'd285,17'd285,17'd980,17'd652,17'd289,17'd289,17'd3595,17'd3254,17'd2940,17'd3253,17'd2262,17'd2939,17'd2121,17'd1839,17'd1422,17'd41008,17'd2267,17'd37171,17'd2786,17'd31732,17'd3603,17'd49408,17'd26739,17'd49409,17'd49410,17'd49411,17'd49412,17'd14330,17'd27600,17'd49198,17'd45406,17'd19006,17'd19893,17'd17689,17'd17206,17'd18656,17'd17204,17'd12680,17'd13094,17'd12955,17'd13209,17'd13209,17'd13462,17'd13597,17'd14344,17'd14344,17'd12062,17'd12677,17'd13211,17'd28554,17'd19891,17'd17319,17'd17448,17'd17575,17'd15902,17'd14473,17'd49303,17'd48820,17'd49200,17'd48299,17'd14220,17'd10429,17'd11088,17'd9574,17'd8369,17'd8369,17'd6625,17'd7085,17'd49201,17'd8847,17'd7423,17'd48302,17'd49413,17'd49414,17'd48304,17'd42507,17'd42938,17'd48824,17'd49017,17'd49304,17'd49415,17'd49305,17'd49416,17'd49417,17'd49418,17'd28443,17'd49419,17'd49420,17'd49421,17'd49422,17'd49423,17'd49424,17'd49026,17'd48837,17'd47684,17'd49425,17'd49426,17'd49427,17'd49428,17'd44874,17'd8243,17'd11403,17'd8874,17'd18556,17'd11671,17'd11400,17'd11524,17'd14673,17'd19158,17'd22472,17'd26258,17'd24993,17'd24706,17'd36348,17'd36072,17'd34205,17'd36349,17'd34205,17'd43622,17'd11523,17'd19533,17'd49220,17'd13135,17'd12419,17'd12256,17'd12997,17'd12418,17'd12417,17'd12417,17'd14003,17'd16556,17'd28572,17'd30677,17'd33875,17'd49033,17'd49033,17'd33720,17'd33568,17'd33568,17'd34835,17'd30834,17'd34551,17'd29778,17'd23515,17'd16325,17'd16068,17'd11524,17'd12423,17'd11132,17'd11133,17'd10166,17'd17719,17'd9479,17'd9340,17'd22812,17'd17232,17'd19279,17'd14383,17'd16070,17'd16070,17'd33722,17'd49429,17'd49430,17'd49431,17'd49432,17'd49433,17'd49434,17'd49241,17'd49435,17'd49436,17'd49437,17'd49438,17'd49439,17'd49339,17'd49231,17'd49440,17'd49046,17'd49335,17'd49441,17'd49336,17'd49442,17'd49443,17'd49444,17'd49445,17'd49446,17'd49447,17'd49448,17'd49449,17'd49450,17'd49451,17'd49452,17'd49453,17'd49454,17'd49455,17'd49456,17'd49456,17'd49457,17'd49458,17'd49459,17'd49460,17'd49458,17'd42423,17'd48770,17'd46739,17'd49061,17'd49061,17'd40805,17'd40805,17'd48236,17'd49461,17'd40501,17'd46530,17'd47520,17'd34419,17'd34419,17'd46928,17'd48775,17'd47323,17'd49462,17'd33765,17'd33616,17'd49463,17'd49464,17'd35543,17'd36112,17'd49465,17'd49466,17'd49467,17'd49468,17'd49469,17'd49268,17'd49470,17'd49471,17'd49472,17'd49473,17'd49375,17'd40957,17'd46555,17'd49474,17'd44590,17'd42437,17'd33642,17'd32658,17'd43978,17'd43550,17'd39591,17'd25438,17'd28480,17'd31520,17'd28597,17'd28484,17'd39591,17'd32668,17'd35159,17'd30275,17'd30275,17'd24087,17'd23918,17'd29376,17'd23387,17'd29374,17'd29376,17'd29528,17'd33652,17'd49475,17'd46202,17'd49377,17'd49377,17'd49476,17'd46954,17'd48610,17'd42295,17'd40956,17'd49477,17'd49380,17'd48446,17'd48153,17'd43281,17'd49478,17'd49479,17'd43147,17'd49480,17'd43692,17'd33791,17'd38025,17'd31352,17'd28727,17'd26901,17'd26174,17'd25567,17'd25320,17'd28718,17'd28975,17'd28852,17'd25180,17'd25320,17'd27764,17'd49481,17'd33484,17'd27766,17'd27027,17'd31354,17'd49482,17'd36848,17'd29831,17'd30884,17'd29979,17'd29978,17'd36132,17'd36132,17'd49386,17'd34285,17'd35150,17'd44361,17'd39583,17'd41862,17'd49387,17'd47339,17'd49483,17'd48363,17'd49484,17'd49485,17'd49485,17'd49486,17'd48708,17'd49391,17'd48536,17'd47737,17'd49392,17'd44355,17'd42599,17'd26902,17'd28725,17'd26530,17'd28602,17'd25709,17'd24252,17'd23386,17'd35017,17'd48794,17'd45265,17'd23044,17'd31660,17'd31658,17'd32350,17'd40523,17'd32190,17'd23393,17'd32013,17'd31497,17'd49487,17'd48624,17'd33649,17'd33480,17'd22159,17'd22507,17'd31660,17'd48631,17'd33161,17'd48457,17'd48370,17'd22682,17'd30276,17'd22505,17'd49488,17'd49489,17'd49490,17'd49491,17'd49492,17'd49493,17'd49494,17'd19469,17'd26948,17'd49495,17'd23975,17'd5482,17'd5332,17'd8154,17'd27815,17'd28057,17'd11316,17'd11316,17'd28305,17'd27932,17'd8780,17'd37031,17'd5762,17'd4842,17'd4842,17'd5329,17'd4845,17'd4686,17'd4840,17'd4996,17'd38442,17'd5144,17'd6067,17'd4682,17'd4683,17'd4841,17'd28418,17'd28536,17'd30637,17'd5160,17'd5002,17'd27570,17'd34656,17'd33841,17'd42180,17'd4017,17'd4016,17'd5476,17'd42630,17'd4671,17'd4831,17'd4017,17'd4515,17'd34157,17'd33838,17'd49496,17'd49497,17'd49498,17'd49499,17'd4205,17'd36037,17'd49500,17'd49501,17'd49502,17'd49503,17'd49504,17'd41480,17'd3869,17'd49505,17'd5494,17'd40099,17'd41159,17'd10388,17'd39032,17'd11048,17'd11867,17'd41481,17'd12913,17'd38072,17'd13420,17'd37959,17'd6095,17'd4713,17'd4713,17'd5630,17'd5630,17'd4713,17'd4882,17'd4713,17'd4729,17'd4729,17'd4713,17'd6415,17'd5371,17'd604,17'd425,17'd3899,17'd256,17'd2255,17'd2420,17'd591,17'd612
},
'{
17'd27713,17'd4243,17'd2593,17'd2422,17'd1831,17'd1127,17'd1277,17'd18,17'd2938,17'd652,17'd286,17'd286,17'd285,17'd467,17'd285,17'd286,17'd652,17'd652,17'd29,17'd289,17'd3595,17'd3254,17'd2940,17'd3253,17'd3103,17'd3103,17'd2600,17'd2121,17'd1702,17'd41008,17'd2267,17'd37171,17'd2786,17'd33542,17'd3603,17'd49506,17'd26981,17'd49507,17'd49508,17'd49411,17'd49412,17'd14330,17'd27600,17'd49509,17'd45406,17'd19006,17'd19893,17'd17689,17'd17206,17'd25512,17'd19006,17'd12680,17'd13094,17'd12955,17'd13209,17'd13209,17'd13968,17'd13597,17'd14344,17'd14344,17'd12062,17'd12677,17'd13211,17'd22630,17'd19891,17'd16289,17'd17448,17'd17810,17'd24348,17'd14473,17'd49303,17'd48820,17'd49200,17'd48299,17'd14220,17'd15898,17'd20426,17'd9702,17'd8369,17'd8369,17'd6625,17'd7085,17'd9985,17'd8847,17'd7423,17'd48302,17'd49413,17'd40271,17'd48304,17'd42507,17'd42938,17'd48824,17'd49017,17'd49304,17'd49415,17'd49510,17'd49511,17'd49512,17'd49418,17'd49513,17'd29461,17'd49514,17'd49515,17'd49516,17'd49517,17'd49518,17'd49519,17'd49520,17'd48093,17'd49521,17'd49522,17'd49523,17'd49524,17'd44408,17'd8243,17'd30671,17'd9189,17'd17717,17'd16561,17'd11670,17'd10476,17'd11274,17'd19158,17'd16442,17'd24706,17'd24993,17'd24858,17'd23513,17'd12583,17'd34205,17'd36349,17'd34205,17'd43622,17'd11523,17'd19533,17'd41343,17'd16325,17'd14130,17'd19032,17'd13884,17'd12859,17'd12418,17'd12417,17'd14003,17'd21504,17'd28348,17'd30073,17'd34203,17'd49525,17'd49033,17'd49032,17'd33720,17'd33568,17'd33568,17'd32283,17'd39211,17'd30830,17'd27347,17'd22992,17'd11521,17'd25280,17'd12584,17'd11399,17'd11132,17'd10166,17'd17719,17'd9741,17'd9620,17'd23679,17'd17232,17'd16549,17'd19279,17'd14928,17'd14928,17'd10479,17'd49526,17'd49527,17'd49528,17'd49529,17'd49530,17'd49531,17'd49448,17'd49532,17'd49533,17'd49534,17'd49332,17'd49535,17'd49536,17'd49537,17'd49538,17'd49539,17'd49540,17'd15680,17'd15805,17'd49541,17'd49542,17'd49543,17'd49544,17'd49545,17'd49546,17'd49547,17'd49548,17'd49549,17'd49550,17'd49551,17'd49552,17'd49553,17'd49554,17'd49555,17'd48768,17'd49556,17'd49557,17'd49558,17'd43678,17'd47907,17'd49559,17'd49559,17'd46522,17'd39411,17'd39411,17'd39411,17'd44919,17'd49560,17'd46927,17'd42284,17'd46529,17'd40501,17'd41565,17'd41565,17'd48973,17'd48876,17'd49067,17'd49561,17'd46929,17'd47519,17'd47124,17'd35543,17'd49562,17'd35973,17'd49563,17'd49564,17'd49565,17'd49566,17'd49567,17'd49568,17'd49569,17'd49570,17'd49571,17'd49572,17'd49375,17'd48523,17'd49275,17'd41583,17'd43838,17'd45749,17'd28483,17'd32658,17'd32996,17'd29970,17'd27511,17'd25177,17'd28480,17'd31520,17'd25567,17'd25317,17'd41730,17'd38808,17'd30431,17'd23384,17'd23565,17'd32186,17'd23918,17'd29376,17'd23923,17'd29374,17'd30127,17'd24087,17'd33482,17'd49171,17'd49378,17'd49275,17'd48898,17'd46756,17'd41106,17'd43423,17'd49379,17'd49573,17'd49574,17'd49380,17'd48709,17'd48262,17'd48363,17'd49575,17'd49479,17'd49576,17'd48147,17'd42600,17'd31352,17'd35570,17'd29245,17'd28727,17'd27027,17'd27766,17'd27882,17'd29976,17'd29100,17'd30275,17'd24902,17'd32007,17'd25177,17'd33803,17'd49577,17'd25567,17'd25707,17'd31035,17'd28258,17'd49578,17'd36132,17'd29979,17'd49579,17'd30131,17'd30280,17'd36132,17'd36132,17'd34286,17'd29107,17'd37248,17'd44361,17'd39583,17'd41862,17'd49387,17'd49580,17'd49581,17'd49184,17'd49582,17'd49583,17'd49583,17'd49584,17'd49585,17'd49391,17'd48708,17'd49586,17'd48899,17'd44821,17'd42599,17'd26902,17'd28725,17'd28482,17'd26064,17'd25709,17'd24252,17'd29826,17'd35017,17'd48794,17'd49587,17'd33798,17'd31346,17'd32502,17'd23926,17'd34107,17'd39281,17'd32503,17'd32829,17'd31344,17'd49487,17'd49588,17'd33649,17'd32502,17'd22683,17'd32829,17'd49589,17'd48625,17'd32499,17'd33162,17'd22683,17'd22681,17'd30276,17'd46454,17'd47840,17'd49590,17'd49591,17'd49592,17'd49593,17'd19302,17'd22901,17'd49594,17'd49595,17'd49596,17'd6211,17'd5482,17'd5332,17'd8154,17'd10515,17'd28057,17'd11316,17'd11037,17'd28305,17'd10897,17'd28058,17'd37031,17'd5336,17'd28418,17'd28418,17'd5329,17'd4845,17'd4686,17'd4840,17'd4996,17'd38442,17'd5144,17'd6067,17'd4995,17'd5328,17'd5328,17'd28418,17'd28418,17'd30637,17'd5160,17'd5002,17'd5329,17'd34921,17'd4999,17'd34157,17'd33839,17'd4356,17'd42772,17'd4185,17'd45393,17'd4017,17'd33839,17'd34157,17'd33992,17'd33841,17'd49597,17'd49598,17'd49599,17'd49600,17'd36738,17'd36037,17'd49601,17'd49602,17'd49603,17'd49604,17'd49504,17'd3562,17'd4054,17'd18756,17'd5025,17'd40099,17'd41159,17'd10388,17'd10790,17'd39181,17'd39483,17'd38580,17'd12913,17'd38072,17'd38072,17'd37959,17'd37959,17'd4883,17'd4713,17'd5630,17'd5630,17'd4713,17'd4882,17'd4713,17'd4729,17'd4729,17'd4713,17'd6415,17'd5957,17'd411,17'd643,17'd261,17'd1097,17'd1093,17'd2420,17'd591,17'd462
},
'{
17'd27713,17'd25384,17'd2784,17'd3250,17'd1831,17'd466,17'd18,17'd18,17'd1278,17'd980,17'd286,17'd1833,17'd467,17'd285,17'd285,17'd26,17'd980,17'd652,17'd289,17'd289,17'd3595,17'd3255,17'd2941,17'd2943,17'd2262,17'd3103,17'd1973,17'd19874,17'd41008,17'd41008,17'd3107,17'd37171,17'd4259,17'd33542,17'd3603,17'd49506,17'd26980,17'd49605,17'd49606,17'd49607,17'd49608,17'd23667,17'd28800,17'd49609,17'd25658,17'd12681,17'd17204,17'd17689,17'd27461,17'd18655,17'd12681,17'd12218,17'd12955,17'd12679,17'd13209,17'd13092,17'd13462,17'd13597,17'd14344,17'd13461,17'd10937,17'd12677,17'd12955,17'd14471,17'd19753,17'd18656,17'd19257,17'd17810,17'd24348,17'd14347,17'd48641,17'd49610,17'd49200,17'd47866,17'd14220,17'd10565,17'd11088,17'd11088,17'd46366,17'd6143,17'd6625,17'd10946,17'd9985,17'd8074,17'd7423,17'd49611,17'd6641,17'd40271,17'd48304,17'd42215,17'd49612,17'd48824,17'd49613,17'd49304,17'd49113,17'd49614,17'd6953,17'd37843,17'd33395,17'd49615,17'd28085,17'd49616,17'd9456,17'd49617,17'd49618,17'd49619,17'd49620,17'd49621,17'd49622,17'd48651,17'd48571,17'd49623,17'd49624,17'd49625,17'd8094,17'd8408,17'd8720,17'd9479,17'd12116,17'd26152,17'd19282,17'd14931,17'd13762,17'd18443,17'd22472,17'd21363,17'd26258,17'd44982,17'd18326,17'd11668,17'd13368,17'd34205,17'd11668,17'd25280,17'd24029,17'd48101,17'd17604,17'd12110,17'd13513,17'd12997,17'd16799,17'd14523,17'd21207,17'd21207,17'd12416,17'd27234,17'd29482,17'd34835,17'd31590,17'd49525,17'd49032,17'd33875,17'd33568,17'd34203,17'd31127,17'd30834,17'd36777,17'd28230,17'd21671,17'd15185,17'd11522,17'd11668,17'd28463,17'd21206,17'd19282,17'd10165,17'd17719,17'd10992,17'd9340,17'd9345,17'd22814,17'd33083,17'd15048,17'd9739,17'd10164,17'd48849,17'd49626,17'd49627,17'd49628,17'd49629,17'd49630,17'd49631,17'd49632,17'd49633,17'd49634,17'd49635,17'd49636,17'd49637,17'd49638,17'd49639,17'd49045,17'd49540,17'd49640,17'd15805,17'd49641,17'd49642,17'd49643,17'd49644,17'd49645,17'd49646,17'd49647,17'd49648,17'd49649,17'd49650,17'd49651,17'd45316,17'd49652,17'd49653,17'd49654,17'd49655,17'd49656,17'd49657,17'd46312,17'd49658,17'd46826,17'd48431,17'd48019,17'd43408,17'd49659,17'd49660,17'd49661,17'd34728,17'd49662,17'd49463,17'd42580,17'd42580,17'd40805,17'd47213,17'd44688,17'd49663,17'd45859,17'd49664,17'd49364,17'd49665,17'd49666,17'd48882,17'd49667,17'd49668,17'd49669,17'd49670,17'd49671,17'd49672,17'd49673,17'd47624,17'd49674,17'd49675,17'd49676,17'd49677,17'd49678,17'd49572,17'd46663,17'd49679,17'd44589,17'd45749,17'd47438,17'd28721,17'd27765,17'd27765,17'd28369,17'd25438,17'd27512,17'd27512,17'd28717,17'd28717,17'd27511,17'd32353,17'd30126,17'd29972,17'd29242,17'd29528,17'd23732,17'd23918,17'd23566,17'd29975,17'd29827,17'd23734,17'd33652,17'd49680,17'd49274,17'd49377,17'd48614,17'd46435,17'd46952,17'd40048,17'd42435,17'd40819,17'd47641,17'd49576,17'd49681,17'd47343,17'd49091,17'd49682,17'd49683,17'd49684,17'd42144,17'd49685,17'd32184,17'd27885,17'd31503,17'd29245,17'd26901,17'd27259,17'd28720,17'd25177,17'd28851,17'd30879,17'd23918,17'd31033,17'd25032,17'd25438,17'd33803,17'd31520,17'd28602,17'd28724,17'd28727,17'd33485,17'd49686,17'd36132,17'd29979,17'd49687,17'd33489,17'd34117,17'd30130,17'd31038,17'd48991,17'd30740,17'd49688,17'd44234,17'd44593,17'd41862,17'd49689,17'd49690,17'd48360,17'd49682,17'd49691,17'd49692,17'd49693,17'd49485,17'd49682,17'd49694,17'd48536,17'd47641,17'd49695,17'd49696,17'd47927,17'd27027,17'd27640,17'd26062,17'd30606,17'd25438,17'd34467,17'd29686,17'd33795,17'd48996,17'd32012,17'd33798,17'd47834,17'd39745,17'd44360,17'd40523,17'd23926,17'd32666,17'd31497,17'd23041,17'd32501,17'd49487,17'd32013,17'd32502,17'd35153,17'd23222,17'd35156,17'd48631,17'd35295,17'd33162,17'd23742,17'd22860,17'd35016,17'd33480,17'd49697,17'd49698,17'd49699,17'd49700,17'd49701,17'd49702,17'd22374,17'd48171,17'd21609,17'd10198,17'd5479,17'd5330,17'd6388,17'd8154,17'd10515,17'd28183,17'd11316,17'd10642,17'd27931,17'd8780,17'd49703,17'd34334,17'd5329,17'd28418,17'd5005,17'd5329,17'd4686,17'd4841,17'd4840,17'd5153,17'd5145,17'd5144,17'd4682,17'd4839,17'd4995,17'd5328,17'd4842,17'd28536,17'd30637,17'd25627,17'd5329,17'd4845,17'd4529,17'd4999,17'd42180,17'd33839,17'd4356,17'd41455,17'd4017,17'd4357,17'd33839,17'd42180,17'd34157,17'd41891,17'd49704,17'd4369,17'd49705,17'd49706,17'd49707,17'd49708,17'd49709,17'd4039,17'd49710,17'd49711,17'd3559,17'd3702,17'd49712,17'd3868,17'd40410,17'd5025,17'd3709,17'd39947,17'd10388,17'd10906,17'd38458,17'd11867,17'd41481,17'd44019,17'd38072,17'd38072,17'd38459,17'd4868,17'd4713,17'd4713,17'd5630,17'd5630,17'd4882,17'd4713,17'd4729,17'd4729,17'd4713,17'd4713,17'd5372,17'd5957,17'd1823,17'd970,17'd258,17'd802,17'd49713,17'd461,17'd612,17'd462
},
'{
17'd27713,17'd4892,17'd2782,17'd3250,17'd1831,17'd1127,17'd16,17'd18,17'd1278,17'd980,17'd286,17'd1833,17'd467,17'd285,17'd285,17'd286,17'd652,17'd652,17'd289,17'd289,17'd3595,17'd3255,17'd2941,17'd2943,17'd2262,17'd3103,17'd1973,17'd1973,17'd1840,17'd41008,17'd3107,17'd2608,17'd4259,17'd33542,17'd3603,17'd49506,17'd26980,17'd5394,17'd20877,17'd49714,17'd49715,17'd23667,17'd28800,17'd49609,17'd25658,17'd22630,17'd19006,17'd17941,17'd18774,17'd18774,17'd12681,17'd12956,17'd11626,17'd12679,17'd13092,17'd12678,17'd13597,17'd13597,17'd14344,17'd14216,17'd11084,17'd12677,17'd12955,17'd14471,17'd19753,17'd17206,17'd19257,17'd19257,17'd17319,17'd14219,17'd48641,17'd49610,17'd49200,17'd47866,17'd14220,17'd15766,17'd20426,17'd9702,17'd7418,17'd5837,17'd6140,17'd10695,17'd9985,17'd8074,17'd7423,17'd49611,17'd6641,17'd40271,17'd49716,17'd42064,17'd43891,17'd48824,17'd49613,17'd44284,17'd46900,17'd49717,17'd49718,17'd38488,17'd49719,17'd49720,17'd9025,17'd49721,17'd49722,17'd49723,17'd49724,17'd49725,17'd49726,17'd49727,17'd49728,17'd48743,17'd49729,17'd49730,17'd49731,17'd49732,17'd49733,17'd49734,17'd9044,17'd9480,17'd9741,17'd10167,17'd19532,17'd10990,17'd13762,17'd16442,17'd22472,17'd21362,17'd33084,17'd44982,17'd37196,17'd28463,17'd34205,17'd34205,17'd11668,17'd25280,17'd24029,17'd41343,17'd30083,17'd14130,17'd19032,17'd12997,17'd13134,17'd14523,17'd21057,17'd21057,17'd12416,17'd16557,17'd28945,17'd30677,17'd33875,17'd34545,17'd34545,17'd33875,17'd33720,17'd34037,17'd32920,17'd32283,17'd31764,17'd36629,17'd24030,17'd18198,17'd14264,17'd11398,17'd11668,17'd11399,17'd19282,17'd10165,17'd10329,17'd21503,17'd9341,17'd9345,17'd15569,17'd16065,17'd15048,17'd9739,17'd10326,17'd29068,17'd49735,17'd49736,17'd49737,17'd49738,17'd49739,17'd49740,17'd49741,17'd49742,17'd49743,17'd49744,17'd49745,17'd49746,17'd49050,17'd48593,17'd48959,17'd49539,17'd22132,17'd49747,17'd15680,17'd49748,17'd49749,17'd49750,17'd49751,17'd49752,17'd47693,17'd49753,17'd49754,17'd48866,17'd49755,17'd49756,17'd49757,17'd49758,17'd49759,17'd49760,17'd49761,17'd49762,17'd47028,17'd49763,17'd49764,17'd46523,17'd49765,17'd49766,17'd49767,17'd49768,17'd49769,17'd47124,17'd49770,17'd49771,17'd39719,17'd47615,17'd46927,17'd47213,17'd40032,17'd40501,17'd46531,17'd46929,17'd39259,17'd44687,17'd48680,17'd49772,17'd49773,17'd49774,17'd49775,17'd49776,17'd47230,17'd49777,17'd49778,17'd49779,17'd49780,17'd49781,17'd49782,17'd49783,17'd49784,17'd49785,17'd46201,17'd44228,17'd44934,17'd33156,17'd44359,17'd29970,17'd33000,17'd27882,17'd25438,17'd27512,17'd27512,17'd25177,17'd28717,17'd28717,17'd29103,17'd25031,17'd34467,17'd29972,17'd34137,17'd33794,17'd29241,17'd23918,17'd23386,17'd29374,17'd31502,17'd29528,17'd30424,17'd49786,17'd46325,17'd49377,17'd49275,17'd46663,17'd47636,17'd39432,17'd41414,17'd49477,17'd49576,17'd49576,17'd48617,17'd47344,17'd49288,17'd49787,17'd49788,17'd49391,17'd40510,17'd43973,17'd33791,17'd33319,17'd29379,17'd31035,17'd26902,17'd25833,17'd28130,17'd28254,17'd24415,17'd24086,17'd23734,17'd24087,17'd25031,17'd27511,17'd31520,17'd28598,17'd25949,17'd27027,17'd37513,17'd32505,17'd49789,17'd29978,17'd49790,17'd34461,17'd33488,17'd33323,17'd30130,17'd29978,17'd33166,17'd49791,17'd49792,17'd44361,17'd44593,17'd41862,17'd49181,17'd49793,17'd48535,17'd49583,17'd49794,17'd49794,17'd49693,17'd49693,17'd49582,17'd49694,17'd48536,17'd47446,17'd48531,17'd40364,17'd43838,17'd26902,17'd27883,17'd26062,17'd30606,17'd25177,17'd24415,17'd29374,17'd33795,17'd43985,17'd40369,17'd32012,17'd32502,17'd30728,17'd44360,17'd32190,17'd23926,17'd32346,17'd48912,17'd33648,17'd32501,17'd49487,17'd32009,17'd23220,17'd35153,17'd48912,17'd49795,17'd48631,17'd48796,17'd49487,17'd22682,17'd30276,17'd39281,17'd35456,17'd49796,17'd49797,17'd49798,17'd49799,17'd49800,17'd49801,17'd49802,17'd49803,17'd21610,17'd7165,17'd5610,17'd5335,17'd6218,17'd9090,17'd10515,17'd28183,17'd11037,17'd10515,17'd27931,17'd9657,17'd5919,17'd41889,17'd5002,17'd28418,17'd5005,17'd5329,17'd4687,17'd4841,17'd4683,17'd5153,17'd5145,17'd5144,17'd4682,17'd4683,17'd5327,17'd5328,17'd28418,17'd28536,17'd30637,17'd25627,17'd5329,17'd5002,17'd4846,17'd41459,17'd46979,17'd33691,17'd39468,17'd41458,17'd4515,17'd4358,17'd42180,17'd4998,17'd33992,17'd34657,17'd49804,17'd4370,17'd49805,17'd38321,17'd49806,17'd49708,17'd35900,17'd49807,17'd49808,17'd49809,17'd49810,17'd3702,17'd49712,17'd40562,17'd6866,17'd5494,17'd3709,17'd41159,17'd48559,17'd10790,17'd39181,17'd38859,17'd38860,17'd38580,17'd38072,17'd38072,17'd38459,17'd38459,17'd4883,17'd4729,17'd5630,17'd5630,17'd4713,17'd4713,17'd4729,17'd4729,17'd4729,17'd4085,17'd5957,17'd5050,17'd1396,17'd259,17'd261,17'd40563,17'd39949,17'd17551,17'd964,17'd462
},
'{
17'd27713,17'd25384,17'd2935,17'd3250,17'd1688,17'd2,17'd19,17'd18,17'd1278,17'd980,17'd286,17'd1833,17'd467,17'd285,17'd285,17'd285,17'd980,17'd652,17'd289,17'd289,17'd3755,17'd3595,17'd3254,17'd2940,17'd3253,17'd3103,17'd2600,17'd19608,17'd1422,17'd41008,17'd2607,17'd2608,17'd4259,17'd33542,17'd3603,17'd28196,17'd26980,17'd49605,17'd49811,17'd49812,17'd24185,17'd49813,17'd22975,17'd23499,17'd23836,17'd16658,17'd12681,17'd19382,17'd18774,17'd17941,17'd11764,17'd13094,17'd12813,17'd12527,17'd13092,17'd15762,17'd13597,17'd14344,17'd14216,17'd14216,17'd11084,17'd12062,17'd13209,17'd14891,17'd20423,17'd18774,17'd27460,17'd19257,17'd17319,17'd14219,17'd49814,17'd48819,17'd33857,17'd14626,17'd14220,17'd10565,17'd10943,17'd11088,17'd9702,17'd6143,17'd6141,17'd10695,17'd9985,17'd8074,17'd7423,17'd49611,17'd6641,17'd39966,17'd40119,17'd40876,17'd42937,17'd43753,17'd49815,17'd43892,17'd44284,17'd49816,17'd49817,17'd46255,17'd35503,17'd8393,17'd27965,17'd29461,17'd49818,17'd49819,17'd27609,17'd49820,17'd24983,17'd49821,17'd49121,17'd49822,17'd49823,17'd49824,17'd49825,17'd49826,17'd49827,17'd49828,17'd49829,17'd9344,17'd9741,17'd21503,17'd10166,17'd10854,17'd11395,17'd15185,17'd16442,17'd22472,17'd22472,17'd18443,17'd30532,17'd22816,17'd13521,17'd13521,17'd11668,17'd25280,17'd11397,17'd14671,17'd18082,17'd11958,17'd12855,17'd13884,17'd14524,17'd14672,17'd14525,17'd14525,17'd14003,17'd19534,17'd28348,17'd29930,17'd34203,17'd31590,17'd34545,17'd33875,17'd33875,17'd34037,17'd34037,17'd33875,17'd31761,17'd29645,17'd24991,17'd21671,17'd16325,17'd11397,17'd18326,17'd11398,17'd11132,17'd11133,17'd10165,17'd17719,17'd27003,17'd27856,17'd15187,17'd16065,17'd15048,17'd9739,17'd10326,17'd10606,17'd28956,17'd49830,17'd49831,17'd49832,17'd49833,17'd49834,17'd49835,17'd49836,17'd49837,17'd49838,17'd49839,17'd49745,17'd49840,17'd48862,17'd49841,17'd49140,17'd49842,17'd49842,17'd49843,17'd49844,17'd49845,17'd49846,17'd49847,17'd49848,17'd49849,17'd49850,17'd49851,17'd49852,17'd49853,17'd49854,17'd49855,17'd49856,17'd49857,17'd49858,17'd49859,17'd49860,17'd41987,17'd49861,17'd49862,17'd49863,17'd47028,17'd47703,17'd49864,17'd49865,17'd39113,17'd46310,17'd46396,17'd49658,17'd49866,17'd43135,17'd44919,17'd49867,17'd34728,17'd47520,17'd38518,17'd39259,17'd49868,17'd34728,17'd49869,17'd49870,17'd35408,17'd49871,17'd49872,17'd49873,17'd49874,17'd49875,17'd49876,17'd49877,17'd49878,17'd49879,17'd49782,17'd47442,17'd49375,17'd49880,17'd48526,17'd43548,17'd33156,17'd49273,17'd42749,17'd25438,17'd28717,17'd28717,17'd25568,17'd28719,17'd27512,17'd25177,17'd25177,17'd27637,17'd29533,17'd28851,17'd24902,17'd29689,17'd23565,17'd31029,17'd29528,17'd34137,17'd29830,17'd29827,17'd29528,17'd29375,17'd33317,17'd49881,17'd49882,17'd46326,17'd49476,17'd47627,17'd49375,17'd42596,17'd47936,17'd49576,17'd48904,17'd49280,17'd49586,17'd47737,17'd49390,17'd49883,17'd49884,17'd49885,17'd49886,17'd45745,17'd37908,17'd40681,17'd29245,17'd30586,17'd28724,17'd32658,17'd27511,17'd24744,17'd28849,17'd23920,17'd23734,17'd24087,17'd29533,17'd28369,17'd31055,17'd27766,17'd26903,17'd33163,17'd29977,17'd36989,17'd49789,17'd29978,17'd49790,17'd34461,17'd49887,17'd33488,17'd30280,17'd29831,17'd29249,17'd49888,17'd36401,17'd41863,17'd44479,17'd45157,17'd48144,17'd49889,17'd48622,17'd49693,17'd49890,17'd49890,17'd49891,17'd49692,17'd49582,17'd49684,17'd48154,17'd47446,17'd43688,17'd46760,17'd33155,17'd28725,17'd27514,17'd26062,17'd27513,17'd25568,17'd30879,17'd37386,17'd33795,17'd43985,17'd40369,17'd32501,17'd33312,17'd31834,17'd33645,17'd44591,17'd30728,17'd32829,17'd33162,17'd31832,17'd49892,17'd31344,17'd32009,17'd32009,17'd31030,17'd36692,17'd32347,17'd48625,17'd32188,17'd47346,17'd22681,17'd30276,17'd35157,17'd23221,17'd47460,17'd46963,17'd49893,17'd35458,17'd44498,17'd45503,17'd21737,17'd49894,17'd26582,17'd7009,17'd5481,17'd27935,17'd6553,17'd9657,17'd27815,17'd27933,17'd11038,17'd10515,17'd9657,17'd8154,17'd5762,17'd5329,17'd29024,17'd4685,17'd5005,17'd5329,17'd4687,17'd4686,17'd4683,17'd5153,17'd5145,17'd5145,17'd4995,17'd4683,17'd5328,17'd5328,17'd37153,17'd37153,17'd30637,17'd25627,17'd5329,17'd4845,17'd4529,17'd4999,17'd34157,17'd42180,17'd33840,17'd33533,17'd4833,17'd33838,17'd33991,17'd41891,17'd41891,17'd5154,17'd49895,17'd49896,17'd49805,17'd49897,17'd49898,17'd36174,17'd49899,17'd49900,17'd49901,17'd42783,17'd49902,17'd41624,17'd40861,17'd8787,17'd6082,17'd5494,17'd3709,17'd41159,17'd48559,17'd10906,17'd38458,17'd11867,17'd38334,17'd38580,17'd38072,17'd38072,17'd4867,17'd4883,17'd4729,17'd4729,17'd8185,17'd5630,17'd4713,17'd4729,17'd4729,17'd4729,17'd4085,17'd4085,17'd2392,17'd1680,17'd1243,17'd271,17'd1097,17'd2255,17'd186,17'd461,17'd2251,17'd2251
},
'{
17'd27713,17'd4892,17'd2593,17'd3250,17'd1688,17'd14,17'd1277,17'd18,17'd1278,17'd980,17'd27,17'd286,17'd467,17'd285,17'd285,17'd286,17'd652,17'd652,17'd289,17'd289,17'd3755,17'd3255,17'd2941,17'd2943,17'd2262,17'd3103,17'd2600,17'd2600,17'd1702,17'd41008,17'd2607,17'd3757,17'd2786,17'd33850,17'd33851,17'd30349,17'd27100,17'd5394,17'd49903,17'd49904,17'd24515,17'd49905,17'd18527,17'd49906,17'd25658,17'd16658,17'd12532,17'd19382,17'd17689,17'd17941,17'd11764,17'd12065,17'd12527,17'd12527,17'd13092,17'd15762,17'd13597,17'd13461,17'd14216,17'd14216,17'd11084,17'd12062,17'd13209,17'd14764,17'd12681,17'd18774,17'd27460,17'd27833,17'd17319,17'd14219,17'd49814,17'd48819,17'd48387,17'd14626,17'd14220,17'd15766,17'd15765,17'd9574,17'd8537,17'd7418,17'd6141,17'd10695,17'd9985,17'd8074,17'd7423,17'd49611,17'd6641,17'd39966,17'd40119,17'd40876,17'd42937,17'd43753,17'd49815,17'd45198,17'd44284,17'd49907,17'd42940,17'd39351,17'd35635,17'd49908,17'd30061,17'd49909,17'd28444,17'd49910,17'd49911,17'd49912,17'd24202,17'd26616,17'd26487,17'd49314,17'd49913,17'd49914,17'd49915,17'd49916,17'd49917,17'd49918,17'd49919,17'd9344,17'd12116,17'd10024,17'd26152,17'd19282,17'd14673,17'd13762,17'd16442,17'd22472,17'd22472,17'd18443,17'd22817,17'd19533,17'd13521,17'd13521,17'd11668,17'd11398,17'd11397,17'd19643,17'd49920,17'd17603,17'd12859,17'd13884,17'd14524,17'd14524,17'd14930,17'd14525,17'd14003,17'd21504,17'd27234,17'd28944,17'd34381,17'd34037,17'd31590,17'd34545,17'd33720,17'd34037,17'd31590,17'd33875,17'd31762,17'd34551,17'd28103,17'd20452,17'd11959,17'd19158,17'd21985,17'd25280,17'd10476,17'd11132,17'd19282,17'd10165,17'd46267,17'd27003,17'd10742,17'd11809,17'd15048,17'd14928,17'd10326,17'd11528,17'd46726,17'd49735,17'd49921,17'd49922,17'd49923,17'd49924,17'd49925,17'd49926,17'd49927,17'd49928,17'd49929,17'd49930,17'd49931,17'd49932,17'd49933,17'd49934,17'd49842,17'd49935,17'd49936,17'd49937,17'd49938,17'd49939,17'd49940,17'd49941,17'd49942,17'd49943,17'd49944,17'd49945,17'd49946,17'd49947,17'd49948,17'd35389,17'd49949,17'd49950,17'd49951,17'd49952,17'd49953,17'd49954,17'd49955,17'd49956,17'd47906,17'd46192,17'd49957,17'd49958,17'd49959,17'd45858,17'd46738,17'd48344,17'd42864,17'd48230,17'd49960,17'd49961,17'd49560,17'd40501,17'd49866,17'd49962,17'd44687,17'd39886,17'd49963,17'd47032,17'd49964,17'd49965,17'd49966,17'd49967,17'd49968,17'd49969,17'd49970,17'd49971,17'd49972,17'd49973,17'd49974,17'd49272,17'd46841,17'd49081,17'd49975,17'd46095,17'd43978,17'd32996,17'd25438,17'd33951,17'd25177,17'd27512,17'd28719,17'd28719,17'd25568,17'd25320,17'd29976,17'd24895,17'd28851,17'd30879,17'd29972,17'd23565,17'd23733,17'd23734,17'd29241,17'd23386,17'd29830,17'd29099,17'd32186,17'd30424,17'd49976,17'd49977,17'd49978,17'd46326,17'd46436,17'd47531,17'd48522,17'd49379,17'd49586,17'd48154,17'd49979,17'd49280,17'd47736,17'd43541,17'd49693,17'd49980,17'd49981,17'd48450,17'd44586,17'd41270,17'd31353,17'd37513,17'd28727,17'd27027,17'd25707,17'd25435,17'd25320,17'd28601,17'd29689,17'd23734,17'd24421,17'd24086,17'd25179,17'd25317,17'd28598,17'd25707,17'd28725,17'd30735,17'd33319,17'd34114,17'd32019,17'd29978,17'd30131,17'd33323,17'd49982,17'd33488,17'd30280,17'd29979,17'd36989,17'd49983,17'd38152,17'd41863,17'd44479,17'd40216,17'd48260,17'd48781,17'd43419,17'd49984,17'd49985,17'd49986,17'd49987,17'd49891,17'd49988,17'd49989,17'd49382,17'd48446,17'd43831,17'd47635,17'd44231,17'd28725,17'd27514,17'd26062,17'd27513,17'd27512,17'd28722,17'd37117,17'd31194,17'd43985,17'd31661,17'd49588,17'd46677,17'd31834,17'd35158,17'd44591,17'd30728,17'd33649,17'd33796,17'd35156,17'd33796,17'd21845,17'd23220,17'd32013,17'd21850,17'd21695,17'd49990,17'd48625,17'd49892,17'd32346,17'd30276,17'd30276,17'd23394,17'd49991,17'd46218,17'd46963,17'd49992,17'd49993,17'd29864,17'd49994,17'd19459,17'd22080,17'd10882,17'd27695,17'd5158,17'd27935,17'd8303,17'd10513,17'd27815,17'd27933,17'd11038,17'd27815,17'd9657,17'd6553,17'd5330,17'd4687,17'd37153,17'd4685,17'd5005,17'd5329,17'd4845,17'd4686,17'd5328,17'd5153,17'd4996,17'd5145,17'd4995,17'd4683,17'd5328,17'd5328,17'd37153,17'd37153,17'd5004,17'd25627,17'd5329,17'd5002,17'd4847,17'd41459,17'd33992,17'd42180,17'd33691,17'd33691,17'd4189,17'd4999,17'd41891,17'd33841,17'd5154,17'd41459,17'd49995,17'd49996,17'd49997,17'd4201,17'd49898,17'd36174,17'd49998,17'd49999,17'd50000,17'd47381,17'd2888,17'd41479,17'd50001,17'd50002,17'd40410,17'd3567,17'd3709,17'd41159,17'd10388,17'd45186,17'd39790,17'd39033,17'd38860,17'd38580,17'd38072,17'd38072,17'd4867,17'd4883,17'd4729,17'd4729,17'd8185,17'd5630,17'd4713,17'd4729,17'd4729,17'd4729,17'd4085,17'd4085,17'd445,17'd1680,17'd1243,17'd207,17'd408,17'd2115,17'd405,17'd17551,17'd1822,17'd2251
},
'{
17'd27713,17'd25384,17'd2935,17'd3250,17'd2597,17'd17,17'd19,17'd18,17'd1278,17'd980,17'd27,17'd286,17'd467,17'd285,17'd285,17'd285,17'd27,17'd652,17'd289,17'd289,17'd3755,17'd3595,17'd3254,17'd2941,17'd3253,17'd3103,17'd2600,17'd19608,17'd1422,17'd2607,17'd3597,17'd3915,17'd33378,17'd33542,17'd3758,17'd29306,17'd5066,17'd50003,17'd21175,17'd50004,17'd13824,17'd23497,17'd18527,17'd23499,17'd22117,17'd16765,17'd12532,17'd20423,17'd19382,17'd19382,17'd13969,17'd12065,17'd12527,17'd14469,17'd13462,17'd13597,17'd14344,17'd13461,17'd14216,17'd13460,17'd12355,17'd12215,17'd13092,17'd14621,17'd22630,17'd19128,17'd27460,17'd19257,17'd17319,17'd14220,17'd34178,17'd50005,17'd48387,17'd14626,17'd14220,17'd10565,17'd10944,17'd10943,17'd9702,17'd7418,17'd6141,17'd7085,17'd49201,17'd8846,17'd7756,17'd39646,17'd50006,17'd6483,17'd39813,17'd49716,17'd42064,17'd43891,17'd50007,17'd45198,17'd43892,17'd44760,17'd45411,17'd50008,17'd47874,17'd50009,17'd8393,17'd28672,17'd27841,17'd28330,17'd50010,17'd50011,17'd50012,17'd50013,17'd50014,17'd49728,17'd50015,17'd50016,17'd50017,17'd50018,17'd8714,17'd50019,17'd50020,17'd47889,17'd24037,17'd10856,17'd15300,17'd10472,17'd10737,17'd11395,17'd16204,17'd16204,17'd15185,17'd15185,17'd11964,17'd13645,17'd11130,17'd11130,17'd11275,17'd11808,17'd13645,17'd13645,17'd18082,17'd12581,17'd12575,17'd13884,17'd14524,17'd15687,17'd15811,17'd22297,17'd14003,17'd21504,17'd16557,17'd28350,17'd30073,17'd31288,17'd35644,17'd31590,17'd33875,17'd34037,17'd31590,17'd34545,17'd33720,17'd50021,17'd29480,17'd24704,17'd19407,17'd18197,17'd23169,17'd11397,17'd11399,17'd11132,17'd11130,17'd14132,17'd41036,17'd9612,17'd17011,17'd9619,17'd19279,17'd22131,17'd10330,17'd12863,17'd50022,17'd24543,17'd17123,17'd49325,17'd50023,17'd50024,17'd50025,17'd49628,17'd50026,17'd50027,17'd50028,17'd49838,17'd50029,17'd50030,17'd50031,17'd50032,17'd50033,17'd50034,17'd50035,17'd49541,17'd14929,17'd26497,17'd24034,17'd14803,17'd50036,17'd49332,17'd50037,17'd50038,17'd50039,17'd50040,17'd50041,17'd50042,17'd50043,17'd50044,17'd50045,17'd50046,17'd50047,17'd38385,17'd50048,17'd50049,17'd40031,17'd50050,17'd50051,17'd46410,17'd50052,17'd47028,17'd46925,17'd46925,17'd46528,17'd46926,17'd50053,17'd50054,17'd45974,17'd47028,17'd50055,17'd49962,17'd49463,17'd48976,17'd50056,17'd42865,17'd50057,17'd50058,17'd50059,17'd50060,17'd50061,17'd49876,17'd50062,17'd50063,17'd50064,17'd50065,17'd50066,17'd50067,17'd48614,17'd48445,17'd50068,17'd43285,17'd43549,17'd28850,17'd28974,17'd28596,17'd25178,17'd27764,17'd27764,17'd25568,17'd29244,17'd29976,17'd25032,17'd29688,17'd23731,17'd23384,17'd29687,17'd23918,17'd23920,17'd23733,17'd31502,17'd29830,17'd23386,17'd23734,17'd24087,17'd34883,17'd50069,17'd46434,17'd50070,17'd46326,17'd46663,17'd47048,17'd39581,17'd40819,17'd43147,17'd48536,17'd49382,17'd47736,17'd48909,17'd49289,17'd49890,17'd49683,17'd50071,17'd48149,17'd44476,17'd33309,17'd31353,17'd29246,17'd28979,17'd28853,17'd25565,17'd29825,17'd25030,17'd28975,17'd29689,17'd31502,17'd23387,17'd23564,17'd25179,17'd28130,17'd30606,17'd26903,17'd26782,17'd29245,17'd32192,17'd29833,17'd32019,17'd30131,17'd30131,17'd33489,17'd49982,17'd49887,17'd30280,17'd36132,17'd38026,17'd35706,17'd38152,17'd41863,17'd44479,17'd40216,17'd47341,17'd47735,17'd49289,17'd49984,17'd49986,17'd50072,17'd49985,17'd49890,17'd49794,17'd49989,17'd49382,17'd48446,17'd46438,17'd46433,17'd44231,17'd27259,17'd27514,17'd26062,17'd27513,17'd27512,17'd23732,17'd23216,17'd44360,17'd48996,17'd31661,17'd34455,17'd33945,17'd23926,17'd34278,17'd44591,17'd23393,17'd34455,17'd21695,17'd35156,17'd33162,17'd49488,17'd23220,17'd21845,17'd22013,17'd21696,17'd32828,17'd50073,17'd49588,17'd23393,17'd30276,17'd22681,17'd46677,17'd45373,17'd50074,17'd50075,17'd50076,17'd50077,17'd50078,17'd50079,17'd50080,17'd22241,17'd10198,17'd5612,17'd30638,17'd6554,17'd8303,17'd10513,17'd27815,17'd28183,17'd10778,17'd7669,17'd6219,17'd26218,17'd4845,17'd32552,17'd4847,17'd4685,17'd5005,17'd5329,17'd5002,17'd4686,17'd5327,17'd5153,17'd4996,17'd42910,17'd4995,17'd4683,17'd5328,17'd5328,17'd37153,17'd29024,17'd5004,17'd25627,17'd5329,17'd4845,17'd4689,17'd5155,17'd41891,17'd4998,17'd47660,17'd4998,17'd4525,17'd5000,17'd33841,17'd41459,17'd5154,17'd41459,17'd40397,17'd50081,17'd49805,17'd38447,17'd50082,17'd36314,17'd50083,17'd50084,17'd50085,17'd50086,17'd50087,17'd3217,17'd50088,17'd50002,17'd7191,17'd50089,17'd3709,17'd39947,17'd10790,17'd50090,17'd11867,17'd44742,17'd41481,17'd38580,17'd38072,17'd38072,17'd4867,17'd4883,17'd3744,17'd35907,17'd12026,17'd12496,17'd1946,17'd4085,17'd4085,17'd4085,17'd4422,17'd1810,17'd2417,17'd1262,17'd1243,17'd258,17'd408,17'd2115,17'd405,17'd17551,17'd1822,17'd1822
},
'{
17'd4243,17'd4892,17'd2593,17'd3250,17'd2597,17'd1415,17'd1277,17'd18,17'd1278,17'd980,17'd27,17'd286,17'd285,17'd285,17'd285,17'd286,17'd28,17'd652,17'd289,17'd289,17'd3755,17'd3255,17'd3431,17'd2942,17'd2262,17'd3103,17'd2600,17'd1973,17'd1840,17'd2432,17'd2607,17'd3757,17'd4259,17'd33850,17'd33542,17'd29449,17'd50091,17'd21799,17'd50092,17'd50004,17'd13824,17'd23497,17'd50093,17'd22976,17'd22117,17'd16765,17'd12531,17'd19382,17'd19128,17'd19382,17'd13969,17'd12065,17'd12679,17'd22802,17'd14469,17'd13597,17'd13461,17'd13461,17'd13460,17'd13326,17'd13460,17'd12215,17'd13092,17'd14621,17'd16658,17'd19128,17'd27460,17'd19008,17'd17572,17'd14220,17'd34178,17'd50094,17'd48387,17'd14626,17'd14220,17'd16880,17'd11231,17'd9574,17'd8537,17'd6143,17'd6141,17'd7085,17'd49201,17'd8846,17'd7756,17'd49112,17'd47094,17'd6483,17'd40582,17'd50095,17'd42666,17'd42937,17'd50007,17'd50096,17'd50097,17'd43354,17'd42669,17'd48193,17'd48084,17'd49115,17'd32428,17'd50098,17'd50099,17'd9322,17'd50100,17'd50101,17'd50102,17'd49820,17'd50103,17'd26251,17'd50104,17'd50105,17'd28808,17'd50106,17'd50107,17'd50108,17'd50109,17'd47889,17'd9478,17'd17011,17'd10856,17'd10165,17'd10739,17'd10736,17'd13362,17'd16204,17'd15185,17'd15185,17'd13762,17'd13645,17'd11275,17'd11275,17'd11808,17'd11808,17'd13645,17'd18444,17'd50110,17'd18558,17'd12417,17'd16559,17'd15571,17'd15687,17'd15811,17'd22297,17'd21504,17'd21504,17'd16913,17'd27348,17'd29198,17'd31289,17'd35644,17'd50111,17'd31590,17'd34380,17'd35644,17'd31590,17'd33875,17'd34381,17'd28686,17'd28103,17'd12255,17'd20314,17'd14258,17'd18327,17'd11524,17'd11399,17'd19533,17'd11130,17'd10472,17'd10741,17'd9883,17'd11277,17'd24998,17'd24998,17'd10331,17'd11670,17'd25530,17'd50112,17'd10174,17'd34039,17'd50113,17'd50114,17'd50115,17'd49628,17'd23344,17'd50116,17'd50117,17'd50118,17'd50119,17'd50029,17'd50120,17'd49942,17'd49442,17'd50121,17'd50121,17'd49335,17'd49441,17'd15432,17'd16064,17'd20908,17'd31130,17'd50122,17'd50123,17'd50124,17'd50125,17'd49945,17'd50126,17'd50127,17'd50128,17'd50129,17'd50130,17'd50131,17'd50132,17'd50133,17'd50134,17'd44089,17'd41851,17'd48125,17'd44687,17'd50135,17'd50136,17'd50137,17'd46525,17'd40346,17'd47906,17'd50138,17'd47124,17'd49662,17'd50139,17'd46405,17'd46291,17'd43135,17'd33451,17'd35263,17'd50140,17'd49462,17'd50141,17'd50142,17'd50143,17'd50144,17'd50145,17'd50146,17'd50147,17'd50148,17'd50149,17'd50150,17'd50151,17'd47436,17'd50152,17'd42742,17'd50153,17'd50154,17'd50155,17'd24744,17'd23561,17'd25180,17'd24898,17'd28596,17'd27764,17'd25568,17'd25320,17'd25180,17'd28851,17'd29534,17'd34137,17'd29827,17'd23386,17'd31502,17'd29241,17'd23918,17'd23566,17'd29830,17'd23566,17'd29528,17'd32186,17'd50156,17'd50157,17'd50157,17'd46326,17'd50158,17'd46758,17'd50159,17'd42435,17'd49477,17'd48263,17'd48536,17'd48154,17'd48264,17'd43419,17'd49682,17'd50160,17'd49788,17'd50161,17'd48041,17'd44823,17'd36690,17'd31353,17'd29245,17'd28486,17'd28725,17'd25566,17'd31034,17'd24745,17'd29102,17'd34137,17'd23566,17'd36987,17'd23384,17'd25179,17'd28600,17'd26062,17'd27259,17'd26781,17'd29379,17'd33321,17'd29981,17'd33322,17'd30131,17'd30131,17'd30736,17'd31505,17'd31506,17'd30280,17'd36132,17'd50162,17'd35424,17'd42882,17'd42739,17'd44479,17'd40216,17'd47535,17'd47828,17'd49484,17'd50163,17'd50072,17'd50072,17'd49986,17'd50164,17'd49683,17'd49989,17'd49382,17'd48709,17'd44930,17'd46201,17'd42147,17'd27259,17'd26530,17'd28481,17'd30734,17'd28719,17'd30275,17'd23216,17'd44360,17'd48996,17'd44109,17'd31497,17'd50165,17'd23926,17'd44591,17'd34278,17'd32503,17'd49588,17'd23044,17'd22510,17'd34457,17'd32665,17'd32009,17'd31497,17'd36545,17'd33161,17'd50166,17'd49095,17'd47346,17'd31834,17'd22856,17'd23926,17'd50167,17'd50168,17'd50074,17'd50169,17'd50170,17'd50171,17'd50172,17'd50173,17'd50174,17'd24790,17'd6842,17'd50175,17'd31717,17'd6554,17'd8303,17'd10513,17'd27815,17'd10642,17'd8934,17'd7499,17'd26708,17'd5003,17'd4840,17'd4840,17'd4847,17'd37153,17'd5005,17'd5329,17'd5329,17'd4842,17'd5327,17'd5152,17'd5153,17'd4995,17'd4683,17'd4683,17'd4841,17'd4841,17'd37153,17'd5008,17'd30333,17'd30333,17'd25627,17'd5002,17'd4847,17'd5155,17'd33841,17'd33992,17'd4998,17'd33992,17'd5001,17'd5001,17'd41459,17'd5155,17'd41459,17'd5155,17'd4684,17'd4528,17'd50176,17'd4201,17'd50177,17'd50178,17'd50179,17'd50180,17'd45654,17'd50086,17'd50181,17'd50182,17'd50183,17'd50184,17'd50185,17'd43742,17'd41159,17'd39947,17'd10790,17'd45403,17'd50186,17'd12176,17'd38580,17'd38580,17'd38072,17'd38072,17'd4867,17'd3896,17'd3744,17'd3744,17'd8185,17'd5630,17'd4728,17'd4085,17'd3391,17'd4085,17'd4422,17'd1810,17'd2417,17'd1263,17'd970,17'd261,17'd40563,17'd2115,17'd50187,17'd17551,17'd1822,17'd964
},
'{
17'd4243,17'd25384,17'd2935,17'd2422,17'd2597,17'd17,17'd19,17'd18,17'd1278,17'd980,17'd27,17'd286,17'd285,17'd285,17'd285,17'd285,17'd27,17'd652,17'd289,17'd289,17'd3755,17'd3595,17'd3255,17'd2941,17'd3253,17'd3103,17'd1973,17'd19874,17'd2431,17'd3911,17'd3597,17'd3915,17'd33378,17'd33542,17'd30812,17'd3271,17'd4440,17'd50188,17'd50092,17'd20140,17'd13824,17'd19374,17'd50093,17'd22976,17'd50189,17'd14470,17'd16765,17'd20423,17'd19382,17'd19006,17'd12361,17'd12065,17'd12527,17'd14469,17'd13462,17'd13597,17'd13461,17'd14216,17'd13326,17'd13326,17'd13460,17'd12355,17'd14469,17'd12955,17'd13969,17'd19006,17'd50190,17'd27460,17'd17206,17'd24348,17'd32260,17'd50191,17'd48387,17'd14626,17'd14220,17'd29623,17'd10944,17'd10943,17'd9702,17'd6143,17'd6142,17'd6625,17'd50192,17'd6304,17'd8073,17'd7423,17'd6782,17'd46895,17'd49414,17'd40120,17'd42506,17'd42666,17'd50193,17'd50096,17'd50097,17'd46899,17'd50194,17'd50195,17'd50196,17'd35635,17'd50197,17'd50198,17'd50199,17'd50200,17'd50201,17'd27470,17'd50202,17'd27112,17'd50103,17'd50203,17'd50204,17'd50205,17'd50206,17'd50207,17'd50208,17'd50209,17'd50210,17'd50211,17'd18194,17'd17011,17'd10856,17'd25811,17'd24703,17'd10737,17'd19157,17'd13362,17'd11963,17'd11963,17'd13362,17'd12115,17'd11965,17'd11965,17'd11274,17'd11274,17'd13516,17'd12115,17'd50212,17'd18329,17'd13517,17'd12860,17'd15687,17'd15687,17'd18449,17'd15811,17'd21504,17'd21504,17'd19534,17'd27486,17'd36347,17'd34381,17'd31590,17'd31590,17'd34037,17'd34037,17'd34037,17'd34037,17'd34037,17'd34203,17'd29785,17'd50213,17'd34213,17'd19407,17'd20608,17'd17478,17'd17236,17'd11524,17'd24029,17'd14671,17'd24708,17'd10325,17'd10164,17'd11135,17'd24998,17'd19279,17'd10331,17'd12585,17'd11528,17'd15431,17'd15187,17'd15684,17'd50214,17'd50215,17'd50216,17'd50217,17'd50218,17'd50219,17'd50220,17'd50221,17'd50222,17'd50223,17'd50224,17'd50225,17'd50226,17'd50227,17'd50228,17'd49747,17'd28108,17'd15679,17'd50229,17'd28236,17'd15182,17'd50230,17'd50231,17'd50232,17'd50233,17'd50234,17'd50235,17'd50236,17'd50237,17'd50238,17'd50239,17'd50240,17'd50241,17'd50242,17'd50243,17'd50244,17'd45857,17'd46062,17'd46062,17'd50245,17'd50245,17'd50246,17'd40196,17'd40196,17'd38936,17'd50247,17'd50248,17'd50249,17'd46406,17'd50250,17'd46309,17'd48775,17'd40661,17'd47803,17'd47803,17'd50251,17'd50252,17'd50253,17'd50254,17'd50255,17'd50256,17'd50257,17'd50258,17'd50259,17'd50260,17'd50261,17'd50262,17'd50263,17'd50264,17'd43155,17'd44105,17'd50155,17'd30424,17'd29972,17'd24743,17'd24895,17'd24744,17'd24898,17'd25178,17'd25568,17'd28254,17'd24897,17'd34467,17'd24086,17'd29827,17'd23387,17'd29376,17'd31502,17'd23920,17'd23565,17'd29826,17'd29826,17'd29099,17'd29241,17'd33652,17'd50265,17'd50266,17'd50266,17'd50158,17'd48611,17'd46842,17'd42738,17'd46847,17'd49576,17'd48536,17'd49184,17'd43147,17'd48264,17'd48995,17'd50267,17'd50268,17'd49788,17'd40508,17'd44697,17'd45878,17'd31353,17'd32016,17'd31035,17'd28486,17'd27259,17'd28600,17'd30432,17'd24742,17'd29378,17'd28976,17'd29826,17'd32352,17'd30275,17'd32353,17'd25435,17'd25833,17'd28853,17'd28486,17'd27642,17'd32193,17'd30885,17'd33322,17'd30131,17'd30280,17'd31036,17'd31036,17'd30736,17'd30131,17'd29831,17'd50269,17'd35704,17'd45611,17'd50270,17'd46948,17'd44475,17'd48908,17'd47936,17'd49682,17'd50271,17'd50272,17'd50273,17'd50072,17'd49986,17'd49890,17'd49989,17'd48154,17'd48787,17'd46946,17'd46203,17'd32995,17'd27259,17'd26530,17'd26064,17'd28599,17'd28719,17'd30275,17'd23216,17'd44360,17'd48996,17'd44109,17'd21846,17'd50165,17'd32350,17'd44591,17'd40523,17'd32346,17'd44109,17'd48796,17'd32010,17'd50274,17'd32665,17'd32346,17'd34455,17'd36129,17'd41585,17'd47948,17'd48717,17'd32829,17'd39281,17'd22856,17'd22333,17'd31830,17'd50275,17'd47742,17'd50276,17'd50277,17'd50278,17'd50279,17'd50280,17'd50281,17'd25995,17'd6212,17'd30638,17'd50282,17'd36586,17'd8933,17'd10777,17'd9933,17'd10515,17'd7669,17'd50283,17'd33369,17'd50284,17'd4995,17'd5757,17'd4847,17'd29024,17'd5002,17'd5329,17'd5329,17'd4842,17'd5327,17'd5152,17'd5153,17'd4683,17'd4683,17'd4683,17'd4841,17'd4841,17'd37153,17'd5009,17'd30638,17'd25627,17'd5329,17'd4845,17'd5156,17'd5155,17'd4999,17'd41891,17'd33992,17'd33841,17'd4529,17'd4689,17'd5155,17'd4526,17'd5155,17'd4526,17'd4847,17'd4528,17'd50176,17'd38447,17'd50082,17'd50285,17'd50286,17'd50287,17'd50288,17'd2534,17'd50289,17'd50290,17'd50183,17'd40715,17'd50185,17'd3708,17'd3871,17'd39947,17'd10790,17'd50090,17'd44742,17'd50291,17'd41481,17'd38580,17'd38072,17'd4867,17'd4883,17'd3896,17'd3744,17'd35907,17'd12026,17'd12496,17'd6415,17'd4085,17'd3391,17'd3391,17'd1810,17'd2392,17'd1680,17'd954,17'd1679,17'd1097,17'd2115,17'd2115,17'd50187,17'd17551,17'd431,17'd964
},
'{
17'd4243,17'd25384,17'd2935,17'd2422,17'd2597,17'd1415,17'd1277,17'd18,17'd1278,17'd980,17'd27,17'd286,17'd285,17'd285,17'd285,17'd285,17'd27,17'd652,17'd289,17'd289,17'd3755,17'd3595,17'd3255,17'd2941,17'd3253,17'd3103,17'd1973,17'd2122,17'd1975,17'd2606,17'd2607,17'd3757,17'd33378,17'd33542,17'd30812,17'd29449,17'd4267,17'd12341,17'd50292,17'd20417,17'd50293,17'd19374,17'd50294,17'd22976,17'd50189,17'd14470,17'd12361,17'd20423,17'd19006,17'd12681,17'd12361,17'd11626,17'd12527,17'd22802,17'd14469,17'd13597,17'd13461,17'd14216,17'd13460,17'd13460,17'd13460,17'd12355,17'd14469,17'd13210,17'd12361,17'd19006,17'd50190,17'd41320,17'd17206,17'd15899,17'd32101,17'd34522,17'd48387,17'd15384,17'd14219,17'd16880,17'd11231,17'd10943,17'd46366,17'd6143,17'd6142,17'd6625,17'd50192,17'd6304,17'd8073,17'd7260,17'd47187,17'd46895,17'd49414,17'd40120,17'd50295,17'd42666,17'd41925,17'd50296,17'd42668,17'd46899,17'd50194,17'd45411,17'd39202,17'd48935,17'd50297,17'd50298,17'd50299,17'd27606,17'd50300,17'd50301,17'd50302,17'd50303,17'd49725,17'd50304,17'd25919,17'd50305,17'd50306,17'd50307,17'd50308,17'd50309,17'd50310,17'd50311,17'd18194,17'd9619,17'd25673,17'd10023,17'd16555,17'd10737,17'd11395,17'd15186,17'd11963,17'd11963,17'd13362,17'd12115,17'd11965,17'd10989,17'd13516,17'd13516,17'd13516,17'd12422,17'd50312,17'd50313,17'd17348,17'd12860,17'd14930,17'd15687,17'd18449,17'd50314,17'd21504,17'd21504,17'd21504,17'd16557,17'd50213,17'd30221,17'd33875,17'd31590,17'd31590,17'd31590,17'd34545,17'd34037,17'd34037,17'd31288,17'd30221,17'd30373,17'd37206,17'd24033,17'd26035,17'd23513,17'd25280,17'd11398,17'd24029,17'd14671,17'd25144,17'd10475,17'd19282,17'd12863,17'd16070,17'd11277,17'd17847,17'd12585,17'd10479,17'd15681,17'd34204,17'd9189,17'd16071,17'd13371,17'd50315,17'd50316,17'd50317,17'd50219,17'd50318,17'd50319,17'd50320,17'd50321,17'd50322,17'd49735,17'd50323,17'd50324,17'd49540,17'd50325,17'd14665,17'd15564,17'd15679,17'd13885,17'd13253,17'd16068,17'd20610,17'd50326,17'd50123,17'd50327,17'd50328,17'd50329,17'd50330,17'd50331,17'd49755,17'd50332,17'd50333,17'd50334,17'd50335,17'd50336,17'd50337,17'd40943,17'd50338,17'd50339,17'd50340,17'd50341,17'd50342,17'd40346,17'd46289,17'd50343,17'd50344,17'd50345,17'd50346,17'd41851,17'd43408,17'd50347,17'd46398,17'd48685,17'd47803,17'd50348,17'd50349,17'd50350,17'd50351,17'd50352,17'd50353,17'd50354,17'd50355,17'd50356,17'd50357,17'd50358,17'd50359,17'd50360,17'd50361,17'd50154,17'd50362,17'd50363,17'd29374,17'd32352,17'd24249,17'd24743,17'd28718,17'd25180,17'd30432,17'd25180,17'd24896,17'd24742,17'd30879,17'd28976,17'd23386,17'd23387,17'd31502,17'd31502,17'd23733,17'd29099,17'd29374,17'd23387,17'd29099,17'd23920,17'd50364,17'd50360,17'd50157,17'd49977,17'd48898,17'd46663,17'd47148,17'd42879,17'd48446,17'd48904,17'd48708,17'd48708,17'd48904,17'd48264,17'd49682,17'd49788,17'd50365,17'd49479,17'd40046,17'd50366,17'd32185,17'd29379,17'd29245,17'd31035,17'd28486,17'd26903,17'd28484,17'd25179,17'd24252,17'd29972,17'd23923,17'd37386,17'd50367,17'd30879,17'd29101,17'd27766,17'd28724,17'd27027,17'd28727,17'd30279,17'd33656,17'd31839,17'd50368,17'd30131,17'd30280,17'd31036,17'd31036,17'd30736,17'd49790,17'd29536,17'd50369,17'd37906,17'd45747,17'd47045,17'd44592,17'd43546,17'd47733,17'd47641,17'd49692,17'd50370,17'd50371,17'd50273,17'd50072,17'd49986,17'd49683,17'd49684,17'd48904,17'd46847,17'd44588,17'd46102,17'd33792,17'd27640,17'd28482,17'd30606,17'd31055,17'd25029,17'd30275,17'd23389,17'd46958,17'd48996,17'd45153,17'd32013,17'd46454,17'd32350,17'd44591,17'd34107,17'd32829,17'd49892,17'd34110,17'd32498,17'd41726,17'd21846,17'd32829,17'd34455,17'd22494,17'd33646,17'd48365,17'd48797,17'd32346,17'd30276,17'd22856,17'd22506,17'd47834,17'd50372,17'd50373,17'd50374,17'd50277,17'd50375,17'd50376,17'd50377,17'd50378,17'd49495,17'd5913,17'd30638,17'd6554,17'd32073,17'd8304,17'd10897,17'd9933,17'd10514,17'd7669,17'd6554,17'd32553,17'd50379,17'd42910,17'd5757,17'd4846,17'd4848,17'd5002,17'd5329,17'd5329,17'd4686,17'd5327,17'd5152,17'd5153,17'd4683,17'd4840,17'd5328,17'd4841,17'd28418,17'd37153,17'd5009,17'd30638,17'd30333,17'd25627,17'd5329,17'd4684,17'd4526,17'd5155,17'd34657,17'd34657,17'd5155,17'd34656,17'd4529,17'd5155,17'd4526,17'd4526,17'd40397,17'd4847,17'd4528,17'd50176,17'd38447,17'd50380,17'd37159,17'd50381,17'd50382,17'd42781,17'd50383,17'd50384,17'd50385,17'd50386,17'd50184,17'd4394,17'd40099,17'd48812,17'd39947,17'd10790,17'd45403,17'd50186,17'd12176,17'd38580,17'd38860,17'd38072,17'd4867,17'd4883,17'd3896,17'd3744,17'd5193,17'd8185,17'd5630,17'd6415,17'd3391,17'd3895,17'd3391,17'd1810,17'd2392,17'd1262,17'd427,17'd607,17'd408,17'd2115,17'd804,17'd50187,17'd403,17'd1092,17'd634
},
'{
17'd3428,17'd3428,17'd10546,17'd3429,17'd31,17'd289,17'd287,17'd652,17'd1278,17'd27,17'd21,17'd21,17'd26,17'd285,17'd50387,17'd7385,17'd980,17'd652,17'd4248,17'd4248,17'd4091,17'd3755,17'd3255,17'd2941,17'd2942,17'd3253,17'd2785,17'd2266,17'd2431,17'd2606,17'd50388,17'd3913,17'd33053,17'd30811,17'd30812,17'd50389,17'd50091,17'd21957,17'd21338,17'd21032,17'd50390,17'd13446,17'd15635,17'd22626,17'd18171,17'd15383,17'd12530,17'd11764,17'd50391,17'd13969,17'd12218,17'd34938,17'd12527,17'd19127,17'd14469,17'd14763,17'd14216,17'd13460,17'd13460,17'd13460,17'd13460,17'd12355,17'd13597,17'd13209,17'd14621,17'd22630,17'd19511,17'd18656,17'd21650,17'd16519,17'd17321,17'd32569,17'd16029,17'd15767,17'd14765,17'd16659,17'd10944,17'd10564,17'd9158,17'd8369,17'd8369,17'd6625,17'd50192,17'd6304,17'd8692,17'd7260,17'd49202,17'd46367,17'd50392,17'd40426,17'd50393,17'd42506,17'd41647,17'd50394,17'd50395,17'd50396,17'd49907,17'd50397,17'd40278,17'd50398,17'd50399,17'd50400,17'd50098,17'd28672,17'd50401,17'd9595,17'd50402,17'd50403,17'd50404,17'd50405,17'd49620,17'd26617,17'd50406,17'd50407,17'd50408,17'd50409,17'd50410,17'd50411,17'd25281,17'd9619,17'd9618,17'd26870,17'd10474,17'd11965,17'd11395,17'd11520,17'd13362,17'd11963,17'd11963,17'd19157,17'd12262,17'd12115,17'd17604,17'd17604,17'd12422,17'd12422,17'd18082,17'd50412,17'd12719,17'd12575,17'd13134,17'd14672,17'd22297,17'd15811,17'd14930,17'd14672,17'd15687,17'd50413,17'd29336,17'd29785,17'd33727,17'd36213,17'd31590,17'd31590,17'd31590,17'd31590,17'd32920,17'd31441,17'd31941,17'd31587,17'd28460,17'd23511,17'd25926,17'd24858,17'd44772,17'd11398,17'd11524,17'd14931,17'd10990,17'd10739,17'd10475,17'd10475,17'd11133,17'd10164,17'd11134,17'd11134,17'd19642,17'd16070,17'd9619,17'd9346,17'd8874,17'd23860,17'd50414,17'd50415,17'd50416,17'd50417,17'd23519,17'd50418,17'd50419,17'd50420,17'd28706,17'd50421,17'd48749,17'd50422,17'd50324,17'd50230,17'd49747,17'd50423,17'd15175,17'd15175,17'd13646,17'd11521,17'd17838,17'd50424,17'd50425,17'd50120,17'd50426,17'd50427,17'd48004,17'd50428,17'd50429,17'd50430,17'd50431,17'd50432,17'd50433,17'd50434,17'd50435,17'd50436,17'd39091,17'd50437,17'd50438,17'd50439,17'd50440,17'd46170,17'd50441,17'd50442,17'd50443,17'd50444,17'd50445,17'd47906,17'd50446,17'd50447,17'd50448,17'd50449,17'd48770,17'd50450,17'd50451,17'd50452,17'd50453,17'd50454,17'd50455,17'd50456,17'd50457,17'd50260,17'd50458,17'd50459,17'd50460,17'd50461,17'd50462,17'd50463,17'd50464,17'd23217,17'd33799,17'd32351,17'd23565,17'd23916,17'd35735,17'd31512,17'd36287,17'd30584,17'd23731,17'd24086,17'd23918,17'd29687,17'd29242,17'd23565,17'd23565,17'd23565,17'd31502,17'd23386,17'd36987,17'd38806,17'd23735,17'd44490,17'd50465,17'd50466,17'd49977,17'd49977,17'd49476,17'd46664,17'd47725,17'd49379,17'd47736,17'd49289,17'd50467,17'd48154,17'd47641,17'd48904,17'd49691,17'd50468,17'd49883,17'd49979,17'd50469,17'd50470,17'd33941,17'd29977,17'd38537,17'd39437,17'd26901,17'd26530,17'd25317,17'd25031,17'd23916,17'd29827,17'd50471,17'd50472,17'd29687,17'd28595,17'd25566,17'd27514,17'd25948,17'd25553,17'd26523,17'd29247,17'd29536,17'd30736,17'd31036,17'd33489,17'd31505,17'd31506,17'd32019,17'd31038,17'd49790,17'd29831,17'd36126,17'd38279,17'd50473,17'd44592,17'd45157,17'd41106,17'd47827,17'd43281,17'd50474,17'd50475,17'd50476,17'd50476,17'd50273,17'd50365,17'd49683,17'd49585,17'd40812,17'd50477,17'd48894,17'd42299,17'd31351,17'd27883,17'd28482,17'd26064,17'd33000,17'd24896,17'd29376,17'd22679,17'd36427,17'd31662,17'd48794,17'd30728,17'd39281,17'd40523,17'd40523,17'd23393,17'd48912,17'd23044,17'd45265,17'd48912,17'd31658,17'd21845,17'd23041,17'd33648,17'd33161,17'd35855,17'd50478,17'd46849,17'd35292,17'd22851,17'd50479,17'd46099,17'd48161,17'd46341,17'd50480,17'd50481,17'd50482,17'd50483,17'd50484,17'd50485,17'd49595,17'd9503,17'd5913,17'd5158,17'd32243,17'd50486,17'd50487,17'd10897,17'd10515,17'd8780,17'd6221,17'd5335,17'd31716,17'd47174,17'd4683,17'd4683,17'd4842,17'd30637,17'd5329,17'd5329,17'd4845,17'd32552,17'd4995,17'd5153,17'd42910,17'd4995,17'd5327,17'd5328,17'd4686,17'd4842,17'd4842,17'd5004,17'd30333,17'd30638,17'd5160,17'd5005,17'd4684,17'd40397,17'd34791,17'd41459,17'd34657,17'd40397,17'd34921,17'd4846,17'd4684,17'd4684,17'd28778,17'd4846,17'd4528,17'd50488,17'd50489,17'd50490,17'd50491,17'd50492,17'd47267,17'd50493,17'd44849,17'd50494,17'd3061,17'd50495,17'd19360,17'd50496,17'd5494,17'd49196,17'd50497,17'd39947,17'd10790,17'd50498,17'd50291,17'd12176,17'd38860,17'd38203,17'd37709,17'd4867,17'd4575,17'd3423,17'd3391,17'd3391,17'd4085,17'd5372,17'd5372,17'd5371,17'd3391,17'd4085,17'd3423,17'd1119,17'd446,17'd623,17'd783,17'd211,17'd1095,17'd186,17'd186,17'd404,17'd593,17'd593
},
'{
17'd3428,17'd3428,17'd10546,17'd2597,17'd30,17'd289,17'd287,17'd28,17'd1278,17'd27,17'd21,17'd21,17'd26,17'd285,17'd21631,17'd7385,17'd27,17'd652,17'd4430,17'd4248,17'd4091,17'd3755,17'd3255,17'd3254,17'd2940,17'd3253,17'd2785,17'd2263,17'd1974,17'd2606,17'd50388,17'd3913,17'd32730,17'd30811,17'd30812,17'd50389,17'd4267,17'd50499,17'd50500,17'd50501,17'd20020,17'd13446,17'd15635,17'd22626,17'd50502,17'd15383,17'd12530,17'd11478,17'd14471,17'd13969,17'd12218,17'd23154,17'd12813,17'd12679,17'd14469,17'd50503,17'd13460,17'd13460,17'd13460,17'd13460,17'd12355,17'd12355,17'd13597,17'd13209,17'd14621,17'd22630,17'd19511,17'd18656,17'd21808,17'd19255,17'd18414,17'd24521,17'd16029,17'd15767,17'd15386,17'd17322,17'd11231,17'd10564,17'd9158,17'd9573,17'd8369,17'd6625,17'd50192,17'd6304,17'd8692,17'd7260,17'd49202,17'd46367,17'd48822,17'd39816,17'd50393,17'd40585,17'd50504,17'd50394,17'd50505,17'd50506,17'd49816,17'd50397,17'd47001,17'd50507,17'd38100,17'd50508,17'd50509,17'd28672,17'd50200,17'd50510,17'd26991,17'd24690,17'd50511,17'd24202,17'd50512,17'd50513,17'd50514,17'd50515,17'd50516,17'd50517,17'd50518,17'd50519,17'd50520,17'd25673,17'd33876,17'd26870,17'd10474,17'd11808,17'd11395,17'd11807,17'd11963,17'd11963,17'd19157,17'd19157,17'd12262,17'd17604,17'd19411,17'd18806,17'd12422,17'd12422,17'd18082,17'd17604,17'd12581,17'd12109,17'd13884,17'd14672,17'd15811,17'd15811,17'd14525,17'd14930,17'd15811,17'd50521,17'd36488,17'd30373,17'd34381,17'd34037,17'd31590,17'd50111,17'd50111,17'd50111,17'd31589,17'd31943,17'd31287,17'd30676,17'd28571,17'd28230,17'd23682,17'd21362,17'd23513,17'd12583,17'd11524,17'd13886,17'd10990,17'd10990,17'd20910,17'd20910,17'd10475,17'd10472,17'd10326,17'd10479,17'd11277,17'd16070,17'd22131,17'd10743,17'd9346,17'd9039,17'd50522,17'd47599,17'd50523,17'd50418,17'd24044,17'd24044,17'd23864,17'd50524,17'd50525,17'd50526,17'd33877,17'd50527,17'd48579,17'd15940,17'd16199,17'd22132,17'd13764,17'd13366,17'd13520,17'd11807,17'd12720,17'd13001,17'd15806,17'd50528,17'd50529,17'd50530,17'd48666,17'd50531,17'd50532,17'd50533,17'd50534,17'd50043,17'd50535,17'd50536,17'd50537,17'd50538,17'd50539,17'd40030,17'd50540,17'd50541,17'd46065,17'd45829,17'd50542,17'd50543,17'd50544,17'd46525,17'd50545,17'd46411,17'd50546,17'd50547,17'd50548,17'd48126,17'd50549,17'd50550,17'd50551,17'd50552,17'd50553,17'd50554,17'd50555,17'd50556,17'd50557,17'd50558,17'd50559,17'd50560,17'd50561,17'd50562,17'd49786,17'd50563,17'd22502,17'd42000,17'd39742,17'd22501,17'd23920,17'd23916,17'd33666,17'd36287,17'd30895,17'd25439,17'd23733,17'd31502,17'd23566,17'd23386,17'd23918,17'd23918,17'd29376,17'd29099,17'd35865,17'd29975,17'd32191,17'd23388,17'd50564,17'd50565,17'd50069,17'd50566,17'd46434,17'd49977,17'd46436,17'd46954,17'd48893,17'd48910,17'd48363,17'd48995,17'd50567,17'd43147,17'd47641,17'd48154,17'd49890,17'd50568,17'd50569,17'd49083,17'd42146,17'd40959,17'd39437,17'd33952,17'd27642,17'd31353,17'd26902,17'd25949,17'd28850,17'd32007,17'd24249,17'd23388,17'd34108,17'd33159,17'd29689,17'd28719,17'd25707,17'd26782,17'd25560,17'd26524,17'd26277,17'd28257,17'd29690,17'd30736,17'd31505,17'd33489,17'd49982,17'd31506,17'd50570,17'd31038,17'd49790,17'd29979,17'd50571,17'd38279,17'd50473,17'd45872,17'd43546,17'd39902,17'd50572,17'd49289,17'd50573,17'd43011,17'd50476,17'd50273,17'd50273,17'd50574,17'd49788,17'd50467,17'd40206,17'd43688,17'd50575,17'd46753,17'd28252,17'd27883,17'd28482,17'd30606,17'd31366,17'd24417,17'd23387,17'd22678,17'd36427,17'd48996,17'd40679,17'd23926,17'd48913,17'd40523,17'd34107,17'd45986,17'd21694,17'd35295,17'd50576,17'd31344,17'd32013,17'd21845,17'd33162,17'd22338,17'd33797,17'd47939,17'd50478,17'd50577,17'd22159,17'd23219,17'd22674,17'd46099,17'd47840,17'd50578,17'd50579,17'd50580,17'd50581,17'd50582,17'd50583,17'd27912,17'd50584,17'd23975,17'd5914,17'd5761,17'd32243,17'd50486,17'd50487,17'd10897,17'd28184,17'd28058,17'd5615,17'd5002,17'd5152,17'd47174,17'd4683,17'd5328,17'd5005,17'd5004,17'd5329,17'd5330,17'd4845,17'd32552,17'd4995,17'd42910,17'd42910,17'd5327,17'd5327,17'd5328,17'd4842,17'd4842,17'd4842,17'd5004,17'd30638,17'd28185,17'd5160,17'd5004,17'd37153,17'd4684,17'd40397,17'd34791,17'd50585,17'd4684,17'd27697,17'd5157,17'd4684,17'd4684,17'd34791,17'd4846,17'd50586,17'd50587,17'd50588,17'd50490,17'd39780,17'd50589,17'd50590,17'd50493,17'd43739,17'd50494,17'd2893,17'd50591,17'd50592,17'd50496,17'd5025,17'd50593,17'd50497,17'd39947,17'd10790,17'd11587,17'd12318,17'd39033,17'd38860,17'd38203,17'd37709,17'd4867,17'd3897,17'd3423,17'd3895,17'd3391,17'd4085,17'd4085,17'd5371,17'd3391,17'd3391,17'd4085,17'd3423,17'd1119,17'd446,17'd623,17'd609,17'd211,17'd1095,17'd639,17'd1682,17'd403,17'd1540,17'd452
},
'{
17'd3428,17'd3251,17'd3752,17'd2597,17'd809,17'd289,17'd287,17'd28,17'd1278,17'd27,17'd285,17'd285,17'd285,17'd285,17'd21631,17'd7385,17'd27,17'd652,17'd4430,17'd4248,17'd4091,17'd4091,17'd3595,17'd3254,17'd2940,17'd3253,17'd2263,17'd2265,17'd2606,17'd2606,17'd50388,17'd3913,17'd32730,17'd30811,17'd30812,17'd50389,17'd50594,17'd50595,17'd21481,17'd50501,17'd20020,17'd13446,17'd17310,17'd20584,17'd50502,17'd19005,17'd12530,17'd11478,17'd13969,17'd13969,17'd12218,17'd11626,17'd12527,17'd14469,17'd14344,17'd13461,17'd13460,17'd13460,17'd13460,17'd13460,17'd12355,17'd12355,17'd14344,17'd13968,17'd13210,17'd13969,17'd25258,17'd18174,17'd21649,17'd21185,17'd22980,17'd24685,17'd14893,17'd15767,17'd14766,17'd16769,17'd16410,17'd10944,17'd9158,17'd9573,17'd8369,17'd6625,17'd6465,17'd6138,17'd8692,17'd7260,17'd49202,17'd6640,17'd46895,17'd6485,17'd40272,17'd40428,17'd50504,17'd41784,17'd50505,17'd50506,17'd44633,17'd50596,17'd50597,17'd50598,17'd38742,17'd37463,17'd50599,17'd30207,17'd27466,17'd9454,17'd50510,17'd50600,17'd50403,17'd9859,17'd50601,17'd26251,17'd50602,17'd50603,17'd50604,17'd50605,17'd9603,17'd50606,17'd50607,17'd50608,17'd9617,17'd26034,17'd10472,17'd16320,17'd11395,17'd11963,17'd11963,17'd11963,17'd19157,17'd15810,17'd12262,17'd12422,17'd18806,17'd12582,17'd12582,17'd12582,17'd17723,17'd12261,17'd17843,17'd12995,17'd16799,17'd14672,17'd15811,17'd22297,17'd14525,17'd14930,17'd15687,17'd50314,17'd37611,17'd31294,17'd30221,17'd31288,17'd31590,17'd35239,17'd50111,17'd50111,17'd31590,17'd34380,17'd31288,17'd30677,17'd29198,17'd28229,17'd24537,17'd23170,17'd23167,17'd11397,17'd11524,17'd11524,17'd10990,17'd10990,17'd10737,17'd10737,17'd10739,17'd10855,17'd10326,17'd11528,17'd11277,17'd14928,17'd14928,17'd17011,17'd9345,17'd24361,17'd17231,17'd28582,17'd8887,17'd19780,17'd8580,17'd8580,17'd8249,17'd9196,17'd35797,17'd23517,17'd50609,17'd33083,17'd16070,17'd20756,17'd15052,17'd15432,17'd13764,17'd13764,17'd11806,17'd11667,17'd16069,17'd13138,17'd26630,17'd28576,17'd15051,17'd28831,17'd50610,17'd50611,17'd50612,17'd50613,17'd50614,17'd50615,17'd50616,17'd50617,17'd50618,17'd50619,17'd50620,17'd50621,17'd50622,17'd50623,17'd50624,17'd50624,17'd40803,17'd50625,17'd50626,17'd50627,17'd50628,17'd50629,17'd50630,17'd50631,17'd50632,17'd50633,17'd50634,17'd50635,17'd50636,17'd50637,17'd50638,17'd50639,17'd50640,17'd50641,17'd50642,17'd50643,17'd50644,17'd50645,17'd50646,17'd50647,17'd50648,17'd39280,17'd36984,17'd50649,17'd22858,17'd23215,17'd31033,17'd29240,17'd24896,17'd25180,17'd34467,17'd29689,17'd29099,17'd35865,17'd23386,17'd23566,17'd23734,17'd29827,17'd30579,17'd31828,17'd29974,17'd32667,17'd23569,17'd29829,17'd23567,17'd50650,17'd49881,17'd49881,17'd50651,17'd50652,17'd46756,17'd39582,17'd50653,17'd40206,17'd48536,17'd49184,17'd48708,17'd43281,17'd48909,17'd49184,17'd50365,17'd50365,17'd50654,17'd50655,17'd46327,17'd32184,17'd27642,17'd29977,17'd36127,17'd30735,17'd28725,17'd27766,17'd27511,17'd28977,17'd24087,17'd23215,17'd32503,17'd50656,17'd30275,17'd27511,17'd31351,17'd27027,17'd27369,17'd27768,17'd28854,17'd28372,17'd29979,17'd31036,17'd31505,17'd33489,17'd49887,17'd33489,17'd30738,17'd30130,17'd49790,17'd36132,17'd50657,17'd38536,17'd47045,17'd38971,17'd41415,17'd50658,17'd46321,17'd49093,17'd50659,17'd50660,17'd50661,17'd50273,17'd50476,17'd50370,17'd49788,17'd49093,17'd39122,17'd42879,17'd46433,17'd43979,17'd25707,17'd26530,17'd26062,17'd30606,17'd33484,17'd23561,17'd29686,17'd34458,17'd32661,17'd48794,17'd31348,17'd48913,17'd48913,17'd32190,17'd32350,17'd32666,17'd32498,17'd32347,17'd32012,17'd31497,17'd21845,17'd31346,17'd32498,17'd32663,17'd42603,17'd42441,17'd48456,17'd45373,17'd22160,17'd22332,17'd32344,17'd32502,17'd38173,17'd50662,17'd50663,17'd50664,17'd50665,17'd50666,17'd50667,17'd50668,17'd50669,17'd6211,17'd50670,17'd28056,17'd26708,17'd8933,17'd9933,17'd27815,17'd8780,17'd6392,17'd5336,17'd28536,17'd47174,17'd42910,17'd4995,17'd4841,17'd5004,17'd25627,17'd5330,17'd5330,17'd4845,17'd4686,17'd4995,17'd42910,17'd5152,17'd5328,17'd4841,17'd28418,17'd4842,17'd4842,17'd4842,17'd5329,17'd5335,17'd28185,17'd5335,17'd5002,17'd4846,17'd4684,17'd40397,17'd34791,17'd28778,17'd4846,17'd42031,17'd4848,17'd4684,17'd40397,17'd34791,17'd4846,17'd50671,17'd49997,17'd50672,17'd50673,17'd50674,17'd37812,17'd3365,17'd21621,17'd44514,17'd50675,17'd38329,17'd50676,17'd50592,17'd50677,17'd7191,17'd50678,17'd50497,17'd39947,17'd10790,17'd50090,17'd44742,17'd38334,17'd37958,17'd38203,17'd37709,17'd4867,17'd3897,17'd3246,17'd3895,17'd3391,17'd4085,17'd4085,17'd3391,17'd3895,17'd3391,17'd3897,17'd3423,17'd228,17'd227,17'd782,17'd3100,17'd2420,17'd253,17'd182,17'd182,17'd805,17'd634,17'd1547
},
'{
17'd3428,17'd3251,17'd3752,17'd2597,17'd809,17'd289,17'd287,17'd28,17'd1278,17'd27,17'd285,17'd285,17'd285,17'd285,17'd21631,17'd7385,17'd27,17'd652,17'd4430,17'd4248,17'd4091,17'd3755,17'd3255,17'd3254,17'd2940,17'd3253,17'd2263,17'd2263,17'd1975,17'd50679,17'd13820,17'd3913,17'd32730,17'd30811,17'd30812,17'd50389,17'd50594,17'd50595,17'd21481,17'd50501,17'd20020,17'd13446,17'd17310,17'd20584,17'd18170,17'd19005,17'd12530,17'd11627,17'd12361,17'd12361,17'd12218,17'd17096,17'd12954,17'd13092,17'd13597,17'd12355,17'd13460,17'd13460,17'd13460,17'd13460,17'd12355,17'd12355,17'd13461,17'd13462,17'd13210,17'd13969,17'd19753,17'd18174,17'd21649,17'd17206,17'd47863,17'd24192,17'd14892,17'd15767,17'd14766,17'd22631,17'd10565,17'd10944,17'd11232,17'd9573,17'd8369,17'd6141,17'd6465,17'd6138,17'd8690,17'd7259,17'd49202,17'd6640,17'd46799,17'd6485,17'd40272,17'd40428,17'd50504,17'd41647,17'd50394,17'd41501,17'd43892,17'd43354,17'd44284,17'd50680,17'd39651,17'd50681,17'd50682,17'd50198,17'd50683,17'd50684,17'd9454,17'd27223,17'd27608,17'd50511,17'd50685,17'd9719,17'd50686,17'd50687,17'd50688,17'd28677,17'd50689,17'd50690,17'd10010,17'd50691,17'd9617,17'd26034,17'd10325,17'd10738,17'd15810,17'd11963,17'd11963,17'd11963,17'd19157,17'd13362,17'd12422,17'd16204,17'd12582,17'd18917,17'd18917,17'd18917,17'd18328,17'd50313,17'd12421,17'd15685,17'd12859,17'd14672,17'd15811,17'd22297,17'd14525,17'd14523,17'd14672,17'd18449,17'd37739,17'd37855,17'd36937,17'd31288,17'd35644,17'd35239,17'd35239,17'd50111,17'd31590,17'd35644,17'd34037,17'd31289,17'd30073,17'd28461,17'd28816,17'd23512,17'd21361,17'd18327,17'd25280,17'd11524,17'd10990,17'd10990,17'd10737,17'd10737,17'd10990,17'd16555,17'd19282,17'd11133,17'd10479,17'd14928,17'd12116,17'd9741,17'd16549,17'd33083,17'd24040,17'd29637,17'd26039,17'd19923,17'd18919,17'd21208,17'd8578,17'd8577,17'd8574,17'd8409,17'd50692,17'd25814,17'd19279,17'd16070,17'd14518,17'd17121,17'd16064,17'd16323,17'd11961,17'd11806,17'd11667,17'd16069,17'd13138,17'd20610,17'd21205,17'd25409,17'd50693,17'd50694,17'd50695,17'd50696,17'd50697,17'd50698,17'd50699,17'd50700,17'd50701,17'd50702,17'd50703,17'd50704,17'd50705,17'd50706,17'd50707,17'd45698,17'd50708,17'd50709,17'd50710,17'd50711,17'd50712,17'd50713,17'd50714,17'd49766,17'd50715,17'd50716,17'd50717,17'd50718,17'd50719,17'd50720,17'd50721,17'd50722,17'd50723,17'd50724,17'd50725,17'd50726,17'd50727,17'd50728,17'd50729,17'd50730,17'd39440,17'd31496,17'd50731,17'd36130,17'd22506,17'd32191,17'd23731,17'd23561,17'd24896,17'd24742,17'd29243,17'd29687,17'd35865,17'd35865,17'd23566,17'd31502,17'd23736,17'd37117,17'd50732,17'd45746,17'd22328,17'd41419,17'd29974,17'd38806,17'd50733,17'd50734,17'd49881,17'd50466,17'd49880,17'd48524,17'd46842,17'd42881,17'd40956,17'd50735,17'd50567,17'd50567,17'd49382,17'd48909,17'd49183,17'd50267,17'd50736,17'd50468,17'd50737,17'd45879,17'd41864,17'd38025,17'd33001,17'd32354,17'd35570,17'd33163,17'd26903,17'd28720,17'd29244,17'd30733,17'd30127,17'd30129,17'd42601,17'd50738,17'd23731,17'd29970,17'd29535,17'd28486,17'd27368,17'd27884,17'd29104,17'd28728,17'd29978,17'd31036,17'd31505,17'd33489,17'd49887,17'd33489,17'd30738,17'd29978,17'd49790,17'd36132,17'd36402,17'd38665,17'd47045,17'd45609,17'd41415,17'd43544,17'd47343,17'd49682,17'd50370,17'd50739,17'd50476,17'd50273,17'd50476,17'd50370,17'd49980,17'd48995,17'd48910,17'd43422,17'd48698,17'd45749,17'd26903,17'd26530,17'd26062,17'd27638,17'd28480,17'd34884,17'd29828,17'd23573,17'd40679,17'd48794,17'd33944,17'd23391,17'd23391,17'd32190,17'd33944,17'd32829,17'd22510,17'd32499,17'd32501,17'd21846,17'd31497,17'd23041,17'd32010,17'd41728,17'd50740,17'd42603,17'd32187,17'd41726,17'd31834,17'd22506,17'd22159,17'd47834,17'd50741,17'd50742,17'd50743,17'd50744,17'd36570,17'd50745,17'd50746,17'd50747,17'd22244,17'd6212,17'd5915,17'd28304,17'd50486,17'd8304,17'd9933,17'd28184,17'd28058,17'd6392,17'd25627,17'd50748,17'd4996,17'd42910,17'd4995,17'd4686,17'd25627,17'd30638,17'd5335,17'd5330,17'd4845,17'd4686,17'd4683,17'd42910,17'd5327,17'd4841,17'd4842,17'd4842,17'd5005,17'd4842,17'd5005,17'd5160,17'd28185,17'd27935,17'd5335,17'd25627,17'd29024,17'd4847,17'd40397,17'd34791,17'd34791,17'd5157,17'd42031,17'd4848,17'd4684,17'd40397,17'd4684,17'd4846,17'd50671,17'd50176,17'd50749,17'd50673,17'd50750,17'd50751,17'd3365,17'd50752,17'd44514,17'd41622,17'd50753,17'd50754,17'd50592,17'd50677,17'd5932,17'd50755,17'd50497,17'd39947,17'd10790,17'd11587,17'd50756,17'd39033,17'd39484,17'd38203,17'd37709,17'd37709,17'd3423,17'd3246,17'd229,17'd3391,17'd4085,17'd4085,17'd3895,17'd3895,17'd3423,17'd3423,17'd3246,17'd228,17'd231,17'd428,17'd429,17'd211,17'd2420,17'd182,17'd181,17'd1091,17'd634,17'd1547
},
'{
17'd3251,17'd3251,17'd10268,17'd2597,17'd809,17'd289,17'd287,17'd27,17'd980,17'd27,17'd286,17'd286,17'd285,17'd467,17'd7555,17'd7385,17'd27,17'd980,17'd4430,17'd4430,17'd4091,17'd4091,17'd3595,17'd3254,17'd2940,17'd2940,17'd2602,17'd2265,17'd2606,17'd50679,17'd50757,17'd4092,17'd32409,17'd30654,17'd3920,17'd50758,17'd50594,17'd22454,17'd50759,17'd23320,17'd20020,17'd50760,17'd17435,17'd19751,17'd50761,17'd19125,17'd12814,17'd11627,17'd12361,17'd12361,17'd14621,17'd13093,17'd13092,17'd14469,17'd14344,17'd12355,17'd13460,17'd13460,17'd13596,17'd13596,17'd13460,17'd14620,17'd13461,17'd13462,17'd13209,17'd14764,17'd32261,17'd25258,17'd17689,17'd19007,17'd19385,17'd22980,17'd14892,17'd15641,17'd14346,17'd16769,17'd16410,17'd10944,17'd9574,17'd7418,17'd8369,17'd6141,17'd5689,17'd5253,17'd5251,17'd7422,17'd6938,17'd50762,17'd46367,17'd49015,17'd39814,17'd39967,17'd40585,17'd50763,17'd50764,17'd50765,17'd45198,17'd43892,17'd50396,17'd50766,17'd50767,17'd50768,17'd50769,17'd8707,17'd50770,17'd50771,17'd50684,17'd27222,17'd27469,17'd50403,17'd21197,17'd50772,17'd50203,17'd50602,17'd50773,17'd50774,17'd50775,17'd50776,17'd34824,17'd35087,17'd9614,17'd9737,17'd50777,17'd33082,17'd18560,17'd13362,17'd28938,17'd11805,17'd11963,17'd11963,17'd16204,17'd16204,17'd18917,17'd18917,17'd18917,17'd18917,17'd12581,17'd12421,17'd50778,17'd50779,17'd12418,17'd12415,17'd15811,17'd24855,17'd21207,17'd14809,17'd14930,17'd15811,17'd50521,17'd38908,17'd29646,17'd31289,17'd34380,17'd35644,17'd35239,17'd35239,17'd35239,17'd35644,17'd35644,17'd33875,17'd34381,17'd30220,17'd28460,17'd25672,17'd23170,17'd16442,17'd11396,17'd11274,17'd11808,17'd11808,17'd10989,17'd10737,17'd10990,17'd11131,17'd11669,17'd19282,17'd11528,17'd10479,17'd9883,17'd9740,17'd11277,17'd19279,17'd34382,17'd16553,17'd23861,17'd8731,17'd9483,17'd14812,17'd21987,17'd24862,17'd8413,17'd8409,17'd29637,17'd16553,17'd16065,17'd22131,17'd17720,17'd10603,17'd16435,17'd15175,17'd11961,17'd11961,17'd11961,17'd13253,17'd11807,17'd14673,17'd11274,17'd33714,17'd50780,17'd50781,17'd50425,17'd50782,17'd50783,17'd50784,17'd50785,17'd50786,17'd50787,17'd50788,17'd50789,17'd50790,17'd50791,17'd50621,17'd50792,17'd50793,17'd50794,17'd50795,17'd50796,17'd50797,17'd50798,17'd50799,17'd46925,17'd50800,17'd50801,17'd50802,17'd50803,17'd50804,17'd50805,17'd50806,17'd50807,17'd50808,17'd50809,17'd50810,17'd50811,17'd50812,17'd50813,17'd50814,17'd50815,17'd45874,17'd22861,17'd50816,17'd50817,17'd50818,17'd22333,17'd23923,17'd29100,17'd23561,17'd24742,17'd29378,17'd48257,17'd30128,17'd23567,17'd23736,17'd29099,17'd30127,17'd23215,17'd23389,17'd45746,17'd22500,17'd32344,17'd22332,17'd29974,17'd24421,17'd50819,17'd50820,17'd49881,17'd49881,17'd50821,17'd48443,17'd41106,17'd49172,17'd47737,17'd48263,17'd50567,17'd48793,17'd43147,17'd43541,17'd50822,17'd49986,17'd50272,17'd49788,17'd48449,17'd44475,17'd41111,17'd30279,17'd33164,17'd32017,17'd36127,17'd27372,17'd25707,17'd27765,17'd27637,17'd33482,17'd29974,17'd42000,17'd50823,17'd33799,17'd23916,17'd33643,17'd27146,17'd28727,17'd47633,17'd28010,17'd28257,17'd29831,17'd30131,17'd31505,17'd31505,17'd33489,17'd31506,17'd33489,17'd30738,17'd29978,17'd49790,17'd31038,17'd50824,17'd41998,17'd46948,17'd44936,17'd39737,17'd43015,17'd47538,17'd49582,17'd42874,17'd43012,17'd50661,17'd50273,17'd50661,17'd50370,17'd49980,17'd48263,17'd41267,17'd42881,17'd50825,17'd44231,17'd27515,17'd26530,17'd26062,17'd28598,17'd27764,17'd28852,17'd37117,17'd36009,17'd50826,17'd31499,17'd32190,17'd47159,17'd45754,17'd32190,17'd32503,17'd31497,17'd22338,17'd32663,17'd33162,17'd31658,17'd31346,17'd33162,17'd22337,17'd33481,17'd41584,17'd48162,17'd50827,17'd44701,17'd22334,17'd46958,17'd45986,17'd50828,17'd50829,17'd50830,17'd50831,17'd50832,17'd36293,17'd50484,17'd19458,17'd50833,17'd47467,17'd5913,17'd5761,17'd28304,17'd50486,17'd50834,17'd9933,17'd8780,17'd28058,17'd27081,17'd4842,17'd30030,17'd4996,17'd42910,17'd5327,17'd5002,17'd5160,17'd28185,17'd5335,17'd5330,17'd4845,17'd4686,17'd5328,17'd5327,17'd5327,17'd4841,17'd4842,17'd5005,17'd5004,17'd30637,17'd5004,17'd5335,17'd28185,17'd27935,17'd5336,17'd25627,17'd4848,17'd37153,17'd4685,17'd37433,17'd37432,17'd5162,17'd5161,17'd29024,17'd4685,17'd4685,17'd4847,17'd50671,17'd50835,17'd50176,17'd50836,17'd50490,17'd50837,17'd48552,17'd50838,17'd44964,17'd44514,17'd20559,17'd50839,17'd50840,17'd2895,17'd50677,17'd50841,17'd50842,17'd50497,17'd39947,17'd10790,17'd50090,17'd11867,17'd38202,17'd39327,17'd38203,17'd37709,17'd3896,17'd3423,17'd3099,17'd3099,17'd3423,17'd3897,17'd3897,17'd3895,17'd3895,17'd3246,17'd3423,17'd50843,17'd4229,17'd3426,17'd447,17'd429,17'd2420,17'd182,17'd182,17'd1822,17'd933,17'd964,17'd454
},
'{
17'd3251,17'd3251,17'd10268,17'd2257,17'd289,17'd653,17'd1833,17'd27,17'd980,17'd27,17'd286,17'd286,17'd285,17'd467,17'd7555,17'd7385,17'd27,17'd980,17'd4430,17'd4430,17'd4091,17'd4091,17'd3595,17'd3254,17'd2941,17'd2940,17'd2602,17'd2264,17'd14600,17'd50679,17'd50757,17'd4092,17'd32409,17'd30654,17'd30348,17'd50758,17'd4749,17'd50844,17'd50759,17'd23146,17'd50845,17'd50760,17'd18403,17'd16876,17'd50761,17'd19125,17'd12814,17'd11627,17'd12361,17'd12361,17'd14621,17'd17096,17'd12954,17'd12678,17'd13597,17'd13461,17'd13460,17'd13460,17'd13596,17'd13596,17'd13460,17'd14620,17'd13461,17'd13597,17'd13209,17'd14764,17'd32261,17'd19753,17'd19893,17'd18774,17'd20149,17'd17690,17'd14892,17'd15641,17'd14346,17'd22631,17'd10565,17'd10428,17'd9159,17'd7418,17'd8369,17'd6142,17'd5837,17'd5253,17'd5087,17'd8070,17'd7420,17'd50762,17'd46367,17'd49015,17'd39814,17'd39967,17'd40585,17'd41332,17'd50846,17'd50847,17'd50096,17'd50097,17'd50506,17'd50848,17'd39350,17'd38609,17'd50849,17'd50850,17'd50851,17'd50852,17'd50684,17'd27110,17'd27223,17'd50853,17'd50854,17'd10001,17'd50855,17'd50686,17'd50856,17'd50857,17'd50858,17'd50859,17'd50860,17'd34954,17'd9872,17'd9737,17'd10161,17'd10601,17'd18445,17'd19157,17'd11805,17'd11805,17'd11962,17'd11963,17'd16204,17'd16204,17'd18917,17'd15053,17'd15053,17'd15053,17'd12719,17'd18558,17'd50861,17'd50862,17'd14003,17'd12415,17'd22297,17'd21057,17'd14526,17'd14809,17'd14525,17'd15811,17'd50521,17'd38908,17'd30373,17'd34381,17'd34037,17'd35644,17'd50863,17'd35239,17'd35239,17'd35239,17'd35239,17'd31590,17'd33568,17'd30221,17'd28686,17'd29778,17'd24031,17'd21363,17'd23167,17'd11396,17'd24029,17'd11808,17'd11965,17'd10989,17'd14931,17'd10854,17'd21206,17'd11132,17'd12863,17'd11528,17'd10479,17'd9883,17'd17719,17'd12116,17'd24037,17'd28815,17'd9194,17'd50864,17'd10607,17'd18201,17'd12586,17'd8413,17'd8413,17'd8572,17'd8569,17'd15684,17'd25814,17'd15298,17'd17839,17'd17720,17'd10604,17'd11395,17'd13253,17'd11961,17'd11961,17'd11961,17'd13520,17'd15185,17'd17478,17'd23337,17'd33714,17'd50865,17'd50866,17'd49439,17'd50867,17'd50868,17'd50869,17'd50870,17'd50871,17'd50872,17'd50873,17'd50874,17'd50875,17'd50876,17'd50877,17'd50878,17'd50879,17'd39234,17'd47026,17'd50880,17'd50341,17'd50799,17'd47027,17'd50881,17'd50882,17'd50883,17'd50884,17'd50885,17'd50886,17'd50887,17'd50888,17'd50889,17'd50890,17'd50891,17'd50892,17'd50893,17'd50894,17'd50895,17'd50896,17'd23222,17'd50818,17'd50897,17'd50898,17'd22494,17'd22860,17'd35865,17'd23732,17'd30879,17'd30275,17'd30278,17'd29973,17'd29974,17'd38806,17'd24421,17'd29099,17'd23387,17'd36426,17'd45874,17'd47457,17'd30427,17'd37659,17'd22860,17'd29974,17'd24421,17'd50899,17'd50900,17'd50901,17'd46434,17'd50902,17'd47049,17'd43690,17'd40509,17'd48363,17'd49390,17'd50567,17'd49382,17'd47736,17'd43419,17'd49891,17'd50736,17'd50272,17'd49479,17'd39735,17'd50903,17'd33791,17'd33164,17'd33321,17'd33654,17'd39437,17'd27372,17'd38538,17'd25709,17'd24898,17'd29375,17'd22331,17'd50904,17'd50905,17'd32504,17'd32007,17'd49273,17'd35011,17'd29379,17'd27761,17'd28371,17'd28857,17'd29978,17'd30280,17'd31837,17'd31505,17'd33489,17'd31506,17'd31506,17'd30280,17'd29978,17'd49790,17'd50906,17'd35989,17'd41998,17'd46948,17'd45039,17'd39902,17'd46845,17'd48909,17'd49988,17'd50907,17'd43146,17'd50661,17'd50476,17'd50661,17'd50574,17'd49683,17'd43147,17'd41579,17'd39582,17'd50908,17'd42147,17'd27515,17'd26530,17'd26064,17'd28597,17'd28974,17'd29378,17'd29973,17'd22858,17'd43985,17'd42601,17'd45492,17'd45379,17'd45754,17'd32190,17'd36427,17'd34455,17'd35295,17'd32011,17'd48912,17'd31658,17'd48912,17'd48457,17'd35855,17'd42151,17'd41112,17'd35710,17'd50909,17'd50910,17'd30728,17'd36566,17'd45986,17'd50911,17'd50912,17'd50913,17'd21712,17'd50914,17'd50915,17'd45772,17'd20086,17'd25994,17'd29022,17'd5914,17'd5761,17'd50916,17'd8933,17'd50487,17'd9933,17'd8780,17'd6221,17'd5336,17'd5152,17'd50917,17'd5153,17'd4995,17'd5328,17'd5329,17'd28185,17'd28185,17'd5335,17'd5160,17'd5002,17'd4686,17'd5328,17'd5327,17'd5328,17'd4842,17'd5005,17'd5005,17'd5004,17'd5004,17'd5004,17'd27935,17'd31717,17'd6554,17'd27935,17'd5160,17'd5008,17'd29024,17'd37153,17'd4685,17'd4685,17'd5161,17'd5162,17'd37153,17'd37153,17'd37153,17'd5157,17'd50671,17'd50918,17'd49997,17'd50919,17'd39020,17'd47264,17'd50920,17'd50921,17'd50922,17'd2536,17'd50923,17'd50924,17'd50840,17'd2895,17'd50925,17'd40715,17'd50842,17'd50497,17'd39947,17'd10790,17'd11587,17'd45291,17'd38859,17'd39484,17'd38203,17'd37709,17'd3896,17'd3246,17'd3099,17'd3099,17'd3423,17'd3897,17'd3423,17'd3895,17'd3246,17'd3246,17'd3246,17'd4712,17'd1825,17'd1264,17'd447,17'd210,17'd211,17'd1682,17'd182,17'd1822,17'd431,17'd962,17'd248
},
'{
17'd3251,17'd14070,17'd2596,17'd2257,17'd289,17'd653,17'd1833,17'd27,17'd980,17'd27,17'd286,17'd286,17'd285,17'd467,17'd7555,17'd7385,17'd27,17'd980,17'd4430,17'd4430,17'd4091,17'd4091,17'd3595,17'd3255,17'd2941,17'd2940,17'd2601,17'd2604,17'd25902,17'd25902,17'd50757,17'd4092,17'd33052,17'd30654,17'd30348,17'd50758,17'd50926,17'd50844,17'd24513,17'd21802,17'd20141,17'd50927,17'd18403,17'd16876,17'd18169,17'd50928,17'd12814,17'd11763,17'd12530,17'd12361,17'd14621,17'd13093,17'd12678,17'd12357,17'd14344,17'd13461,17'd13460,17'd13460,17'd13595,17'd13595,17'd13596,17'd13837,17'd13460,17'd14344,17'd13209,17'd14621,17'd50391,17'd20423,17'd19006,17'd19128,17'd28668,17'd19385,17'd16987,17'd14892,17'd14346,17'd15899,17'd16410,17'd10944,17'd15517,17'd7418,17'd9573,17'd8368,17'd6141,17'd5254,17'd6627,17'd8690,17'd7099,17'd50929,17'd50930,17'd46895,17'd50392,17'd39816,17'd50931,17'd50932,17'd50933,17'd50846,17'd42216,17'd41648,17'd50934,17'd50935,17'd50767,17'd38609,17'd50936,17'd50937,17'd50938,17'd50939,17'd50940,17'd27109,17'd27222,17'd9595,17'd50853,17'd50941,17'd49725,17'd50942,17'd50943,17'd50944,17'd50945,17'd50946,17'd30966,17'd50947,17'd50948,17'd50949,17'd10161,17'd10601,17'd42810,17'd19157,17'd16797,17'd16797,17'd11805,17'd28938,17'd18447,17'd18447,17'd12260,17'd12858,17'd11958,17'd12420,17'd12106,17'd17603,17'd50950,17'd50862,17'd13515,17'd12416,17'd24855,17'd21207,17'd14526,17'd14526,17'd14525,17'd15811,17'd16556,17'd35101,17'd36347,17'd29785,17'd31289,17'd34037,17'd35644,17'd35239,17'd50951,17'd50952,17'd50952,17'd35239,17'd33875,17'd34835,17'd31587,17'd29480,17'd25672,17'd22819,17'd21361,17'd16326,17'd11397,17'd24029,17'd11808,17'd11274,17'd11274,17'd11808,17'd10854,17'd11132,17'd12863,17'd11527,17'd11133,17'd10326,17'd10166,17'd17719,17'd9739,17'd33722,17'd15569,17'd16553,17'd9040,17'd8410,17'd30969,17'd11404,17'd8572,17'd8730,17'd8724,17'd9621,17'd10174,17'd16065,17'd15048,17'd25675,17'd19156,17'd10852,17'd11395,17'd11667,17'd20313,17'd20313,17'd11806,17'd13135,17'd13520,17'd14264,17'd17343,17'd24035,17'd31130,17'd50953,17'd50954,17'd50955,17'd50956,17'd50957,17'd50958,17'd50959,17'd50960,17'd50961,17'd50962,17'd50963,17'd50964,17'd50965,17'd50966,17'd50967,17'd50968,17'd50969,17'd50342,17'd46524,17'd50546,17'd45594,17'd50970,17'd50971,17'd50972,17'd50973,17'd50974,17'd50975,17'd50976,17'd50977,17'd50978,17'd50979,17'd50980,17'd50981,17'd50982,17'd50983,17'd50984,17'd42441,17'd50985,17'd50986,17'd47066,17'd50987,17'd47457,17'd31655,17'd31502,17'd29099,17'd23217,17'd32830,17'd36986,17'd39440,17'd40960,17'd31502,17'd50988,17'd50989,17'd50990,17'd50991,17'd38172,17'd45876,17'd31496,17'd22330,17'd37511,17'd50733,17'd50992,17'd50993,17'd50266,17'd46662,17'd50994,17'd50995,17'd42596,17'd49574,17'd49390,17'd49485,17'd50567,17'd49979,17'd48909,17'd49289,17'd49985,17'd50272,17'd50996,17'd41098,17'd44473,17'd46425,17'd27642,17'd32193,17'd33486,17'd33654,17'd31353,17'd27146,17'd25708,17'd28717,17'd24898,17'd29528,17'd22159,17'd50997,17'd50998,17'd29376,17'd41730,17'd27260,17'd37908,17'd29977,17'd28981,17'd29537,17'd29690,17'd30280,17'd31506,17'd31837,17'd31036,17'd30280,17'd31505,17'd30736,17'd30738,17'd29979,17'd29979,17'd50906,17'd35989,17'd41998,17'd44592,17'd44101,17'd50658,17'd41414,17'd48263,17'd49794,17'd50907,17'd43146,17'd50661,17'd50661,17'd50273,17'd50574,17'd49691,17'd47736,17'd42295,17'd47052,17'd42300,17'd31351,17'd27514,17'd26062,17'd28594,17'd25709,17'd23561,17'd23385,17'd39131,17'd35296,17'd50826,17'd31348,17'd31500,17'd24094,17'd44591,17'd23926,17'd49094,17'd31659,17'd32347,17'd22511,17'd31831,17'd31192,17'd31660,17'd32011,17'd35154,17'd42152,17'd50999,17'd35155,17'd51000,17'd51001,17'd23393,17'd51002,17'd51003,17'd50168,17'd51004,17'd51005,17'd51006,17'd51007,17'd51008,17'd51009,17'd20836,17'd26582,17'd7494,17'd50670,17'd6389,17'd26708,17'd8933,17'd50487,17'd8780,17'd28058,17'd26828,17'd5002,17'd29594,17'd47471,17'd5153,17'd4995,17'd4841,17'd5330,17'd28185,17'd28185,17'd5335,17'd5160,17'd5002,17'd4842,17'd5328,17'd5327,17'd28418,17'd4842,17'd5005,17'd5004,17'd25627,17'd25627,17'd25627,17'd5336,17'd28185,17'd6554,17'd27935,17'd5335,17'd5004,17'd30637,17'd37029,17'd37288,17'd37029,17'd5167,17'd5009,17'd37288,17'd29024,17'd4848,17'd5161,17'd5006,17'd49996,17'd51010,17'd51011,17'd51012,17'd48805,17'd51013,17'd44848,17'd51014,17'd51015,17'd51016,17'd51017,17'd40097,17'd51018,17'd51019,17'd50184,17'd50842,17'd50497,17'd39947,17'd10790,17'd39032,17'd11867,17'd39948,17'd39327,17'd37709,17'd3423,17'd3423,17'd3246,17'd3099,17'd2586,17'd3247,17'd3423,17'd3423,17'd2586,17'd2586,17'd2586,17'd50843,17'd3898,17'd3426,17'd1264,17'd447,17'd210,17'd2420,17'd639,17'd182,17'd2251,17'd2251,17'd432,17'd51020
},
'{
17'd3251,17'd14070,17'd2596,17'd1414,17'd289,17'd653,17'd1833,17'd27,17'd980,17'd27,17'd286,17'd286,17'd285,17'd467,17'd7555,17'd7385,17'd27,17'd980,17'd4430,17'd4430,17'd4431,17'd4091,17'd3595,17'd3255,17'd2941,17'd2940,17'd2601,17'd2601,17'd2945,17'd25902,17'd50757,17'd4092,17'd33052,17'd30654,17'd30348,17'd50758,17'd50926,17'd51021,17'd12342,17'd13194,17'd13700,17'd50927,17'd18403,17'd16876,17'd18169,17'd50928,17'd12814,17'd11627,17'd12361,17'd12361,17'd14621,17'd23325,17'd12812,17'd12678,17'd13597,17'd13461,17'd13460,17'd13460,17'd13595,17'd13595,17'd13596,17'd13837,17'd13460,17'd14344,17'd13092,17'd13211,17'd14471,17'd20423,17'd18884,17'd19382,17'd19511,17'd19008,17'd16987,17'd14768,17'd14219,17'd15899,17'd16410,17'd10428,17'd9300,17'd7418,17'd9573,17'd8368,17'd6141,17'd5254,17'd6627,17'd8541,17'd7421,17'd40873,17'd46489,17'd46895,17'd50392,17'd39816,17'd39649,17'd6646,17'd50932,17'd41332,17'd51022,17'd51023,17'd50934,17'd50935,17'd50767,17'd51024,17'd51025,17'd35922,17'd50938,17'd51026,17'd51027,17'd51028,17'd27110,17'd27223,17'd51029,17'd51030,17'd51031,17'd50203,17'd50602,17'd51032,17'd51033,17'd51034,17'd51035,17'd51036,17'd51037,17'd9733,17'd10020,17'd50777,17'd51038,17'd11665,17'd16198,17'd16797,17'd11805,17'd28938,17'd18447,17'd18447,17'd12260,17'd12858,17'd12420,17'd12419,17'd12106,17'd17603,17'd50862,17'd15433,17'd13515,17'd14003,17'd24855,17'd21207,17'd51039,17'd45548,17'd15942,17'd21057,17'd21504,17'd51040,17'd39070,17'd29481,17'd30677,17'd34203,17'd35644,17'd35239,17'd35239,17'd50952,17'd50952,17'd50863,17'd34545,17'd34203,17'd30676,17'd31286,17'd27346,17'd23512,17'd21363,17'd18443,17'd18327,17'd24029,17'd11275,17'd11274,17'd14673,17'd11274,17'd10990,17'd10854,17'd10476,17'd12863,17'd10326,17'd10326,17'd10165,17'd10165,17'd9883,17'd17839,17'd48849,17'd9344,17'd9189,17'd29637,17'd9348,17'd8410,17'd24368,17'd33404,17'd9195,17'd8880,17'd9042,17'd24361,17'd16065,17'd33722,17'd45549,17'd29332,17'd14931,17'd11395,17'd16064,17'd20313,17'd20313,17'd11806,17'd13646,17'd13646,17'd11521,17'd13000,17'd17121,17'd22296,17'd51041,17'd51042,17'd50222,17'd51043,17'd51044,17'd51045,17'd51046,17'd51047,17'd43773,17'd51048,17'd51049,17'd50964,17'd51050,17'd50966,17'd46626,17'd49962,17'd50049,17'd46525,17'd51051,17'd51052,17'd51053,17'd51054,17'd51055,17'd51056,17'd51057,17'd51058,17'd51059,17'd51060,17'd51061,17'd22016,17'd51062,17'd51063,17'd51064,17'd51065,17'd51066,17'd51067,17'd51068,17'd51069,17'd22154,17'd51070,17'd51071,17'd37116,17'd32351,17'd30425,17'd31656,17'd34458,17'd22328,17'd31828,17'd40960,17'd23736,17'd40833,17'd35736,17'd34638,17'd51072,17'd51073,17'd50576,17'd32344,17'd22329,17'd31828,17'd51074,17'd50900,17'd50651,17'd51075,17'd46757,17'd49572,17'd51076,17'd46846,17'd50735,17'd51077,17'd49693,17'd50567,17'd48154,17'd48264,17'd49484,17'd50072,17'd50371,17'd51078,17'd51079,17'd44102,17'd32994,17'd40371,17'd33486,17'd29107,17'd28134,17'd29245,17'd28725,17'd28602,17'd28480,17'd25032,17'd33794,17'd22683,17'd51080,17'd23740,17'd30431,17'd43022,17'd32006,17'd39437,17'd33001,17'd29105,17'd29831,17'd49579,17'd33489,17'd31506,17'd31837,17'd31036,17'd30280,17'd31505,17'd31506,17'd30736,17'd29979,17'd29979,17'd50906,17'd35989,17'd51081,17'd44592,17'd46844,17'd51082,17'd46955,17'd49184,17'd49890,17'd50739,17'd43146,17'd50661,17'd50661,17'd50907,17'd49986,17'd49682,17'd47641,17'd42595,17'd46665,17'd46753,17'd25707,17'd27514,17'd26062,17'd28130,17'd25178,17'd24090,17'd29830,17'd34458,17'd35429,17'd43840,17'd30881,17'd51083,17'd24094,17'd40523,17'd30728,17'd47346,17'd33648,17'd32499,17'd22510,17'd31831,17'd31345,17'd32662,17'd32187,17'd42747,17'd51084,17'd51085,17'd35015,17'd22671,17'd51086,17'd36289,17'd51087,17'd44000,17'd45374,17'd47353,17'd51088,17'd51089,17'd51090,17'd51091,17'd24780,17'd21299,17'd12884,17'd6844,17'd5761,17'd6389,17'd51092,17'd51093,17'd50487,17'd8780,17'd28058,17'd26949,17'd4841,17'd47471,17'd47471,17'd42910,17'd5327,17'd4842,17'd5335,17'd28185,17'd31717,17'd28185,17'd5160,17'd5002,17'd28418,17'd5328,17'd5327,17'd4842,17'd5005,17'd30637,17'd5004,17'd5160,17'd5160,17'd25627,17'd27935,17'd31717,17'd6390,17'd5614,17'd28185,17'd25627,17'd5004,17'd5008,17'd37029,17'd5009,17'd5168,17'd5009,17'd37029,17'd5008,17'd4848,17'd42031,17'd5006,17'd50587,17'd51010,17'd51011,17'd51094,17'd51095,17'd51013,17'd44739,17'd51014,17'd2727,17'd39027,17'd51096,17'd40097,17'd51097,17'd50925,17'd50184,17'd8481,17'd4225,17'd39947,17'd10790,17'd11188,17'd51098,17'd39483,17'd39484,17'd38203,17'd37821,17'd3423,17'd3246,17'd3099,17'd2586,17'd3247,17'd3423,17'd3246,17'd3247,17'd2586,17'd50843,17'd4712,17'd3898,17'd795,17'd447,17'd226,17'd1094,17'd211,17'd186,17'd964,17'd2251,17'd27948,17'd455,17'd51099
},
'{
17'd14188,17'd2422,17'd2596,17'd1414,17'd289,17'd652,17'd27,17'd286,17'd26,17'd26,17'd286,17'd286,17'd467,17'd467,17'd7555,17'd7555,17'd27,17'd980,17'd4430,17'd4430,17'd4091,17'd4091,17'd3907,17'd3595,17'd3254,17'd2941,17'd2601,17'd2604,17'd25902,17'd13819,17'd4432,17'd3912,17'd33052,17'd31259,17'd30348,17'd50758,17'd23492,17'd50844,17'd24513,17'd21802,17'd20418,17'd50927,17'd16155,17'd19750,17'd17935,17'd32896,17'd12955,17'd12065,17'd12530,17'd12362,17'd13211,17'd13093,17'd12678,17'd12062,17'd12355,17'd12355,17'd13460,17'd13460,17'd13595,17'd13595,17'd12212,17'd12212,17'd13460,17'd13461,17'd13597,17'd13210,17'd13969,17'd12681,17'd12532,17'd18884,17'd19892,17'd25512,17'd18776,17'd16987,17'd16033,17'd15899,17'd16410,17'd10945,17'd15517,17'd7418,17'd9573,17'd7087,17'd6468,17'd5689,17'd6306,17'd8690,17'd8375,17'd51100,17'd6635,17'd46999,17'd51101,17'd6485,17'd38891,17'd6788,17'd51102,17'd50933,17'd51103,17'd51104,17'd50765,17'd51105,17'd51106,17'd51024,17'd51107,17'd51108,17'd33394,17'd51026,17'd50940,17'd51028,17'd27331,17'd50510,17'd26991,17'd51109,17'd51110,17'd51111,17'd51112,17'd17336,17'd51113,17'd51114,17'd51115,17'd10452,17'd51116,17'd10313,17'd50949,17'd50777,17'd10470,17'd25278,17'd11665,17'd21982,17'd11805,17'd11805,17'd28938,17'd21822,17'd19412,17'd11957,17'd12857,17'd11958,17'd16321,17'd16321,17'd15433,17'd15433,17'd34558,17'd13515,17'd14003,17'd13515,17'd14526,17'd45548,17'd50862,17'd34558,17'd14003,17'd16556,17'd35101,17'd51117,17'd29785,17'd34381,17'd34037,17'd51118,17'd50863,17'd35239,17'd50951,17'd50863,17'd51118,17'd34037,17'd31941,17'd31587,17'd28345,17'd25927,17'd24209,17'd21361,17'd18327,17'd11397,17'd11808,17'd11808,17'd14931,17'd14931,17'd10737,17'd14931,17'd13886,17'd10476,17'd11132,17'd19282,17'd19532,17'd10326,17'd10165,17'd9883,17'd20756,17'd15048,17'd15187,17'd10174,17'd15684,17'd9195,17'd8729,17'd8729,17'd26154,17'd16317,17'd10336,17'd8874,17'd9344,17'd17011,17'd29199,17'd16908,17'd10603,17'd10738,17'd10737,17'd16064,17'd28108,17'd13764,17'd13253,17'd13253,17'd11667,17'd11520,17'd12720,17'd17715,17'd51119,17'd32123,17'd51120,17'd51121,17'd50320,17'd51122,17'd51123,17'd51124,17'd51125,17'd51126,17'd51127,17'd51128,17'd45856,17'd51129,17'd47122,17'd51130,17'd51131,17'd50246,17'd51132,17'd51133,17'd51134,17'd51135,17'd51136,17'd51137,17'd51138,17'd51139,17'd51140,17'd51141,17'd51142,17'd51143,17'd51144,17'd51145,17'd51146,17'd47067,17'd51147,17'd51148,17'd51149,17'd51150,17'd48716,17'd51151,17'd51152,17'd22504,17'd22858,17'd36009,17'd22858,17'd22331,17'd23388,17'd34112,17'd41587,17'd22503,17'd44360,17'd49094,17'd47949,17'd32348,17'd51153,17'd32997,17'd36566,17'd23570,17'd34894,17'd50899,17'd51154,17'd51075,17'd50821,17'd47436,17'd51155,17'd48707,17'd49586,17'd48995,17'd51156,17'd49987,17'd49093,17'd43281,17'd48363,17'd49691,17'd51157,17'd50160,17'd51158,17'd51159,17'd44477,17'd37908,17'd32192,17'd32018,17'd37250,17'd30279,17'd28486,17'd28725,17'd30734,17'd28480,17'd25032,17'd51160,17'd49096,17'd46322,17'd32191,17'd32668,17'd28253,17'd34637,17'd27884,17'd28855,17'd29106,17'd29979,17'd33323,17'd33489,17'd31505,17'd31837,17'd31036,17'd30280,17'd33489,17'd33489,17'd30280,17'd29978,17'd29981,17'd51161,17'd35705,17'd51081,17'd45872,17'd44474,17'd51162,17'd43830,17'd49583,17'd50574,17'd50661,17'd43146,17'd51163,17'd50661,17'd50476,17'd49985,17'd49390,17'd47343,17'd42738,17'd47925,17'd45749,17'd27515,17'd26062,17'd30606,17'd25317,17'd25030,17'd28849,17'd29828,17'd23038,17'd35711,17'd42601,17'd34278,17'd31663,17'd45379,17'd23391,17'd32346,17'd49588,17'd33796,17'd32664,17'd22864,17'd41726,17'd31660,17'd32010,17'd48162,17'd51164,17'd51084,17'd46217,17'd48456,17'd51165,17'd51166,17'd36427,17'd51167,17'd51168,17'd51169,17'd51170,17'd51171,17'd51172,17'd51173,17'd51174,17'd47757,17'd25219,17'd8913,17'd5914,17'd5331,17'd6389,17'd8303,17'd8780,17'd8780,17'd6220,17'd27081,17'd33692,17'd30485,17'd38317,17'd38442,17'd4996,17'd5327,17'd5002,17'd5335,17'd27935,17'd6554,17'd28185,17'd5160,17'd5002,17'd4842,17'd5328,17'd5328,17'd28536,17'd4842,17'd5004,17'd25627,17'd30333,17'd30638,17'd30638,17'd28185,17'd6554,17'd6390,17'd5614,17'd27935,17'd5160,17'd5004,17'd5004,17'd5004,17'd37030,17'd5165,17'd51175,17'd37029,17'd38059,17'd5011,17'd4849,17'd51176,17'd50587,17'd51177,17'd51178,17'd50674,17'd51179,17'd51180,17'd45782,17'd51181,17'd51182,17'd50924,17'd51096,17'd40560,17'd51018,17'd50677,17'd51183,17'd41000,17'd4225,17'd39947,17'd45186,17'd39032,17'd11048,17'd38202,17'd37957,17'd37821,17'd3423,17'd3246,17'd1119,17'd228,17'd1119,17'd2586,17'd2586,17'd2586,17'd50843,17'd50843,17'd5195,17'd3898,17'd4398,17'd4398,17'd2587,17'd234,17'd244,17'd212,17'd963,17'd1822,17'd462,17'd931,17'd613,17'd51184
},
'{
17'd14188,17'd2422,17'd2596,17'd1414,17'd289,17'd652,17'd27,17'd286,17'd26,17'd26,17'd286,17'd1833,17'd467,17'd467,17'd7555,17'd7555,17'd286,17'd980,17'd4430,17'd4430,17'd4091,17'd4091,17'd3907,17'd3595,17'd3254,17'd2941,17'd3105,17'd2601,17'd3106,17'd13187,17'd4432,17'd3912,17'd33052,17'd31259,17'd30348,17'd50758,17'd23492,17'd6609,17'd22974,17'd13194,17'd13700,17'd50927,17'd16155,17'd18166,17'd17935,17'd32896,17'd12955,17'd12065,17'd12218,17'd12362,17'd13211,17'd13093,17'd12678,17'd12062,17'd13461,17'd12355,17'd13460,17'd13460,17'd13595,17'd13595,17'd12212,17'd12212,17'd13460,17'd12355,17'd13597,17'd13210,17'd13969,17'd12681,17'd12532,17'd12532,17'd19382,17'd27461,17'd18776,17'd16290,17'd16033,17'd15899,17'd16410,17'd10945,17'd10429,17'd7418,17'd9573,17'd6769,17'd5409,17'd5689,17'd6306,17'd8541,17'd43069,17'd51100,17'd6635,17'd46999,17'd51101,17'd6485,17'd38891,17'd38482,17'd51185,17'd50932,17'd51186,17'd50847,17'd50765,17'd51105,17'd51106,17'd50767,17'd38609,17'd37060,17'd51187,17'd51188,17'd51189,17'd27605,17'd27331,17'd27110,17'd50510,17'd50402,17'd26861,17'd51190,17'd51191,17'd51192,17'd51193,17'd51194,17'd51195,17'd30521,17'd10589,17'd51196,17'd50949,17'd50777,17'd10324,17'd26869,17'd32590,17'd21982,17'd28812,17'd11805,17'd28938,17'd16548,17'd16548,17'd11957,17'd12857,17'd11958,17'd16321,17'd16321,17'd15433,17'd15433,17'd48846,17'd13515,17'd14003,17'd13517,17'd21506,17'd45548,17'd50862,17'd15433,17'd13515,17'd21504,17'd16557,17'd37206,17'd29201,17'd36937,17'd34203,17'd34380,17'd51118,17'd50863,17'd50952,17'd50952,17'd50863,17'd35644,17'd31287,17'd30676,17'd28461,17'd28103,17'd24030,17'd21363,17'd23513,17'd18327,17'd11397,17'd11808,17'd11274,17'd14931,17'd10737,17'd10737,17'd10990,17'd10476,17'd11132,17'd19282,17'd19282,17'd19532,17'd10165,17'd10165,17'd11670,17'd10479,17'd15048,17'd9345,17'd10174,17'd15684,17'd25677,17'd26259,17'd38904,17'd16440,17'd17480,17'd17480,17'd10173,17'd15187,17'd15048,17'd25675,17'd22296,17'd10603,17'd16320,17'd10736,17'd29331,17'd13885,17'd13885,17'd16064,17'd11667,17'd13137,17'd15182,17'd13001,17'd21205,17'd33237,17'd25408,17'd17347,17'd51197,17'd51121,17'd51198,17'd51199,17'd51200,17'd51201,17'd51202,17'd51203,17'd51204,17'd46304,17'd44462,17'd51205,17'd51206,17'd51207,17'd51208,17'd51209,17'd51210,17'd51211,17'd51212,17'd51213,17'd51214,17'd51215,17'd51216,17'd51217,17'd51218,17'd51219,17'd51219,17'd51220,17'd51221,17'd51222,17'd51223,17'd51224,17'd51225,17'd51226,17'd51227,17'd51228,17'd51151,17'd30580,17'd32345,17'd31657,17'd36009,17'd51229,17'd35865,17'd23736,17'd22680,17'd37510,17'd21845,17'd32662,17'd51230,17'd51231,17'd33647,17'd32997,17'd32350,17'd43843,17'd51232,17'd51233,17'd51154,17'd50263,17'd51234,17'd49473,17'd48047,17'd48049,17'd48154,17'd49682,17'd49984,17'd49891,17'd48995,17'd43419,17'd49093,17'd49575,17'd50160,17'd49787,17'd48450,17'd49079,17'd45878,17'd30279,17'd32507,17'd36989,17'd33320,17'd31503,17'd26901,17'd26903,17'd30734,17'd27511,17'd28851,17'd38806,17'd22861,17'd37249,17'd30127,17'd39443,17'd28252,17'd37908,17'd28133,17'd28856,17'd29536,17'd30131,17'd33323,17'd33488,17'd31505,17'd31837,17'd31036,17'd30280,17'd33323,17'd33489,17'd30131,17'd29979,17'd29833,17'd51235,17'd35705,17'd45747,17'd38971,17'd43545,17'd40047,17'd39575,17'd49692,17'd50907,17'd51236,17'd43146,17'd51163,17'd50476,17'd50072,17'd49987,17'd49289,17'd48700,17'd43832,17'd48145,17'd32995,17'd27514,17'd26062,17'd28720,17'd27511,17'd24416,17'd29242,17'd23216,17'd23573,17'd35711,17'd39282,17'd32015,17'd44110,17'd34453,17'd39281,17'd48911,17'd49588,17'd31832,17'd34456,17'd51237,17'd41726,17'd32662,17'd35015,17'd35154,17'd51238,17'd46456,17'd51239,17'd49795,17'd22848,17'd51086,17'd48911,17'd37534,17'd51240,17'd51241,17'd51242,17'd51243,17'd51244,17'd51245,17'd26097,17'd51246,17'd25622,17'd7166,17'd5915,17'd26218,17'd26708,17'd8933,17'd7668,17'd8780,17'd6391,17'd26828,17'd4686,17'd38058,17'd38441,17'd4991,17'd5145,17'd5328,17'd5329,17'd28185,17'd6554,17'd6554,17'd28185,17'd30638,17'd5004,17'd4842,17'd5328,17'd5328,17'd28418,17'd4842,17'd5004,17'd25627,17'd30638,17'd30638,17'd30638,17'd28185,17'd6554,17'd6390,17'd5614,17'd27935,17'd30638,17'd5004,17'd5004,17'd25627,17'd37030,17'd5165,17'd51175,17'd51175,17'd38059,17'd5011,17'd4849,17'd51247,17'd51248,17'd4372,17'd51249,17'd50750,17'd51179,17'd51180,17'd20859,17'd51250,17'd2540,17'd51096,17'd2900,17'd40560,17'd51018,17'd51251,17'd51252,17'd41000,17'd4225,17'd39947,17'd45186,17'd40716,17'd51253,17'd38859,17'd38334,17'd37957,17'd37821,17'd3246,17'd228,17'd228,17'd1119,17'd2586,17'd2586,17'd2586,17'd50843,17'd50843,17'd5195,17'd1824,17'd4398,17'd1120,17'd226,17'd234,17'd633,17'd246,17'd212,17'd964,17'd441,17'd1238,17'd18515,17'd51254
},
'{
17'd14188,17'd1831,17'd1414,17'd1416,17'd653,17'd652,17'd286,17'd286,17'd26,17'd26,17'd285,17'd467,17'd467,17'd467,17'd7555,17'd7385,17'd286,17'd980,17'd4430,17'd4430,17'd4091,17'd4091,17'd3907,17'd3595,17'd3255,17'd2941,17'd3105,17'd4739,17'd5805,17'd14192,17'd5219,17'd5217,17'd32088,17'd31259,17'd30348,17'd29043,17'd23492,17'd22619,17'd23829,17'd51255,17'd21644,17'd12797,17'd15756,17'd18166,17'd16762,17'd17571,17'd12679,17'd12065,17'd12218,17'd13094,17'd12955,17'd13093,17'd12678,17'd12357,17'd13461,17'd13461,17'd13460,17'd13460,17'd13595,17'd13595,17'd12212,17'd12212,17'd13596,17'd13838,17'd12356,17'd13599,17'd12530,17'd11764,17'd12361,17'd16765,17'd19006,17'd18655,17'd16519,17'd15902,17'd16034,17'd20585,17'd17318,17'd10945,17'd10429,17'd7418,17'd9573,17'd9701,17'd7418,17'd5255,17'd7252,17'd5251,17'd5085,17'd7097,17'd6637,17'd46489,17'd51256,17'd49015,17'd39504,17'd38482,17'd38603,17'd6646,17'd41783,17'd51103,17'd50847,17'd51105,17'd51257,17'd51258,17'd51259,17'd51260,17'd51261,17'd8861,17'd51262,17'd29460,17'd51263,17'd27110,17'd9454,17'd51264,17'd50011,17'd50405,17'd51265,17'd18434,17'd51266,17'd15931,17'd51267,17'd10586,17'd10588,17'd51268,17'd9734,17'd10161,17'd32777,17'd51269,17'd51270,17'd32590,17'd16313,17'd11804,17'd11956,17'd37741,17'd37741,17'd29492,17'd47110,17'd12998,17'd13136,17'd13252,17'd15433,17'd51271,17'd48846,17'd13515,17'd12417,17'd13517,17'd15685,17'd50779,17'd50779,17'd15685,17'd17348,17'd19407,17'd23855,17'd27121,17'd28460,17'd28686,17'd30221,17'd31288,17'd51118,17'd50863,17'd50952,17'd50952,17'd51272,17'd51118,17'd31288,17'd34381,17'd29198,17'd28818,17'd24856,17'd24992,17'd24706,17'd23513,17'd11397,17'd11808,17'd11808,17'd11274,17'd10737,17'd10737,17'd10737,17'd10990,17'd10854,17'd11131,17'd11132,17'd19282,17'd19532,17'd19532,17'd24996,17'd12863,17'd11528,17'd12116,17'd9345,17'd24361,17'd23859,17'd16317,17'd17607,17'd16440,17'd17480,17'd26153,17'd10335,17'd9344,17'd10742,17'd9740,17'd29199,17'd25928,17'd10477,17'd10739,17'd16320,17'd51273,17'd16792,17'd15432,17'd16068,17'd13000,17'd16068,17'd14931,17'd17838,17'd26630,17'd26759,17'd18080,17'd17346,17'd51274,17'd51275,17'd49239,17'd51276,17'd51277,17'd51278,17'd51279,17'd51280,17'd51281,17'd51282,17'd51283,17'd51284,17'd51285,17'd51286,17'd51287,17'd51288,17'd51289,17'd51290,17'd51291,17'd51292,17'd51293,17'd51294,17'd51295,17'd51296,17'd51297,17'd51295,17'd51298,17'd51299,17'd51300,17'd51300,17'd51301,17'd46679,17'd51302,17'd48161,17'd31830,17'd22005,17'd22167,17'd22165,17'd31657,17'd22679,17'd41587,17'd34894,17'd30277,17'd31031,17'd41726,17'd21853,17'd51303,17'd51304,17'd51305,17'd51302,17'd31346,17'd51306,17'd37116,17'd51307,17'd51308,17'd51309,17'd51310,17'd51311,17'd51312,17'd51313,17'd47737,17'd48708,17'd50267,17'd49987,17'd49891,17'd49289,17'd48995,17'd49691,17'd49980,17'd49980,17'd48793,17'd48040,17'd46660,17'd36542,17'd28134,17'd36989,17'd32018,17'd39910,17'd31352,17'd26902,17'd25833,17'd28598,17'd31034,17'd34467,17'd29829,17'd37659,17'd51314,17'd50364,17'd28721,17'd27258,17'd32356,17'd28256,17'd30587,17'd36132,17'd30280,17'd33489,17'd33488,17'd31505,17'd31036,17'd30738,17'd30130,17'd30131,17'd33489,17'd30131,17'd29979,17'd30434,17'd51235,17'd51315,17'd40519,17'd44828,17'd43153,17'd45478,17'd49289,17'd49987,17'd50273,17'd51236,17'd51236,17'd51163,17'd50476,17'd49986,17'd49988,17'd43419,17'd45151,17'd49696,17'd49474,17'd28252,17'd26530,17'd28602,17'd28484,17'd27637,17'd28975,17'd29826,17'd30425,17'd36009,17'd35711,17'd35736,17'd23570,17'd33511,17'd34453,17'd31834,17'd47346,17'd31659,17'd33798,17'd35295,17'd51316,17'd32997,17'd32010,17'd35710,17'd51066,17'd46678,17'd51164,17'd50166,17'd46849,17'd31030,17'd51317,17'd32829,17'd46561,17'd51318,17'd51319,17'd51320,17'd51321,17'd51322,17'd51323,17'd51324,17'd51325,17'd49398,17'd7166,17'd5916,17'd5159,17'd26708,17'd8304,17'd7499,17'd28058,17'd6392,17'd27571,17'd30486,17'd38441,17'd4186,17'd5754,17'd5144,17'd4841,17'd5160,17'd28185,17'd6554,17'd6554,17'd28185,17'd5160,17'd5002,17'd4842,17'd28418,17'd28536,17'd28418,17'd4842,17'd5004,17'd25627,17'd30638,17'd30638,17'd30638,17'd28185,17'd6554,17'd6390,17'd6390,17'd27935,17'd30638,17'd30333,17'd30333,17'd30638,17'd36887,17'd5165,17'd51175,17'd51175,17'd5010,17'd5011,17'd4849,17'd51247,17'd51326,17'd51327,17'd51328,17'd39171,17'd51329,17'd51330,17'd2881,17'd51331,17'd41312,17'd51332,17'd22262,17'd51333,17'd40860,17'd51251,17'd51252,17'd51334,17'd3870,17'd39947,17'd10790,17'd10906,17'd11048,17'd38202,17'd37957,17'd37821,17'd2586,17'd1119,17'd228,17'd228,17'd1119,17'd2586,17'd50843,17'd50843,17'd50843,17'd50843,17'd3898,17'd1825,17'd38071,17'd1120,17'd1122,17'd234,17'd633,17'd453,17'd592,17'd612,17'd51335,17'd51336,17'd434,17'd51337
},
'{
17'd14188,17'd3252,17'd2596,17'd1414,17'd289,17'd652,17'd286,17'd286,17'd26,17'd26,17'd285,17'd467,17'd2937,17'd467,17'd7555,17'd7385,17'd286,17'd980,17'd4430,17'd4430,17'd4091,17'd4091,17'd3755,17'd3595,17'd3255,17'd3255,17'd3104,17'd3105,17'd25790,17'd14192,17'd5219,17'd4092,17'd33052,17'd31259,17'd30348,17'd29043,17'd23492,17'd6609,17'd51338,17'd13077,17'd51339,17'd12797,17'd15756,17'd18166,17'd16762,17'd17571,17'd12679,17'd24345,17'd12065,17'd13094,17'd12955,17'd13093,17'd12678,17'd12062,17'd13461,17'd13461,17'd13460,17'd13460,17'd13595,17'd12212,17'd12212,17'd12212,17'd13596,17'd13838,17'd12215,17'd13599,17'd12530,17'd11764,17'd12361,17'd12361,17'd12681,17'd18774,17'd16519,17'd15902,17'd16034,17'd17319,17'd17206,17'd10945,17'd10429,17'd9440,17'd46366,17'd6142,17'd7750,17'd5255,17'd7252,17'd5250,17'd6933,17'd7258,17'd6637,17'd46489,17'd51256,17'd49015,17'd39504,17'd6645,17'd38603,17'd6788,17'd51340,17'd40879,17'd50847,17'd50765,17'd51105,17'd51341,17'd38894,17'd38487,17'd37060,17'd34369,17'd30060,17'd28929,17'd51342,17'd27331,17'd27110,17'd27724,17'd50511,17'd24202,17'd51343,17'd51191,17'd51192,17'd51344,17'd10449,17'd51345,17'd32588,17'd10589,17'd9874,17'd9881,17'd51346,17'd51269,17'd11518,17'd29493,17'd11956,17'd11804,17'd11956,17'd51347,17'd17837,17'd29492,17'd47110,17'd12998,17'd13365,17'd13517,17'd34558,17'd48846,17'd48846,17'd13515,17'd13517,17'd13517,17'd15685,17'd50779,17'd50779,17'd50779,17'd17603,17'd17474,17'd12108,17'd24991,17'd28103,17'd35372,17'd30220,17'd34835,17'd34380,17'd51118,17'd50863,17'd50952,17'd51272,17'd50863,17'd34380,17'd34203,17'd30221,17'd30373,17'd28104,17'd24856,17'd25926,17'd24858,17'd18327,17'd24029,17'd24029,17'd11274,17'd10989,17'd10989,17'd14262,17'd10989,17'd10990,17'd10854,17'd10476,17'd11132,17'd19282,17'd19282,17'd24996,17'd11132,17'd10478,17'd10479,17'd17011,17'd9345,17'd15944,17'd17480,17'd10336,17'd10336,17'd22813,17'd9743,17'd9743,17'd9340,17'd9479,17'd9619,17'd14928,17'd29068,17'd15181,17'd14518,17'd10326,17'd10855,17'd16320,17'd15052,17'd17236,17'd17236,17'd17236,17'd11523,17'd24210,17'd14803,17'd45549,17'd51348,17'd51349,17'd51350,17'd51351,17'd51352,17'd51353,17'd50611,17'd51354,17'd50699,17'd42238,17'd51355,17'd51356,17'd51357,17'd51358,17'd51359,17'd51360,17'd51361,17'd51362,17'd51363,17'd51364,17'd51365,17'd51366,17'd51367,17'd51368,17'd51369,17'd51370,17'd51371,17'd51372,17'd51373,17'd22667,17'd51374,17'd51375,17'd51376,17'd51377,17'd51378,17'd51316,17'd32662,17'd51379,17'd51380,17'd46428,17'd22161,17'd45616,17'd50732,17'd22325,17'd32345,17'd50274,17'd51381,17'd51382,17'd51383,17'd51384,17'd46861,17'd51385,17'd31497,17'd32999,17'd46096,17'd50899,17'd51386,17'd51387,17'd51388,17'd51389,17'd48047,17'd46199,17'd48263,17'd50467,17'd50267,17'd49683,17'd49692,17'd49389,17'd49484,17'd49890,17'd51390,17'd49989,17'd51391,17'd45984,17'd40825,17'd36127,17'd32355,17'd29107,17'd32505,17'd32506,17'd30586,17'd28978,17'd25565,17'd28369,17'd29976,17'd23732,17'd29829,17'd40962,17'd32680,17'd51392,17'd25708,17'd27027,17'd32832,17'd29247,17'd31504,17'd29978,17'd30280,17'd33489,17'd49887,17'd31505,17'd31036,17'd30738,17'd30131,17'd33323,17'd33489,17'd30131,17'd29978,17'd30740,17'd51393,17'd36401,17'd40519,17'd44936,17'd43544,17'd48534,17'd49390,17'd50271,17'd50661,17'd51236,17'd51163,17'd50272,17'd50072,17'd50164,17'd49582,17'd48264,17'd48781,17'd46760,17'd47334,17'd25707,17'd28482,17'd28594,17'd29101,17'd24897,17'd29378,17'd29374,17'd39131,17'd35296,17'd35429,17'd35017,17'd46570,17'd46570,17'd46669,17'd33480,17'd49487,17'd43982,17'd45265,17'd21695,17'd50984,17'd50984,17'd22511,17'd42440,17'd51238,17'd51394,17'd42152,17'd49990,17'd46106,17'd44701,17'd21848,17'd30880,17'd45990,17'd51395,17'd51396,17'd51397,17'd51398,17'd51399,17'd51400,17'd51401,17'd51402,17'd27197,17'd6845,17'd5916,17'd50175,17'd26708,17'd8304,17'd9091,17'd28058,17'd6392,17'd33692,17'd38317,17'd40081,17'd43584,17'd5477,17'd5144,17'd4686,17'd5335,17'd28185,17'd6390,17'd6554,17'd28185,17'd30638,17'd5004,17'd4842,17'd28418,17'd28536,17'd28418,17'd4842,17'd5004,17'd5160,17'd30638,17'd30638,17'd28185,17'd28185,17'd6554,17'd6390,17'd6219,17'd6390,17'd28185,17'd30638,17'd30638,17'd28185,17'd36887,17'd5165,17'd5164,17'd5164,17'd5011,17'd5012,17'd4849,17'd51247,17'd51326,17'd51403,17'd51404,17'd51405,17'd51329,17'd51406,17'd2881,17'd51407,17'd51408,17'd51409,17'd22262,17'd51410,17'd40860,17'd51411,17'd51412,17'd51334,17'd3870,17'd39947,17'd10790,17'd40716,17'd51413,17'd38202,17'd37957,17'd37821,17'd2586,17'd1119,17'd228,17'd228,17'd1119,17'd2586,17'd50843,17'd50843,17'd4712,17'd4712,17'd3898,17'd795,17'd628,17'd628,17'd1122,17'd234,17'd245,17'd51414,17'd1547,17'd441,17'd1238,17'd21467,17'd766,17'd18867
},
'{
17'd14188,17'd10535,17'd2257,17'd1416,17'd653,17'd652,17'd286,17'd285,17'd26,17'd285,17'd467,17'd2937,17'd2937,17'd467,17'd21631,17'd7385,17'd7061,17'd27444,17'd4430,17'd4430,17'd4091,17'd4091,17'd3755,17'd3595,17'd3255,17'd3255,17'd3435,17'd4250,17'd5805,17'd14192,17'd5219,17'd51415,17'd32088,17'd25792,17'd4097,17'd29043,17'd4266,17'd51416,17'd51338,17'd13077,17'd51339,17'd12797,17'd15756,17'd51417,17'd16762,17'd51418,17'd12679,17'd24345,17'd12065,17'd12814,17'd12955,17'd12679,17'd12357,17'd12062,17'd12355,17'd12355,17'd13596,17'd13596,17'd13595,17'd12212,17'd13837,17'd13837,17'd13596,17'd13838,17'd12215,17'd13093,17'd12530,17'd11764,17'd12530,17'd12361,17'd16658,17'd19382,17'd21185,17'd17320,17'd17445,17'd17319,17'd17206,17'd10945,17'd10429,17'd8537,17'd9158,17'd9701,17'd8537,17'd5255,17'd7252,17'd5250,17'd4923,17'd7258,17'd6637,17'd46489,17'd51256,17'd49203,17'd51419,17'd6645,17'd38603,17'd6788,17'd51340,17'd6789,17'd50764,17'd51420,17'd51105,17'd51421,17'd40429,17'd38355,17'd51260,17'd51422,17'd50198,17'd51423,17'd51342,17'd51424,17'd51425,17'd27332,17'd50403,17'd50404,17'd51426,17'd17222,17'd51427,17'd51428,17'd15798,17'd51429,17'd31938,17'd10454,17'd51430,17'd9875,17'd10019,17'd38112,17'd38111,17'd37988,17'd28680,17'd17597,17'd17597,17'd51431,17'd51347,17'd40746,17'd47199,17'd15809,17'd13365,17'd12995,17'd15570,17'd48846,17'd48846,17'd34558,17'd13517,17'd13517,17'd15433,17'd50862,17'd17603,17'd17967,17'd17967,17'd17967,17'd17348,17'd12255,17'd28107,17'd30222,17'd28686,17'd31765,17'd31288,17'd35644,17'd50863,17'd50863,17'd50952,17'd51272,17'd51432,17'd33243,17'd34381,17'd29785,17'd28571,17'd28816,17'd24705,17'd24993,17'd23169,17'd22817,17'd24029,17'd11274,17'd10989,17'd18560,17'd14262,17'd14262,17'd14931,17'd10990,17'd10476,17'd11132,17'd11132,17'd11132,17'd19282,17'd19282,17'd11132,17'd11527,17'd14928,17'd9479,17'd15807,17'd14674,17'd15807,17'd15807,17'd10173,17'd9346,17'd23679,17'd9340,17'd9480,17'd9741,17'd11277,17'd25675,17'd15943,17'd25812,17'd10479,17'd17124,17'd10166,17'd11133,17'd10606,17'd11527,17'd14134,17'd16687,17'd17236,17'd13001,17'd16908,17'd50953,17'd49637,17'd49746,17'd51433,17'd51434,17'd51435,17'd51436,17'd51437,17'd51438,17'd51439,17'd51440,17'd51441,17'd51442,17'd51443,17'd51444,17'd51445,17'd51446,17'd51447,17'd51448,17'd51449,17'd51450,17'd51451,17'd51452,17'd51453,17'd51454,17'd51455,17'd51456,17'd51457,17'd51458,17'd51459,17'd51460,17'd51461,17'd51462,17'd51463,17'd51464,17'd51065,17'd42002,17'd41585,17'd51465,17'd51466,17'd33650,17'd51229,17'd22504,17'd31831,17'd35155,17'd51467,17'd51468,17'd51469,17'd51470,17'd51471,17'd51067,17'd51472,17'd32013,17'd22327,17'd51473,17'd51233,17'd51474,17'd51310,17'd51475,17'd49374,17'd51476,17'd49091,17'd49184,17'd49478,17'd49575,17'd49794,17'd49583,17'd50822,17'd49692,17'd50574,17'd51390,17'd50654,17'd48259,17'd44476,17'd36690,17'd32831,17'd32018,17'd29536,17'd28371,17'd47440,17'd25702,17'd31351,17'd25435,17'd29103,17'd28851,17'd23565,17'd37386,17'd51477,17'd38669,17'd33157,17'd27515,17'd28979,17'd28258,17'd28257,17'd31196,17'd29978,17'd30736,17'd31506,17'd49887,17'd31506,17'd31036,17'd30130,17'd30131,17'd34460,17'd32021,17'd31838,17'd29981,17'd51478,17'd50824,17'd36537,17'd50473,17'd44932,17'd39581,17'd48360,17'd49693,17'd42874,17'd43012,17'd51236,17'd51236,17'd51163,17'd50072,17'd49890,17'd49682,17'd48535,17'd49889,17'd46433,17'd43838,17'd27515,17'd26062,17'd27765,17'd29103,17'd28718,17'd29377,17'd23217,17'd22859,17'd37659,17'd35296,17'd35455,17'd44233,17'd46570,17'd45492,17'd32013,17'd31659,17'd49892,17'd43158,17'd33648,17'd50984,17'd34457,17'd35015,17'd51479,17'd46775,17'd51394,17'd51226,17'd51480,17'd45990,17'd44701,17'd50987,17'd21850,17'd45373,17'd51481,17'd46568,17'd51482,17'd51483,17'd51484,17'd51485,17'd51486,17'd51487,17'd29022,17'd5915,17'd5332,17'd50175,17'd6390,17'd7668,17'd9091,17'd28058,17'd26828,17'd4841,17'd51488,17'd33208,17'd5604,17'd33041,17'd38442,17'd4686,17'd28185,17'd6554,17'd6390,17'd6554,17'd28185,17'd25627,17'd5002,17'd4842,17'd28418,17'd28536,17'd28418,17'd5005,17'd25627,17'd5160,17'd30638,17'd30638,17'd28185,17'd28185,17'd6554,17'd6390,17'd6219,17'd6390,17'd28185,17'd30638,17'd30638,17'd28185,17'd36887,17'd5165,17'd5164,17'd5165,17'd5012,17'd5012,17'd5007,17'd51247,17'd51326,17'd51489,17'd51490,17'd51491,17'd51329,17'd48468,17'd51492,17'd42042,17'd51493,17'd21783,17'd51494,17'd2730,17'd51495,17'd50496,17'd41478,17'd3562,17'd4056,17'd39947,17'd10790,17'd10906,17'd5355,17'd38202,17'd37957,17'd37821,17'd1119,17'd228,17'd228,17'd228,17'd4712,17'd50843,17'd50843,17'd50843,17'd4712,17'd4400,17'd1824,17'd795,17'd628,17'd629,17'd798,17'd451,17'd245,17'd1547,17'd454,17'd432,17'd39034,17'd21324,17'd51496,17'd51497
},
'{
17'd14188,17'd3252,17'd2597,17'd1414,17'd289,17'd28,17'd286,17'd285,17'd285,17'd285,17'd467,17'd467,17'd2937,17'd467,17'd21631,17'd7385,17'd7061,17'd27444,17'd4430,17'd4430,17'd4091,17'd4091,17'd3755,17'd3595,17'd3255,17'd3255,17'd3435,17'd3104,17'd25790,17'd14192,17'd5219,17'd51415,17'd32088,17'd25792,17'd4097,17'd29043,17'd4266,17'd51416,17'd51338,17'd51498,17'd51339,17'd12797,17'd15756,17'd51417,17'd51499,17'd51418,17'd12527,17'd24345,17'd12065,17'd12814,17'd12955,17'd12679,17'd12357,17'd12062,17'd12355,17'd12355,17'd13596,17'd13596,17'd13595,17'd13595,17'd13837,17'd13837,17'd13596,17'd12355,17'd10937,17'd13093,17'd12530,17'd11764,17'd12530,17'd12362,17'd16765,17'd19006,17'd21185,17'd17320,17'd17445,17'd17319,17'd17206,17'd20023,17'd10429,17'd9440,17'd9702,17'd6142,17'd7750,17'd4767,17'd7751,17'd4924,17'd4923,17'd7584,17'd6638,17'd50930,17'd46999,17'd49203,17'd51419,17'd39057,17'd38350,17'd38482,17'd40586,17'd6789,17'd50764,17'd51420,17'd51105,17'd51105,17'd40429,17'd51500,17'd51259,17'd51501,17'd50298,17'd51502,17'd30662,17'd27723,17'd51424,17'd51503,17'd51504,17'd50511,17'd51505,17'd20599,17'd51506,17'd51507,17'd51508,17'd51509,17'd28452,17'd32757,17'd51510,17'd9876,17'd10019,17'd38112,17'd36079,17'd36357,17'd51431,17'd28680,17'd17597,17'd28680,17'd51347,17'd40746,17'd51511,17'd15809,17'd13365,17'd13517,17'd13515,17'd34558,17'd48846,17'd34558,17'd13517,17'd13517,17'd15433,17'd15433,17'd17603,17'd17967,17'd17843,17'd17843,17'd17603,17'd19407,17'd23511,17'd28230,17'd31286,17'd39211,17'd33568,17'd34037,17'd35644,17'd50863,17'd50951,17'd51512,17'd51513,17'd35100,17'd34203,17'd34381,17'd31587,17'd28344,17'd27483,17'd26495,17'd24858,17'd24994,17'd22817,17'd13516,17'd18560,17'd18560,17'd13762,17'd11964,17'd14673,17'd14931,17'd13886,17'd10476,17'd10476,17'd10476,17'd10476,17'd19282,17'd19282,17'd14518,17'd11528,17'd9741,17'd9480,17'd15187,17'd15569,17'd15569,17'd15569,17'd15187,17'd9480,17'd9480,17'd9742,17'd9742,17'd14928,17'd11277,17'd10479,17'd15943,17'd15943,17'd11134,17'd10327,17'd21503,17'd9473,17'd12116,17'd27490,17'd19779,17'd10331,17'd26037,17'd51514,17'd45934,17'd50953,17'd51515,17'd51516,17'd51433,17'd51517,17'd51518,17'd51519,17'd51520,17'd51521,17'd51522,17'd51523,17'd51524,17'd51525,17'd51526,17'd45217,17'd51527,17'd51528,17'd51529,17'd51530,17'd51531,17'd51532,17'd51533,17'd51534,17'd21522,17'd51535,17'd51536,17'd51537,17'd51538,17'd51539,17'd51540,17'd51301,17'd51541,17'd51542,17'd21532,17'd51164,17'd51543,17'd51544,17'd22002,17'd49096,17'd36846,17'd22505,17'd36691,17'd51464,17'd51545,17'd51546,17'd51547,17'd51548,17'd51549,17'd51550,17'd51551,17'd34457,17'd30728,17'd51552,17'd51553,17'd51554,17'd50263,17'd51555,17'd51556,17'd47724,17'd51557,17'd43419,17'd50267,17'd49787,17'd49787,17'd49582,17'd49582,17'd49583,17'd49890,17'd50273,17'd50568,17'd49084,17'd47345,17'd42741,17'd31503,17'd32505,17'd34285,17'd28857,17'd28371,17'd27368,17'd25948,17'd35012,17'd28369,17'd25030,17'd24249,17'd29376,17'd51558,17'd51559,17'd37512,17'd28366,17'd27371,17'd29246,17'd33485,17'd28372,17'd28857,17'd30130,17'd31036,17'd31506,17'd49887,17'd31506,17'd30736,17'd30130,17'd30131,17'd34460,17'd32021,17'd31838,17'd31037,17'd51560,17'd50824,17'd36537,17'd46950,17'd44587,17'd42596,17'd49091,17'd49988,17'd50907,17'd43146,17'd51236,17'd51163,17'd50272,17'd50574,17'd49794,17'd49289,17'd46199,17'd49287,17'd51561,17'd45749,17'd27514,17'd26062,17'd27765,17'd25179,17'd34884,17'd29687,17'd41273,17'd22858,17'd31657,17'd31343,17'd40833,17'd36414,17'd43986,17'd48913,17'd31344,17'd33648,17'd50576,17'd50576,17'd23041,17'd31831,17'd21693,17'd35294,17'd51562,17'd51563,17'd46775,17'd42439,17'd50073,17'd34455,17'd47358,17'd22013,17'd21843,17'd51564,17'd51565,17'd51566,17'd51567,17'd51568,17'd51569,17'd41883,17'd51570,17'd50669,17'd30331,17'd51571,17'd5761,17'd5159,17'd6219,17'd7668,17'd9091,17'd6391,17'd5336,17'd4996,17'd51572,17'd51573,17'd51574,17'd43584,17'd38442,17'd4686,17'd28185,17'd6390,17'd6390,17'd6554,17'd28185,17'd30333,17'd5004,17'd4842,17'd28418,17'd28536,17'd28418,17'd5005,17'd25627,17'd5160,17'd30638,17'd30638,17'd28185,17'd27935,17'd6554,17'd6390,17'd6219,17'd6390,17'd28185,17'd30638,17'd28185,17'd27935,17'd36887,17'd5165,17'd5164,17'd37030,17'd5012,17'd5012,17'd5007,17'd51247,17'd51326,17'd49599,17'd51575,17'd47564,17'd37812,17'd51576,17'd51014,17'd38713,17'd51577,17'd51578,17'd2899,17'd51579,17'd51495,17'd51580,17'd51581,17'd3702,17'd5493,17'd39947,17'd10790,17'd40716,17'd51253,17'd38202,17'd37957,17'd5939,17'd1119,17'd228,17'd1260,17'd228,17'd4712,17'd50843,17'd4712,17'd4712,17'd4400,17'd4400,17'd1825,17'd1264,17'd628,17'd629,17'd451,17'd242,17'd1540,17'd247,17'd248,17'd31099,17'd21944,17'd51582,17'd20265,17'd51497
},
'{
17'd14188,17'd3252,17'd2597,17'd1414,17'd289,17'd27,17'd285,17'd285,17'd285,17'd467,17'd467,17'd467,17'd467,17'd467,17'd21631,17'd50387,17'd7385,17'd27444,17'd4430,17'd4430,17'd4091,17'd4091,17'd3755,17'd3595,17'd3255,17'd3255,17'd3435,17'd4250,17'd5805,17'd5805,17'd4742,17'd4744,17'd32088,17'd25792,17'd4097,17'd29043,17'd6448,17'd12042,17'd23665,17'd51498,17'd51339,17'd12665,17'd20581,17'd19749,17'd51499,17'd51418,17'd12527,17'd24345,17'd11626,17'd12065,17'd12528,17'd12679,17'd12357,17'd12062,17'd13461,17'd13461,17'd13596,17'd13596,17'd13596,17'd13596,17'd13837,17'd13837,17'd13596,17'd13838,17'd12215,17'd12813,17'd12530,17'd11913,17'd12218,17'd13094,17'd12362,17'd18884,17'd16986,17'd17207,17'd17207,17'd17319,17'd17206,17'd20023,17'd10429,17'd9702,17'd9158,17'd9573,17'd8537,17'd4927,17'd51583,17'd4924,17'd4923,17'd7584,17'd6638,17'd51584,17'd51585,17'd51586,17'd49015,17'd39057,17'd38890,17'd40275,17'd51185,17'd6949,17'd51587,17'd50764,17'd50505,17'd50765,17'd51588,17'd40277,17'd51589,17'd51590,17'd8083,17'd51591,17'd51592,17'd29766,17'd27466,17'd27467,17'd27469,17'd25807,17'd51593,17'd51594,17'd17222,17'd51595,17'd26360,17'd51596,17'd28093,17'd51597,17'd51598,17'd51599,17'd28682,17'd10731,17'd35655,17'd29938,17'd30216,17'd28567,17'd51600,17'd28567,17'd51431,17'd51347,17'd21819,17'd18077,17'd13365,17'd12856,17'd12417,17'd13515,17'd34558,17'd13515,17'd13517,17'd12995,17'd15570,17'd15433,17'd17603,17'd12581,17'd18328,17'd17843,17'd18197,17'd20314,17'd23512,17'd25672,17'd51601,17'd36777,17'd31773,17'd33875,17'd35644,17'd50863,17'd50951,17'd51512,17'd51602,17'd51603,17'd33243,17'd31289,17'd30972,17'd30370,17'd32435,17'd34962,17'd51604,17'd23513,17'd21985,17'd13516,17'd18560,17'd18560,17'd12262,17'd13762,17'd14673,17'd14931,17'd13886,17'd14134,17'd14134,17'd12721,17'd11399,17'd11669,17'd10475,17'd14518,17'd15943,17'd14928,17'd9479,17'd9620,17'd9478,17'd24037,17'd23857,17'd23857,17'd9619,17'd17011,17'd9885,17'd10992,17'd11671,17'd9884,17'd11671,17'd17599,17'd26037,17'd10478,17'd10329,17'd18916,17'd48577,17'd12117,17'd15807,17'd37336,17'd17473,17'd33237,17'd51605,17'd17715,17'd14803,17'd15940,17'd15681,17'd49324,17'd51519,17'd51606,17'd51519,17'd51607,17'd51608,17'd51609,17'd51610,17'd51611,17'd51612,17'd51613,17'd51614,17'd51615,17'd51616,17'd51617,17'd51618,17'd20928,17'd51619,17'd51620,17'd51621,17'd51622,17'd51623,17'd51624,17'd51625,17'd51626,17'd51627,17'd51628,17'd51629,17'd51630,17'd51468,17'd51631,17'd51632,17'd46678,17'd51633,17'd51634,17'd51635,17'd51228,17'd49487,17'd22686,17'd51636,17'd51637,17'd51638,17'd51639,17'd51640,17'd21227,17'd51641,17'd51642,17'd31344,17'd45379,17'd51232,17'd50646,17'd51643,17'd51644,17'd51645,17'd51389,17'd51646,17'd48153,17'd49682,17'd49788,17'd51647,17'd49787,17'd49682,17'd51648,17'd49988,17'd50365,17'd51236,17'd50568,17'd51649,17'd49085,17'd40520,17'd28373,17'd32507,17'd34285,17'd30884,17'd28372,17'd25558,17'd25703,17'd28253,17'd25178,17'd28008,17'd30275,17'd35865,17'd51558,17'd35022,17'd51650,17'd25707,17'd34767,17'd29977,17'd32505,17'd29537,17'd29536,17'd29978,17'd31036,17'd31506,17'd31506,17'd30736,17'd30736,17'd30130,17'd29979,17'd34460,17'd32021,17'd31838,17'd30434,17'd51560,17'd50824,17'd38665,17'd51651,17'd46947,17'd48358,17'd43419,17'd49890,17'd50739,17'd43144,17'd51652,17'd51236,17'd50661,17'd49985,17'd49691,17'd48622,17'd49581,17'd47638,17'd51653,17'd33642,17'd26530,17'd28481,17'd28369,17'd24898,17'd29102,17'd48257,17'd32830,17'd35711,17'd37659,17'd22506,17'd46115,17'd36414,17'd23570,17'd40523,17'd31659,17'd48457,17'd43158,17'd49892,17'd31346,17'd31660,17'd22510,17'd42603,17'd46775,17'd51654,17'd51655,17'd41112,17'd33798,17'd34455,17'd50987,17'd51656,17'd51657,17'd22512,17'd51658,17'd34641,17'd51659,17'd51660,17'd51661,17'd23772,17'd26212,17'd11013,17'd6844,17'd6552,17'd5158,17'd5159,17'd6219,17'd6391,17'd6220,17'd6221,17'd5329,17'd51662,17'd40396,17'd33207,17'd33040,17'd43584,17'd5145,17'd4845,17'd28185,17'd32073,17'd6390,17'd6554,17'd28185,17'd25627,17'd5002,17'd5005,17'd28418,17'd28536,17'd28418,17'd5005,17'd25627,17'd5160,17'd30638,17'd28185,17'd28185,17'd27935,17'd6390,17'd6219,17'd6219,17'd6390,17'd28185,17'd30638,17'd28185,17'd27935,17'd36887,17'd5165,17'd5164,17'd37030,17'd5169,17'd5012,17'd51663,17'd51326,17'd51177,17'd51664,17'd51665,17'd47374,17'd3540,17'd51666,17'd51667,17'd51668,17'd51669,17'd51578,17'd2899,17'd51579,17'd51670,17'd9100,17'd51581,17'd3562,17'd4056,17'd39947,17'd10790,17'd10906,17'd11048,17'd38202,17'd5938,17'd51671,17'd228,17'd228,17'd446,17'd625,17'd4712,17'd4712,17'd4712,17'd4400,17'd4229,17'd1824,17'd1402,17'd447,17'd629,17'd629,17'd451,17'd243,17'd792,17'd38862,17'd51672,17'd455,17'd51336,17'd36907,17'd51673,17'd51674
},
'{
17'd14188,17'd3252,17'd2597,17'd1414,17'd653,17'd27,17'd286,17'd286,17'd1833,17'd467,17'd467,17'd467,17'd467,17'd1691,17'd21631,17'd7385,17'd7061,17'd27444,17'd4430,17'd4430,17'd4091,17'd4091,17'd3755,17'd3595,17'd3255,17'd3255,17'd3435,17'd3104,17'd4739,17'd5805,17'd4742,17'd51415,17'd32088,17'd25792,17'd4097,17'd29043,17'd12041,17'd12042,17'd6916,17'd51498,17'd51339,17'd12665,17'd13082,17'd14203,17'd51499,17'd51418,17'd12527,17'd24345,17'd11626,17'd11626,17'd12528,17'd12679,17'd12357,17'd12062,17'd13461,17'd13461,17'd13596,17'd13596,17'd13596,17'd13596,17'd13837,17'd13837,17'd13596,17'd13461,17'd51675,17'd12527,17'd12218,17'd12361,17'd12218,17'd13094,17'd12362,17'd12531,17'd17205,17'd17319,17'd17207,17'd17319,17'd17206,17'd20023,17'd16410,17'd13471,17'd9702,17'd46366,17'd8537,17'd4927,17'd51583,17'd4126,17'd3950,17'd7584,17'd6476,17'd51584,17'd51585,17'd51676,17'd50392,17'd39057,17'd6643,17'd38890,17'd38603,17'd6949,17'd50933,17'd51677,17'd51678,17'd50765,17'd6790,17'd51679,17'd51680,17'd51681,17'd50682,17'd51682,17'd7929,17'd30662,17'd51683,17'd27467,17'd9595,17'd50853,17'd51684,17'd51685,17'd18072,17'd17002,17'd16787,17'd51686,17'd51687,17'd51688,17'd51689,17'd51690,17'd9878,17'd51691,17'd35807,17'd38111,17'd16906,17'd28567,17'd51600,17'd28567,17'd51431,17'd51347,17'd21819,17'd21502,17'd13365,17'd12856,17'd12417,17'd13517,17'd34558,17'd13515,17'd13517,17'd12995,17'd13517,17'd15685,17'd17603,17'd12581,17'd17843,17'd17843,17'd12582,17'd19409,17'd22819,17'd24859,17'd30525,17'd40439,17'd39211,17'd33568,17'd34380,17'd50863,17'd35239,17'd51692,17'd51693,17'd51694,17'd34705,17'd34037,17'd34381,17'd31587,17'd34696,17'd51695,17'd27122,17'd33084,17'd18681,17'd13516,17'd10989,17'd18560,17'd15810,17'd14262,17'd14262,17'd11274,17'd11524,17'd11524,17'd11524,17'd11524,17'd21206,17'd21206,17'd10739,17'd16320,17'd10477,17'd11528,17'd9741,17'd18442,17'd25281,17'd18080,17'd33083,17'd23857,17'd15048,17'd9740,17'd10856,17'd16796,17'd16796,17'd19278,17'd11276,17'd19642,17'd26037,17'd21205,17'd11132,17'd17719,17'd16554,17'd24039,17'd10336,17'd51696,17'd37850,17'd32123,17'd25146,17'd26630,17'd14134,17'd12721,17'd51697,17'd28578,17'd47407,17'd51698,17'd51699,17'd28707,17'd51700,17'd51701,17'd51702,17'd51703,17'd51704,17'd51705,17'd51706,17'd51707,17'd51708,17'd51709,17'd51710,17'd51711,17'd51712,17'd51713,17'd51714,17'd20767,17'd51715,17'd22148,17'd51716,17'd21222,17'd51717,17'd51718,17'd51719,17'd51720,17'd51721,17'd21541,17'd51722,17'd51394,17'd51723,17'd51724,17'd51725,17'd33648,17'd33646,17'd51726,17'd51727,17'd51728,17'd51729,17'd51730,17'd51731,17'd51732,17'd51147,17'd51733,17'd31658,17'd51734,17'd51735,17'd51736,17'd51737,17'd51738,17'd51739,17'd47534,17'd51740,17'd43281,17'd49794,17'd50568,17'd51390,17'd49683,17'd51648,17'd49691,17'd49890,17'd50268,17'd51741,17'd49883,17'd51742,17'd49177,17'd33790,17'd32505,17'd33321,17'd34285,17'd30884,17'd28257,17'd26279,17'd26168,17'd44229,17'd25031,17'd29532,17'd23385,17'd23566,17'd51743,17'd39292,17'd39449,17'd27640,17'd47145,17'd33319,17'd32505,17'd29536,17'd29690,17'd29979,17'd31036,17'd31506,17'd31506,17'd31506,17'd30736,17'd29978,17'd29979,17'd34460,17'd32021,17'd33167,17'd29981,17'd51478,17'd50824,17'd41998,17'd48705,17'd43543,17'd41579,17'd48995,17'd49986,17'd50661,17'd51744,17'd51745,17'd51236,17'd50661,17'd49985,17'd49682,17'd48535,17'd48621,17'd47339,17'd51746,17'd38538,17'd28482,17'd30606,17'd27882,17'd24417,17'd29972,17'd37386,17'd34458,17'd51747,17'd35296,17'd22331,17'd36414,17'd34452,17'd32513,17'd33944,17'd33796,17'd22510,17'd43158,17'd31659,17'd31497,17'd31659,17'd35295,17'd41584,17'd51067,17'd51748,17'd51655,17'd41584,17'd33796,17'd48912,17'd51749,17'd51656,17'd22494,17'd48269,17'd51750,17'd36154,17'd51751,17'd51752,17'd51753,17'd22050,17'd51754,17'd7165,17'd28532,17'd6552,17'd5612,17'd26218,17'd6219,17'd6391,17'd6391,17'd5919,17'd4686,17'd51755,17'd51756,17'd43585,17'd5910,17'd33041,17'd6067,17'd5002,17'd6554,17'd32073,17'd6219,17'd6554,17'd28185,17'd25627,17'd5002,17'd5005,17'd28418,17'd28536,17'd4842,17'd5005,17'd25627,17'd5160,17'd30638,17'd28185,17'd28185,17'd27935,17'd6390,17'd6219,17'd6219,17'd6390,17'd31717,17'd30638,17'd28185,17'd27935,17'd36887,17'd5164,17'd5164,17'd36887,17'd5169,17'd5012,17'd51663,17'd51326,17'd51010,17'd38706,17'd50750,17'd46987,17'd37296,17'd51757,17'd45184,17'd51758,17'd51759,17'd51578,17'd2899,17'd51579,17'd40999,17'd51183,17'd51760,17'd3562,17'd48811,17'd39947,17'd10790,17'd10906,17'd11048,17'd38202,17'd5938,17'd51761,17'd228,17'd1260,17'd446,17'd446,17'd4400,17'd4712,17'd4712,17'd4400,17'd1824,17'd1824,17'd1402,17'd1264,17'd628,17'd629,17'd451,17'd784,17'd955,17'd248,17'd51762,17'd51763,17'd21467,17'd18759,17'd51764,17'd51765
},
'{
17'd3251,17'd3252,17'd2257,17'd17,17'd653,17'd980,17'd286,17'd1833,17'd286,17'd1833,17'd467,17'd1691,17'd21631,17'd21631,17'd51766,17'd51767,17'd7385,17'd7060,17'd4430,17'd4430,17'd4091,17'd4091,17'd3755,17'd3595,17'd3754,17'd3754,17'd3435,17'd5210,17'd5055,17'd5806,17'd5805,17'd4581,17'd4897,17'd25792,17'd29176,17'd28194,17'd27954,17'd25793,17'd23495,17'd12513,17'd20141,17'd10555,17'd51768,17'd19003,17'd16982,17'd51769,17'd12678,17'd12527,17'd12813,17'd13093,17'd12679,17'd12679,17'd12357,17'd12062,17'd12355,17'd13461,17'd15761,17'd13596,17'd13595,17'd12212,17'd12212,17'd12212,17'd13596,17'd13596,17'd12355,17'd12357,17'd14764,17'd14622,17'd13211,17'd14621,17'd13094,17'd11764,17'd17204,17'd18656,17'd18657,17'd17319,17'd17318,17'd17318,17'd16410,17'd15765,17'd15765,17'd13602,17'd7418,17'd14218,17'd51770,17'd3951,17'd3950,17'd6629,17'd6638,17'd6634,17'd51771,17'd51676,17'd51101,17'd51772,17'd51773,17'd38604,17'd51774,17'd51775,17'd51776,17'd50933,17'd51777,17'd51777,17'd51420,17'd51679,17'd6951,17'd51778,17'd51590,17'd51779,17'd51682,17'd51780,17'd51781,17'd50401,17'd51782,17'd27469,17'd51109,17'd51685,17'd17113,17'd21198,17'd18553,17'd26252,17'd15166,17'd51783,17'd51784,17'd51785,17'd10015,17'd10018,17'd10321,17'd36788,17'd29634,17'd16906,17'd51600,17'd51600,17'd51786,17'd51787,17'd28221,17'd51788,17'd51789,17'd13881,17'd12856,17'd12856,17'd12417,17'd12417,17'd12995,17'd12995,17'd13518,17'd21506,17'd15685,17'd14670,17'd17843,17'd17843,17'd18806,17'd19410,17'd21362,17'd23512,17'd24856,17'd28103,17'd31286,17'd31439,17'd31441,17'd31943,17'd35644,17'd35239,17'd51512,17'd51692,17'd51512,17'd35239,17'd33720,17'd31941,17'd30072,17'd29066,17'd27346,17'd24705,17'd20608,17'd18444,17'd11965,17'd10737,17'd10737,17'd14262,17'd14262,17'd14262,17'd14673,17'd11274,17'd11274,17'd10990,17'd12720,17'd14132,17'd16320,17'd10604,17'd19532,17'd14518,17'd10478,17'd23340,17'd8720,17'd48407,17'd24366,17'd15569,17'd51790,17'd40134,17'd10022,17'd10741,17'd19532,17'd19280,17'd12863,17'd12863,17'd10606,17'd14518,17'd10739,17'd10476,17'd25675,17'd16065,17'd10174,17'd10336,17'd17347,17'd33238,17'd15807,17'd19279,17'd26759,17'd25812,17'd25812,17'd26759,17'd16065,17'd17347,17'd34039,17'd50864,17'd51791,17'd51792,17'd13371,17'd51793,17'd51794,17'd51795,17'd51796,17'd51797,17'd51798,17'd51799,17'd51800,17'd51801,17'd51802,17'd51803,17'd20627,17'd20916,17'd51804,17'd51805,17'd51806,17'd51807,17'd51808,17'd51809,17'd51810,17'd51811,17'd51812,17'd51813,17'd51814,17'd51815,17'd51816,17'd22014,17'd22318,17'd51164,17'd51817,17'd51818,17'd51819,17'd51820,17'd20626,17'd51821,17'd51822,17'd51823,17'd51824,17'd51464,17'd51825,17'd51826,17'd51827,17'd51828,17'd50266,17'd50821,17'd51311,17'd51829,17'd48153,17'd49484,17'd49986,17'd50268,17'd49986,17'd49988,17'd49691,17'd49788,17'd50476,17'd51830,17'd51831,17'd49281,17'd43421,17'd45873,17'd47336,17'd28257,17'd29380,17'd29537,17'd28487,17'd26276,17'd27258,17'd32658,17'd33483,17'd24415,17'd29972,17'd23564,17'd29102,17'd34283,17'd44229,17'd25833,17'd35023,17'd28980,17'd33485,17'd38026,17'd28857,17'd29690,17'd30736,17'd31505,17'd31506,17'd31506,17'd31506,17'd30131,17'd49790,17'd30131,17'd30280,17'd30280,17'd30280,17'd29690,17'd30738,17'd51832,17'd51081,17'd51833,17'd45879,17'd48700,17'd49484,17'd50072,17'd50661,17'd51236,17'd51834,17'd43144,17'd50739,17'd49985,17'd41723,17'd44098,17'd43690,17'd48611,17'd44699,17'd25565,17'd28602,17'd27638,17'd25438,17'd28852,17'd29686,17'd22679,17'd35296,17'd35711,17'd45037,17'd22501,17'd23567,17'd29829,17'd22330,17'd22162,17'd22336,17'd51379,17'd51465,17'd36544,17'd31346,17'd33796,17'd33946,17'd51164,17'd51748,17'd51654,17'd51394,17'd21701,17'd21842,17'd21849,17'd33162,17'd32662,17'd22511,17'd51835,17'd51836,17'd51837,17'd51838,17'd51839,17'd51840,17'd19957,17'd25220,17'd6211,17'd5913,17'd6384,17'd5611,17'd6218,17'd8304,17'd8304,17'd6391,17'd5335,17'd4996,17'd40079,17'd43585,17'd51841,17'd51574,17'd4990,17'd5327,17'd25627,17'd32073,17'd32073,17'd6554,17'd31717,17'd30638,17'd25627,17'd5002,17'd5005,17'd4842,17'd28418,17'd4842,17'd5005,17'd25627,17'd5335,17'd28185,17'd30638,17'd28185,17'd27935,17'd6390,17'd6220,17'd7499,17'd32073,17'd51842,17'd50282,17'd36887,17'd5166,17'd5166,17'd5009,17'd37030,17'd36887,17'd5338,17'd5012,17'd51247,17'd51843,17'd51844,17'd51845,17'd51846,17'd51847,17'd51576,17'd24809,17'd51848,17'd51849,17'd51850,17'd51851,17'd51852,17'd51853,17'd51854,17'd51252,17'd51855,17'd51856,17'd51857,17'd43462,17'd10790,17'd18383,17'd5026,17'd38201,17'd5937,17'd4400,17'd4229,17'd4400,17'd4400,17'd4400,17'd3898,17'd5195,17'd5195,17'd3898,17'd2391,17'd795,17'd1264,17'd232,17'd447,17'd448,17'd1379,17'd24496,17'd31099,17'd21325,17'd51020,17'd433,17'd18515,17'd19492,17'd51858,17'd51859
},
'{
17'd3251,17'd3252,17'd2257,17'd17,17'd653,17'd980,17'd287,17'd2424,17'd287,17'd1833,17'd467,17'd1691,17'd51860,17'd51860,17'd51766,17'd7386,17'd7061,17'd7060,17'd4430,17'd4430,17'd4091,17'd4091,17'd3755,17'd3595,17'd3754,17'd3754,17'd3435,17'd3435,17'd5658,17'd5806,17'd5805,17'd4432,17'd51861,17'd25792,17'd51862,17'd51863,17'd27954,17'd6608,17'd51864,17'd51865,17'd20141,17'd10555,17'd12800,17'd16875,17'd18529,17'd51769,17'd12678,17'd12527,17'd12813,17'd13093,17'd12679,17'd12679,17'd12357,17'd12062,17'd13461,17'd13461,17'd13596,17'd13596,17'd12212,17'd12212,17'd12212,17'd12212,17'd13596,17'd13460,17'd12526,17'd14763,17'd51866,17'd20147,17'd19005,17'd13211,17'd12065,17'd11478,17'd17204,17'd18656,17'd18657,17'd16519,17'd16289,17'd17318,17'd16410,17'd15765,17'd15765,17'd13722,17'd8537,17'd14218,17'd51770,17'd3785,17'd3950,17'd3949,17'd7584,17'd6638,17'd6777,17'd51585,17'd51867,17'd51868,17'd51773,17'd37971,17'd38093,17'd51869,17'd51870,17'd50933,17'd51871,17'd51777,17'd51420,17'd51679,17'd51680,17'd38487,17'd51681,17'd35922,17'd51872,17'd7929,17'd29909,17'd9025,17'd51782,17'd9595,17'd51873,17'd51874,17'd51426,17'd17222,17'd20600,17'd16787,17'd15038,17'd51875,17'd27229,17'd51876,17'd51877,17'd10013,17'd10728,17'd27001,17'd11394,17'd16906,17'd51600,17'd51600,17'd51878,17'd51879,17'd51880,17'd22811,17'd12410,17'd51789,17'd13763,17'd12856,17'd12417,17'd12417,17'd13517,17'd12995,17'd13518,17'd21506,17'd15685,17'd50779,17'd12581,17'd17843,17'd18806,17'd18806,17'd22472,17'd23170,17'd24707,17'd26370,17'd29480,17'd30072,17'd31941,17'd31441,17'd34037,17'd35239,17'd50952,17'd51692,17'd51881,17'd50952,17'd31590,17'd33568,17'd30676,17'd29067,17'd29923,17'd25672,17'd25926,17'd18681,17'd11808,17'd10990,17'd10737,17'd10736,17'd14262,17'd11395,17'd11964,17'd13516,17'd11965,17'd11129,17'd14931,17'd11131,17'd16320,17'd16320,17'd11132,17'd13886,17'd13886,17'd10024,17'd16066,17'd8569,17'd33238,17'd28578,17'd15048,17'd26870,17'd17720,17'd10603,17'd19282,17'd19282,17'd11527,17'd11527,17'd11527,17'd14518,17'd10854,17'd16320,17'd20756,17'd28577,17'd16065,17'd10174,17'd15684,17'd9045,17'd9041,17'd24361,17'd24998,17'd16070,17'd25530,17'd15681,17'd22131,17'd9345,17'd9039,17'd29637,17'd50864,17'd12424,17'd9195,17'd24545,17'd21988,17'd51882,17'd51883,17'd51884,17'd51885,17'd51886,17'd51887,17'd51888,17'd51889,17'd23700,17'd51890,17'd5593,17'd51891,17'd51892,17'd51893,17'd51894,17'd51895,17'd21523,17'd51896,17'd51897,17'd51898,17'd51899,17'd51900,17'd51901,17'd51902,17'd43556,17'd46572,17'd51903,17'd51904,17'd51905,17'd51906,17'd51907,17'd24056,17'd51908,17'd51909,17'd51910,17'd51911,17'd51912,17'd51913,17'd51914,17'd50646,17'd50566,17'd49977,17'd46757,17'd49580,17'd51915,17'd48264,17'd49582,17'd50072,17'd50476,17'd49986,17'd49988,17'd49988,17'd50164,17'd50739,17'd50272,17'd51916,17'd48615,17'd45152,17'd39907,17'd51917,17'd28257,17'd29380,17'd29537,17'd51918,17'd26524,17'd28978,17'd33643,17'd38667,17'd23917,17'd29532,17'd23916,17'd24896,17'd28369,17'd28483,17'd27515,17'd46431,17'd33952,17'd33165,17'd38026,17'd28857,17'd49790,17'd31506,17'd31505,17'd31506,17'd31506,17'd31506,17'd33323,17'd49790,17'd30131,17'd30131,17'd30280,17'd30280,17'd49790,17'd30736,17'd51919,17'd40519,17'd44472,17'd46104,17'd48153,17'd49582,17'd50736,17'd50272,17'd51652,17'd51920,17'd43144,17'd42875,17'd49891,17'd39726,17'd41580,17'd39737,17'd51561,17'd46095,17'd25708,17'd28602,17'd25567,17'd25029,17'd24902,17'd32351,17'd22856,17'd31496,17'd35711,17'd32830,17'd30579,17'd38806,17'd29974,17'd30276,17'd22156,17'd48716,17'd51379,17'd21697,17'd22013,17'd31346,17'd48457,17'd42441,17'd51921,17'd51922,17'd51654,17'd51303,17'd34880,17'd36545,17'd36692,17'd33162,17'd51923,17'd51924,17'd49590,17'd51170,17'd51925,17'd51926,17'd51927,17'd51928,17'd23264,17'd11830,17'd5913,17'd5914,17'd6384,17'd5158,17'd6218,17'd8933,17'd8304,17'd6220,17'd25627,17'd4997,17'd33208,17'd51841,17'd7491,17'd51929,17'd4188,17'd28536,17'd30638,17'd32073,17'd34658,17'd32073,17'd6554,17'd30638,17'd25627,17'd5002,17'd5005,17'd4842,17'd28418,17'd5005,17'd30637,17'd25627,17'd5335,17'd28185,17'd28185,17'd28185,17'd5614,17'd6390,17'd9091,17'd29740,17'd34658,17'd51842,17'd50282,17'd36887,17'd5166,17'd42031,17'd5009,17'd37030,17'd36887,17'd51930,17'd5013,17'd38192,17'd51931,17'd4674,17'd51932,17'd51846,17'd3542,17'd51933,17'd51934,17'd51935,17'd51936,17'd51937,17'd51851,17'd40714,17'd51938,17'd51939,17'd41478,17'd51855,17'd41001,17'd51857,17'd18629,17'd10790,17'd18383,17'd5026,17'd11328,17'd4558,17'd4400,17'd4229,17'd4400,17'd4400,17'd4229,17'd3898,17'd5195,17'd3898,17'd3072,17'd5775,17'd628,17'd2113,17'd1114,17'd959,17'd448,17'd8013,17'd51940,17'd30806,17'd20563,17'd214,17'd18515,17'd51582,17'd20265,17'd51858,17'd51859
},
'{
17'd3251,17'd3252,17'd2257,17'd3905,17'd1278,17'd980,17'd28,17'd287,17'd286,17'd1833,17'd467,17'd1691,17'd51860,17'd51941,17'd51766,17'd7388,17'd7061,17'd7060,17'd4430,17'd4430,17'd4431,17'd4091,17'd3755,17'd3755,17'd3754,17'd3754,17'd12335,17'd5210,17'd5806,17'd5806,17'd14192,17'd4581,17'd5058,17'd32089,17'd51942,17'd51943,17'd51944,17'd51945,17'd8055,17'd51865,17'd20141,17'd51946,17'd12800,17'd19252,17'd17095,17'd16764,17'd12357,17'd22802,17'd12527,17'd13093,17'd13209,17'd13209,17'd12357,17'd12062,17'd13461,17'd13461,17'd13460,17'd13460,17'd12212,17'd12212,17'd12212,17'd12212,17'd13596,17'd13596,17'd14620,17'd14763,17'd51866,17'd15383,17'd19005,17'd19005,17'd13093,17'd12530,17'd19006,17'd25512,17'd19385,17'd17319,17'd17318,17'd17318,17'd17318,17'd15765,17'd11231,17'd11088,17'd9158,17'd51947,17'd47870,17'd51948,17'd4124,17'd3628,17'd7584,17'd7914,17'd6777,17'd51771,17'd51949,17'd51101,17'd51773,17'd37971,17'd38093,17'd6948,17'd51775,17'd50932,17'd41646,17'd51777,17'd51950,17'd51588,17'd51680,17'd6951,17'd36766,17'd51951,17'd36197,17'd51591,17'd49615,17'd27965,17'd51952,17'd27111,17'd26860,17'd20443,17'd19272,17'd18072,17'd18316,17'd51953,17'd51954,17'd15166,17'd27228,17'd51955,17'd51785,17'd10015,17'd29917,17'd10844,17'd29939,17'd29634,17'd28567,17'd16197,17'd28097,17'd51956,17'd51879,17'd27978,17'd18803,17'd51957,17'd30982,17'd13643,17'd12418,17'd12417,17'd13517,17'd13517,17'd21506,17'd21506,17'd15685,17'd15685,17'd12719,17'd12581,17'd12582,17'd18806,17'd14258,17'd21362,17'd23168,17'd24856,17'd35376,17'd31286,17'd39211,17'd30973,17'd34037,17'd50111,17'd50952,17'd51958,17'd51959,17'd51692,17'd50863,17'd34037,17'd34835,17'd31440,17'd30370,17'd28343,17'd24538,17'd21361,17'd11397,17'd11808,17'd10989,17'd10989,17'd14262,17'd11395,17'd13762,17'd13516,17'd11965,17'd11129,17'd10854,17'd14931,17'd10990,17'd10854,17'd11524,17'd17236,17'd11399,17'd11527,17'd9190,17'd15428,17'd16066,17'd25814,17'd33083,17'd15048,17'd51960,17'd10606,17'd10991,17'd10991,17'd11527,17'd11527,17'd11527,17'd10476,17'd10854,17'd16320,17'd25928,17'd25530,17'd16065,17'd17716,17'd17123,17'd8883,17'd16066,17'd9041,17'd16795,17'd22814,17'd32916,17'd28577,17'd33722,17'd16554,17'd9346,17'd9039,17'd23860,17'd51961,17'd17607,17'd8731,17'd51962,17'd51963,17'd51964,17'd51965,17'd51966,17'd51967,17'd51968,17'd51969,17'd22312,17'd16090,17'd134,17'd51970,17'd51971,17'd51972,17'd51973,17'd51974,17'd51975,17'd51976,17'd51977,17'd51717,17'd51978,17'd51979,17'd51980,17'd51981,17'd29867,17'd51982,17'd51983,17'd51984,17'd51985,17'd51986,17'd51907,17'd51987,17'd51988,17'd51989,17'd51990,17'd51991,17'd42439,17'd48912,17'd51992,17'd51993,17'd50992,17'd50157,17'd46554,17'd48443,17'd48046,17'd51994,17'd49093,17'd49890,17'd50736,17'd50736,17'd49890,17'd49988,17'd49794,17'd50568,17'd50272,17'd51995,17'd51996,17'd51997,17'd43974,17'd34104,17'd28010,17'd28257,17'd28372,17'd29537,17'd28133,17'd25698,17'd26903,17'd28721,17'd38808,17'd24902,17'd51998,17'd25179,17'd25709,17'd28483,17'd25565,17'd27514,17'd28979,17'd27885,17'd40050,17'd36848,17'd29536,17'd30130,17'd31036,17'd31506,17'd31506,17'd31506,17'd30280,17'd49790,17'd49579,17'd49790,17'd29981,17'd29981,17'd30130,17'd29978,17'd31838,17'd51999,17'd46950,17'd42878,17'd43542,17'd47937,17'd49794,17'd50371,17'd52000,17'd52001,17'd52001,17'd50661,17'd50370,17'd49693,17'd52002,17'd39901,17'd47050,17'd46102,17'd43978,17'd27766,17'd28602,17'd25709,17'd27763,17'd23384,17'd23218,17'd23573,17'd31657,17'd51314,17'd23217,17'd31341,17'd23567,17'd33158,17'd22333,17'd36984,17'd52003,17'd51465,17'd32662,17'd41726,17'd33162,17'd32010,17'd41112,17'd52004,17'd51922,17'd51748,17'd51479,17'd41275,17'd36545,17'd22011,17'd32498,17'd49795,17'd51924,17'd52005,17'd52006,17'd52007,17'd51322,17'd52008,17'd52009,17'd52010,17'd11548,17'd5914,17'd5758,17'd5610,17'd5331,17'd6218,17'd8933,17'd8304,17'd6219,17'd4842,17'd33532,17'd33208,17'd5910,17'd7821,17'd33041,17'd5144,17'd4842,17'd6554,17'd9091,17'd9091,17'd6390,17'd6554,17'd30638,17'd25627,17'd5002,17'd5005,17'd4842,17'd28418,17'd30637,17'd5004,17'd25627,17'd28185,17'd28185,17'd28185,17'd28185,17'd5614,17'd6390,17'd6219,17'd9091,17'd34658,17'd51842,17'd50282,17'd36887,17'd5166,17'd5166,17'd5009,17'd37030,17'd36887,17'd51930,17'd37697,17'd38192,17'd52011,17'd52012,17'd39779,17'd52013,17'd52014,17'd51933,17'd52015,17'd2530,17'd52016,17'd52017,17'd52018,17'd51852,17'd51938,17'd51939,17'd52019,17'd51855,17'd4224,17'd48811,17'd10388,17'd10906,17'd5495,17'd52020,17'd11049,17'd4712,17'd4400,17'd4229,17'd4229,17'd4229,17'd4229,17'd3898,17'd3898,17'd3898,17'd3072,17'd1120,17'd1121,17'd52021,17'd2113,17'd959,17'd448,17'd8013,17'd22435,17'd928,17'd52022,17'd281,17'd1116,17'd20266,17'd52023,17'd52024,17'd30040
},
'{
17'd3251,17'd3252,17'd2257,17'd17,17'd653,17'd980,17'd28,17'd287,17'd286,17'd1833,17'd467,17'd1691,17'd51860,17'd52025,17'd8047,17'd7388,17'd7061,17'd7060,17'd4430,17'd4430,17'd4431,17'd4431,17'd3755,17'd3755,17'd3754,17'd9816,17'd12335,17'd12335,17'd5658,17'd5806,17'd14192,17'd4432,17'd5057,17'd32409,17'd29176,17'd28194,17'd4265,17'd24335,17'd8055,17'd12513,17'd51339,17'd52026,17'd12800,17'd13964,17'd17200,17'd51769,17'd12678,17'd12527,17'd12813,17'd13093,17'd13209,17'd13209,17'd12357,17'd12062,17'd13461,17'd13461,17'd13460,17'd13460,17'd12212,17'd12212,17'd12212,17'd12212,17'd13837,17'd13460,17'd11473,17'd50503,17'd19890,17'd15383,17'd19005,17'd13211,17'd11626,17'd12956,17'd17317,17'd27461,17'd19385,17'd17319,17'd16410,17'd17318,17'd17318,17'd15765,17'd11231,17'd15517,17'd8537,17'd14218,17'd52027,17'd52028,17'd52029,17'd3949,17'd7254,17'd7914,17'd6475,17'd52030,17'd52031,17'd51101,17'd51773,17'd38483,17'd38351,17'd38221,17'd51869,17'd50932,17'd41646,17'd52032,17'd51678,17'd51420,17'd52033,17'd51680,17'd52034,17'd50849,17'd52035,17'd52036,17'd8393,17'd30662,17'd51263,17'd52037,17'd51029,17'd21811,17'd51685,17'd52038,17'd52039,17'd52040,17'd10448,17'd26361,17'd52041,17'd27229,17'd51876,17'd52042,17'd52043,17'd10596,17'd10845,17'd11517,17'd30216,17'd51600,17'd16197,17'd51956,17'd51880,17'd27978,17'd52044,17'd18803,17'd30982,17'd13643,17'd12418,17'd12418,17'd12417,17'd13517,17'd15942,17'd21506,17'd15685,17'd15685,17'd12719,17'd12581,17'd12582,17'd18806,17'd20609,17'd20450,17'd22818,17'd24537,17'd28230,17'd51601,17'd36777,17'd30834,17'd33875,17'd50111,17'd50952,17'd51958,17'd51959,17'd51959,17'd51272,17'd34380,17'd31289,17'd30677,17'd29330,17'd28344,17'd28105,17'd24362,17'd14264,17'd11397,17'd11965,17'd10989,17'd14262,17'd11395,17'd13762,17'd11964,17'd11965,17'd11129,17'd10854,17'd14810,17'd14931,17'd10990,17'd17236,17'd17236,17'd11399,17'd20610,17'd16680,17'd52045,17'd52046,17'd9621,17'd24361,17'd16065,17'd16070,17'd10479,17'd10606,17'd11527,17'd19155,17'd19155,17'd15176,17'd21206,17'd10854,17'd16320,17'd10477,17'd11528,17'd9741,17'd9345,17'd24361,17'd15684,17'd8878,17'd8878,17'd8885,17'd17480,17'd22814,17'd33083,17'd24998,17'd22131,17'd17011,17'd9344,17'd14811,17'd24212,17'd17607,17'd12425,17'd52047,17'd52048,17'd52049,17'd52050,17'd52051,17'd51966,17'd52052,17'd11977,17'd20188,17'd16090,17'd132,17'd11821,17'd52053,17'd20918,17'd52054,17'd52055,17'd52056,17'd52057,17'd52058,17'd52059,17'd52060,17'd52061,17'd52062,17'd52063,17'd52064,17'd51224,17'd52065,17'd52066,17'd52067,17'd52068,17'd52069,17'd21680,17'd52070,17'd52071,17'd52072,17'd21385,17'd52073,17'd36289,17'd52074,17'd52075,17'd52076,17'd50263,17'd46841,17'd47147,17'd48621,17'd48264,17'd50267,17'd51390,17'd50736,17'd50574,17'd49891,17'd49988,17'd49890,17'd51995,17'd51157,17'd52077,17'd41263,17'd44225,17'd41417,17'd40367,17'd28256,17'd28372,17'd29106,17'd29537,17'd27884,17'd25429,17'd27259,17'd28721,17'd29688,17'd52078,17'd52079,17'd28600,17'd28723,17'd33642,17'd25949,17'd27883,17'd29379,17'd28373,17'd49285,17'd29537,17'd29690,17'd30736,17'd31505,17'd31506,17'd31506,17'd31506,17'd30131,17'd49579,17'd49579,17'd49790,17'd29981,17'd29981,17'd36132,17'd31038,17'd29981,17'd50657,17'd52080,17'd50469,17'd48701,17'd48909,17'd50164,17'd50371,17'd51652,17'd52001,17'd51741,17'd50072,17'd50271,17'd52081,17'd52082,17'd51082,17'd48524,17'd48258,17'd32658,17'd27766,17'd28720,17'd27512,17'd28129,17'd29827,17'd39131,17'd36009,17'd51747,17'd35018,17'd29829,17'd34112,17'd29829,17'd30277,17'd22159,17'd36128,17'd45890,17'd52083,17'd31831,17'd32997,17'd48457,17'd34280,17'd46339,17'd52084,17'd51922,17'd52085,17'd52086,17'd34280,17'd36545,17'd48457,17'd21693,17'd48456,17'd46341,17'd45885,17'd30468,17'd52087,17'd52088,17'd52089,17'd52090,17'd52091,17'd10627,17'd50670,17'd5481,17'd4844,17'd6389,17'd26709,17'd8303,17'd8154,17'd27935,17'd31716,17'd38846,17'd5604,17'd52092,17'd52093,17'd33367,17'd42910,17'd5004,17'd6390,17'd9091,17'd9091,17'd6390,17'd6554,17'd30638,17'd30333,17'd5004,17'd5005,17'd4842,17'd28418,17'd30637,17'd5004,17'd30333,17'd28185,17'd28185,17'd28185,17'd28185,17'd5614,17'd6390,17'd9091,17'd32074,17'd34658,17'd52094,17'd50282,17'd36887,17'd5166,17'd5166,17'd5163,17'd37030,17'd36887,17'd51930,17'd37697,17'd52095,17'd49997,17'd52096,17'd39779,17'd52013,17'd52014,17'd52097,17'd52098,17'd52099,17'd52100,17'd52017,17'd52101,17'd52102,17'd51938,17'd3212,17'd52019,17'd51855,17'd4224,17'd41315,17'd41003,17'd10388,17'd18142,17'd52020,17'd11049,17'd4712,17'd4400,17'd4229,17'd4229,17'd4229,17'd4229,17'd3898,17'd3898,17'd3898,17'd1402,17'd628,17'd1121,17'd52103,17'd52021,17'd959,17'd629,17'd52104,17'd22606,17'd52105,17'd52106,17'd790,17'd787,17'd52107,17'd38073,17'd52024,17'd52108
},
'{
17'd3251,17'd3252,17'd2257,17'd3905,17'd1278,17'd980,17'd6744,17'd6902,17'd286,17'd467,17'd1691,17'd1691,17'd7384,17'd51941,17'd52025,17'd7555,17'd7061,17'd7060,17'd4430,17'd4430,17'd4430,17'd4430,17'd4091,17'd4091,17'd3755,17'd3907,17'd11210,17'd5657,17'd5806,17'd5806,17'd14192,17'd4581,17'd5058,17'd4585,17'd5064,17'd5390,17'd51863,17'd24335,17'd8055,17'd12513,17'd51339,17'd52109,17'd52110,17'd13964,17'd17315,17'd16764,17'd12357,17'd15763,17'd12527,17'd13093,17'd13209,17'd13209,17'd12357,17'd12062,17'd13461,17'd13461,17'd13460,17'd13460,17'd14620,17'd14620,17'd13837,17'd13837,17'd13837,17'd13596,17'd14620,17'd50503,17'd19890,17'd19005,17'd13599,17'd13599,17'd12527,17'd12218,17'd18884,17'd19007,17'd19008,17'd19255,17'd16410,17'd17318,17'd17572,17'd11231,17'd15765,17'd15765,17'd9702,17'd9007,17'd52027,17'd52111,17'd52029,17'd3949,17'd7254,17'd7914,17'd6475,17'd41780,17'd52031,17'd52112,17'd52113,17'd38483,17'd52114,17'd38351,17'd51869,17'd6646,17'd40585,17'd52032,17'd41784,17'd50764,17'd51588,17'd51680,17'd38487,17'd52115,17'd52116,17'd52117,17'd52118,17'd52119,17'd27722,17'd52120,17'd52121,17'd52122,17'd20443,17'd17956,17'd20896,17'd52123,17'd51953,17'd51954,17'd52124,17'd26995,17'd51955,17'd27734,17'd10724,17'd10157,17'd30093,17'd35245,17'd52125,17'd52126,17'd52127,17'd52128,17'd28097,17'd52129,17'd14925,17'd19530,17'd52130,17'd13643,17'd13643,17'd14525,17'd14003,17'd12417,17'd13517,17'd15570,17'd15685,17'd15685,17'd12106,17'd17603,17'd18917,17'd12582,17'd20609,17'd52131,17'd20449,17'd23512,17'd27004,17'd30525,17'd47107,17'd39211,17'd34203,17'd31590,17'd50952,17'd51958,17'd52132,17'd52133,17'd52134,17'd51432,17'd34203,17'd34835,17'd31440,17'd28461,17'd28227,17'd24707,17'd22992,17'd16326,17'd24029,17'd24029,17'd11397,17'd11396,17'd11395,17'd11395,17'd10989,17'd11965,17'd11130,17'd11275,17'd11274,17'd14673,17'd11274,17'd11274,17'd11274,17'd13138,17'd21205,17'd23679,17'd15050,17'd21507,17'd9040,17'd10174,17'd18556,17'd11135,17'd20756,17'd20756,17'd17599,17'd19155,17'd12423,17'd11399,17'd10990,17'd10737,17'd10604,17'd14666,17'd11134,17'd10857,17'd9190,17'd23859,17'd29920,17'd9046,17'd12425,17'd8729,17'd25677,17'd17480,17'd16065,17'd33722,17'd17839,17'd9741,17'd10026,17'd10336,17'd9194,17'd8569,17'd37334,17'd8887,17'd52135,17'd52136,17'd52137,17'd51883,17'd52138,17'd52139,17'd52140,17'd17363,17'd51890,17'd11683,17'd52141,17'd52142,17'd52143,17'd52144,17'd52145,17'd52146,17'd52147,17'd52148,17'd52149,17'd52150,17'd52151,17'd52152,17'd52153,17'd22492,17'd52154,17'd52155,17'd52156,17'd5593,17'd131,17'd52157,17'd52158,17'd52159,17'd51375,17'd52160,17'd43158,17'd24094,17'd52161,17'd52162,17'd51554,17'd52163,17'd47237,17'd47044,17'd49089,17'd49484,17'd50468,17'd50268,17'd50072,17'd49985,17'd49891,17'd49891,17'd49986,17'd51157,17'd50160,17'd52164,17'd52165,17'd44356,17'd41731,17'd32193,17'd28257,17'd28372,17'd28857,17'd29537,17'd31503,17'd26782,17'd27515,17'd28600,17'd29100,17'd52166,17'd28717,17'd31351,17'd28978,17'd28724,17'd26530,17'd26782,17'd27761,17'd28487,17'd36848,17'd28857,17'd29979,17'd30736,17'd31505,17'd33489,17'd31506,17'd33489,17'd30131,17'd49579,17'd32833,17'd32508,17'd29981,17'd29981,17'd36132,17'd49286,17'd29833,17'd52167,17'd47630,17'd39431,17'd52168,17'd48263,17'd49986,17'd52000,17'd51745,17'd52169,17'd51830,17'd50468,17'd49988,17'd52170,17'd40214,17'd40048,17'd50070,17'd43155,17'd28723,17'd28602,17'd27765,17'd24897,17'd29378,17'd32191,17'd31656,17'd35429,17'd39911,17'd39131,17'd24421,17'd31029,17'd29829,17'd36986,17'd22162,17'd41865,17'd52003,17'd52171,17'd31345,17'd31831,17'd42150,17'd52172,17'd52173,17'd52174,17'd51922,17'd52175,17'd52172,17'd51912,17'd22864,17'd22510,17'd42150,17'd48630,17'd46218,17'd52176,17'd50075,17'd52177,17'd52178,17'd52179,17'd52180,17'd52181,17'd10198,17'd50670,17'd5481,17'd4844,17'd6553,17'd26709,17'd8154,17'd6707,17'd25627,17'd4996,17'd38846,17'd33041,17'd51574,17'd33041,17'd5144,17'd4841,17'd30638,17'd6219,17'd9091,17'd9091,17'd6219,17'd6554,17'd28185,17'd25627,17'd5002,17'd5005,17'd5005,17'd4842,17'd5004,17'd5004,17'd30638,17'd28185,17'd28185,17'd30638,17'd28185,17'd5614,17'd26709,17'd8303,17'd9091,17'd34658,17'd36586,17'd31717,17'd30638,17'd25627,17'd5160,17'd25627,17'd37030,17'd52182,17'd37435,17'd37944,17'd51326,17'd52183,17'd52184,17'd52185,17'd52186,17'd52187,17'd52188,17'd52189,17'd37706,17'd52190,17'd52017,17'd52191,17'd52192,17'd51938,17'd52193,17'd50182,17'd52194,17'd4224,17'd41315,17'd48559,17'd18383,17'd18142,17'd52020,17'd11049,17'd4712,17'd4229,17'd1824,17'd1824,17'd1824,17'd1824,17'd3898,17'd5195,17'd3898,17'd1402,17'd796,17'd630,17'd1546,17'd2113,17'd796,17'd629,17'd52104,17'd52195,17'd52196,17'd33539,17'd18633,17'd20266,17'd52197,17'd28427,17'd52108,17'd52198
},
'{
17'd3251,17'd3252,17'd2257,17'd17,17'd653,17'd980,17'd6744,17'd6902,17'd286,17'd1833,17'd467,17'd1691,17'd7384,17'd1690,17'd8047,17'd7555,17'd7061,17'd7060,17'd4430,17'd4430,17'd4430,17'd4430,17'd4431,17'd4091,17'd3755,17'd3907,17'd11210,17'd3756,17'd5658,17'd5806,17'd14192,17'd4742,17'd5218,17'd32409,17'd29176,17'd5390,17'd51863,17'd52199,17'd52200,17'd52201,17'd20284,17'd12939,17'd12516,17'd16649,17'd17315,17'd51769,17'd12678,17'd15516,17'd12527,17'd12813,17'd13209,17'd13092,17'd12357,17'd12062,17'd13461,17'd13461,17'd14216,17'd13460,17'd13460,17'd14620,17'd13837,17'd13837,17'd13837,17'd14620,17'd11473,17'd50503,17'd13210,17'd19005,17'd13599,17'd13599,17'd12527,17'd12065,17'd12531,17'd17689,17'd19383,17'd19255,17'd11231,17'd17318,17'd17572,17'd11231,17'd15765,17'd15517,17'd7418,17'd9007,17'd52202,17'd52203,17'd52029,17'd4462,17'd3949,17'd7584,17'd7094,17'd6474,17'd52204,17'd52112,17'd52113,17'd52205,17'd38483,17'd52206,17'd52207,17'd39058,17'd40585,17'd41176,17'd41647,17'd50394,17'd51588,17'd52033,17'd38487,17'd37188,17'd52208,17'd52209,17'd33395,17'd8393,17'd28929,17'd52210,17'd22805,17'd20598,17'd52211,17'd52212,17'd52213,17'd52039,17'd51595,17'd52214,17'd26361,17'd26865,17'd52215,17'd52216,17'd10153,17'd10462,17'd30386,17'd52217,17'd10847,17'd25277,17'd27852,17'd52128,17'd17008,17'd52218,17'd52219,17'd52044,17'd51957,17'd18684,17'd13643,17'd14525,17'd12416,17'd14003,17'd13517,17'd15570,17'd15685,17'd15685,17'd12106,17'd12106,17'd18917,17'd12582,17'd20609,17'd52220,17'd52221,17'd23514,17'd27347,17'd27346,17'd30830,17'd30527,17'd31941,17'd31590,17'd50952,17'd51958,17'd52132,17'd51959,17'd51693,17'd52134,17'd34380,17'd31288,17'd31765,17'd31587,17'd29328,17'd26872,17'd24209,17'd18443,17'd21985,17'd24029,17'd11397,17'd11397,17'd11395,17'd11395,17'd14262,17'd10989,17'd11130,17'd14381,17'd11275,17'd14673,17'd11274,17'd14673,17'd16068,17'd16068,17'd17236,17'd11134,17'd15682,17'd21507,17'd8879,17'd17607,17'd10026,17'd19531,17'd16070,17'd15688,17'd17599,17'd27488,17'd12584,17'd11398,17'd14931,17'd11519,17'd14810,17'd14810,17'd14666,17'd11528,17'd9341,17'd17600,17'd9621,17'd23861,17'd16205,17'd11966,17'd11966,17'd9195,17'd24361,17'd16065,17'd9739,17'd9739,17'd9620,17'd9743,17'd9040,17'd8723,17'd22473,17'd15429,17'd52222,17'd52223,17'd52224,17'd52225,17'd52226,17'd52227,17'd52228,17'd7979,17'd20628,17'd52229,17'd52230,17'd52231,17'd52232,17'd52233,17'd52234,17'd52235,17'd52236,17'd52237,17'd52238,17'd52239,17'd52240,17'd52241,17'd21381,17'd52242,17'd52243,17'd52244,17'd52245,17'd132,17'd52246,17'd52247,17'd52248,17'd52249,17'd52250,17'd52251,17'd33649,17'd52252,17'd50647,17'd49171,17'd52253,17'd52254,17'd52255,17'd52256,17'd43419,17'd49794,17'd50160,17'd50736,17'd50574,17'd50271,17'd49987,17'd49985,17'd50268,17'd51831,17'd51916,17'd48900,17'd44223,17'd43289,17'd32831,17'd36988,17'd29380,17'd28728,17'd29536,17'd28487,17'd29245,17'd27259,17'd27514,17'd28598,17'd52257,17'd52258,17'd38538,17'd32343,17'd27146,17'd27640,17'd43290,17'd28727,17'd28256,17'd29537,17'd29536,17'd30884,17'd49790,17'd30736,17'd31506,17'd33489,17'd33489,17'd33489,17'd49790,17'd49579,17'd32833,17'd29981,17'd29981,17'd29981,17'd36132,17'd36848,17'd49791,17'd36841,17'd52259,17'd39735,17'd49279,17'd49184,17'd50072,17'd51652,17'd51834,17'd52169,17'd51157,17'd49788,17'd49485,17'd48360,17'd39736,17'd46952,17'd52260,17'd43286,17'd28602,17'd28720,17'd25438,17'd29240,17'd23385,17'd29973,17'd35018,17'd40052,17'd31656,17'd32351,17'd23734,17'd23734,17'd30579,17'd22331,17'd22156,17'd52261,17'd52261,17'd36544,17'd31497,17'd31660,17'd34617,17'd51479,17'd46776,17'd52262,17'd52084,17'd46455,17'd41275,17'd43697,17'd42150,17'd22511,17'd48453,17'd47540,17'd52263,17'd52264,17'd51567,17'd52265,17'd52266,17'd39300,17'd52267,17'd50584,17'd29292,17'd52268,17'd4844,17'd5612,17'd8303,17'd26709,17'd8154,17'd6387,17'd4686,17'd4997,17'd5477,17'd4521,17'd52269,17'd4188,17'd5327,17'd30637,17'd28185,17'd6219,17'd7499,17'd9091,17'd6219,17'd6390,17'd28185,17'd30333,17'd25627,17'd5002,17'd5005,17'd30637,17'd5004,17'd30333,17'd30638,17'd28185,17'd28185,17'd30638,17'd28185,17'd5614,17'd8303,17'd8933,17'd29740,17'd34658,17'd36586,17'd6554,17'd30638,17'd25627,17'd5160,17'd30638,17'd52270,17'd35760,17'd37435,17'd52271,17'd51248,17'd52272,17'd52184,17'd50674,17'd52273,17'd52187,17'd52274,17'd42920,17'd21782,17'd52190,17'd52017,17'd52275,17'd2729,17'd51938,17'd52193,17'd52276,17'd41000,17'd4224,17'd41002,17'd41626,17'd10388,17'd5026,17'd52020,17'd11049,17'd4712,17'd4229,17'd1824,17'd1824,17'd1824,17'd1824,17'd3898,17'd5195,17'd1824,17'd38071,17'd38856,17'd18144,17'd796,17'd2113,17'd796,17'd8314,17'd8788,17'd929,17'd52106,17'd25495,17'd32559,17'd766,17'd19602,17'd52277,17'd52278,17'd52279
},
'{
17'd34512,17'd14070,17'd2257,17'd3905,17'd980,17'd980,17'd286,17'd286,17'd286,17'd467,17'd1691,17'd1691,17'd1691,17'd1690,17'd7555,17'd7555,17'd7061,17'd7060,17'd6744,17'd4430,17'd4430,17'd4430,17'd4431,17'd4091,17'd3755,17'd3907,17'd11210,17'd5657,17'd5806,17'd5806,17'd5806,17'd4742,17'd5218,17'd4585,17'd25650,17'd5390,17'd51863,17'd52199,17'd52200,17'd52201,17'd20284,17'd12664,17'd52280,17'd15508,17'd52281,17'd16763,17'd15762,17'd12678,17'd12678,17'd13092,17'd13209,17'd13092,17'd12357,17'd12062,17'd13461,17'd13461,17'd14216,17'd14216,17'd13460,17'd14620,17'd14620,17'd14620,17'd13837,17'd13837,17'd13460,17'd50503,17'd13210,17'd19005,17'd13599,17'd13599,17'd12527,17'd12065,17'd12531,17'd19893,17'd19383,17'd19255,17'd11231,17'd17318,17'd20425,17'd11231,17'd15765,17'd15765,17'd46366,17'd9007,17'd52282,17'd52283,17'd52284,17'd4122,17'd3783,17'd7584,17'd7914,17'd6474,17'd6479,17'd52112,17'd52285,17'd52286,17'd52205,17'd52114,17'd38351,17'd6645,17'd40274,17'd41176,17'd41647,17'd50394,17'd51588,17'd52287,17'd38894,17'd52288,17'd52289,17'd52290,17'd50297,17'd32428,17'd28329,17'd51263,17'd22805,17'd26249,17'd22123,17'd52291,17'd17956,17'd52292,17'd17114,17'd51507,17'd26748,17'd15416,17'd52293,17'd52294,17'd10969,17'd10724,17'd10157,17'd26868,17'd10982,17'd52128,17'd27852,17'd11955,17'd12103,17'd52295,17'd52296,17'd52297,17'd52298,17'd18322,17'd30231,17'd52299,17'd14525,17'd14525,17'd12417,17'd15570,17'd15433,17'd15433,17'd12106,17'd12106,17'd15053,17'd18917,17'd12582,17'd20047,17'd52131,17'd26035,17'd23682,17'd25672,17'd28816,17'd30831,17'd31761,17'd31442,17'd50863,17'd52300,17'd52301,17'd52302,17'd52303,17'd52304,17'd52305,17'd34380,17'd34203,17'd30221,17'd29067,17'd28229,17'd25925,17'd21505,17'd23169,17'd21985,17'd11397,17'd11397,17'd14673,17'd16068,17'd14810,17'd14810,17'd10854,17'd14132,17'd22647,17'd11274,17'd14673,17'd14673,17'd16068,17'd16069,17'd14262,17'd13886,17'd9344,17'd10027,17'd24368,17'd26259,17'd9042,17'd10173,17'd15048,17'd14928,17'd19642,17'd19155,17'd14134,17'd11524,17'd14673,17'd11395,17'd16068,17'd14673,17'd12862,17'd52306,17'd15943,17'd10857,17'd28820,17'd9045,17'd26038,17'd12425,17'd8412,17'd24368,17'd9041,17'd10174,17'd16554,17'd9619,17'd16554,17'd13887,17'd8875,17'd8723,17'd8878,17'd10338,17'd8412,17'd8576,17'd11406,17'd19035,17'd52307,17'd52308,17'd52309,17'd52310,17'd23017,17'd52311,17'd52312,17'd52313,17'd52314,17'd52315,17'd23886,17'd51537,17'd52316,17'd52317,17'd52318,17'd52319,17'd52320,17'd52321,17'd52322,17'd52323,17'd20768,17'd5593,17'd135,17'd132,17'd20465,17'd52311,17'd52324,17'd52325,17'd52326,17'd42003,17'd52327,17'd52328,17'd52329,17'd50461,17'd52330,17'd52331,17'd52332,17'd40516,17'd49691,17'd50072,17'd50272,17'd50273,17'd50574,17'd50271,17'd49985,17'd50736,17'd50371,17'd52333,17'd52334,17'd48356,17'd39583,17'd37777,17'd32505,17'd37118,17'd30587,17'd28728,17'd29536,17'd28257,17'd30586,17'd25833,17'd26062,17'd39444,17'd52335,17'd27764,17'd52336,17'd34637,17'd27027,17'd33499,17'd26781,17'd27642,17'd28487,17'd29831,17'd29536,17'd29690,17'd30131,17'd31506,17'd33489,17'd33489,17'd30131,17'd30131,17'd29979,17'd29690,17'd32833,17'd29981,17'd29981,17'd29981,17'd29981,17'd36989,17'd52337,17'd52338,17'd52339,17'd52340,17'd48535,17'd49691,17'd50268,17'd51920,17'd52341,17'd52342,17'd50371,17'd49794,17'd49183,17'd51557,17'd47725,17'd49476,17'd52343,17'd37778,17'd28720,17'd27765,17'd28254,17'd28849,17'd32191,17'd41419,17'd39911,17'd40052,17'd30129,17'd23567,17'd29241,17'd23920,17'd23569,17'd30276,17'd22165,17'd52261,17'd31832,17'd41726,17'd31497,17'd33162,17'd52344,17'd52345,17'd52346,17'd21385,17'd52347,17'd46571,17'd51302,17'd43697,17'd50827,17'd22337,17'd48538,17'd47447,17'd52348,17'd47353,17'd52349,17'd51752,17'd52350,17'd52351,17'd46125,17'd46227,17'd7660,17'd52352,17'd4844,17'd5331,17'd8303,17'd50486,17'd6707,17'd5760,17'd4995,17'd4187,17'd5477,17'd4990,17'd4188,17'd5145,17'd28418,17'd30333,17'd6390,17'd7499,17'd6220,17'd6219,17'd6219,17'd6390,17'd28185,17'd30638,17'd25627,17'd5004,17'd5004,17'd5004,17'd5160,17'd30638,17'd28185,17'd6554,17'd6554,17'd31717,17'd6554,17'd6390,17'd8303,17'd8154,17'd7499,17'd32074,17'd32073,17'd6554,17'd30638,17'd5004,17'd30638,17'd30638,17'd50282,17'd35760,17'd37435,17'd52095,17'd51177,17'd52353,17'd52354,17'd52355,17'd51847,17'd36742,17'd52356,17'd52357,17'd52358,17'd52359,17'd52360,17'd52275,17'd52361,17'd52362,17'd52193,17'd50182,17'd40861,17'd5626,17'd41002,17'd18512,17'd18383,17'd5026,17'd52020,17'd11049,17'd5195,17'd1824,17'd1824,17'd1824,17'd1825,17'd1825,17'd1824,17'd3898,17'd1402,17'd447,17'd236,17'd630,17'd959,17'd959,17'd235,17'd52363,17'd38332,17'd1664,17'd52364,17'd52365,17'd52366,17'd52107,17'd52023,17'd52367,17'd52368,17'd52369
},
'{
17'd34512,17'd14070,17'd2257,17'd17,17'd652,17'd27,17'd286,17'd1833,17'd286,17'd1833,17'd467,17'd1691,17'd1691,17'd1691,17'd7555,17'd7385,17'd7061,17'd7060,17'd6744,17'd4430,17'd4430,17'd4430,17'd4431,17'd4431,17'd3755,17'd3755,17'd11210,17'd3756,17'd5658,17'd5806,17'd5806,17'd4742,17'd5218,17'd32409,17'd25502,17'd51862,17'd28194,17'd52370,17'd7234,17'd21481,17'd50501,17'd22796,17'd12345,17'd20420,17'd17933,17'd17685,17'd16282,17'd12678,17'd12678,17'd13092,17'd13092,17'd13092,17'd12357,17'd12062,17'd13461,17'd13461,17'd14466,17'd14216,17'd13460,17'd14620,17'd14620,17'd14620,17'd13837,17'd14620,17'd12526,17'd50503,17'd13210,17'd19005,17'd13599,17'd13599,17'd12527,17'd12065,17'd20424,17'd19893,17'd19383,17'd19255,17'd15765,17'd16410,17'd20425,17'd11231,17'd15765,17'd10429,17'd8537,17'd9007,17'd52371,17'd52372,17'd52373,17'd52374,17'd4128,17'd52375,17'd7254,17'd7913,17'd6776,17'd51949,17'd52285,17'd6641,17'd52376,17'd52377,17'd52378,17'd39200,17'd40428,17'd52379,17'd50504,17'd52380,17'd50764,17'd51420,17'd40429,17'd52381,17'd52382,17'd52383,17'd50297,17'd33395,17'd51423,17'd52384,17'd26991,17'd26249,17'd52122,17'd52385,17'd10302,17'd52386,17'd52387,17'd52388,17'd52389,17'd52390,17'd52391,17'd52392,17'd10968,17'd52393,17'd10462,17'd52394,17'd52395,17'd52396,17'd27852,17'd28455,17'd11126,17'd11125,17'd52397,17'd19640,17'd52398,17'd52399,17'd30983,17'd31774,17'd14930,17'd14930,17'd12417,17'd13517,17'd15433,17'd15433,17'd12106,17'd12106,17'd15053,17'd18917,17'd12582,17'd18806,17'd52220,17'd20450,17'd23514,17'd24859,17'd26370,17'd30218,17'd39211,17'd31442,17'd50863,17'd50952,17'd52400,17'd52401,17'd52402,17'd52303,17'd51272,17'd51118,17'd33875,17'd48660,17'd31439,17'd31768,17'd26757,17'd24030,17'd22472,17'd18327,17'd21985,17'd24029,17'd11274,17'd14673,17'd14810,17'd14810,17'd14810,17'd11131,17'd14381,17'd11275,17'd16068,17'd14673,17'd14673,17'd11520,17'd13362,17'd12720,17'd14383,17'd9045,17'd8412,17'd11966,17'd8878,17'd10336,17'd15187,17'd9619,17'd14928,17'd19642,17'd15176,17'd11399,17'd11274,17'd14262,17'd11522,17'd11521,17'd16069,17'd12720,17'd17121,17'd16908,17'd16319,17'd52403,17'd15684,17'd25677,17'd24368,17'd9886,17'd10338,17'd9041,17'd15430,17'd15180,17'd28815,17'd18080,17'd16318,17'd9044,17'd9621,17'd8878,17'd8725,17'd8413,17'd25679,17'd52404,17'd52405,17'd52307,17'd52406,17'd52407,17'd24877,17'd52408,17'd52409,17'd22148,17'd52410,17'd51715,17'd52411,17'd52412,17'd52413,17'd21073,17'd52414,17'd52415,17'd52416,17'd52417,17'd52418,17'd52419,17'd11683,17'd360,17'd130,17'd5593,17'd51987,17'd52420,17'd52421,17'd52422,17'd46967,17'd22512,17'd52423,17'd52424,17'd52425,17'd52426,17'd51234,17'd52427,17'd52428,17'd41410,17'd49986,17'd51163,17'd51163,17'd50273,17'd50370,17'd49985,17'd50574,17'd51157,17'd50736,17'd49787,17'd42293,17'd44223,17'd43289,17'd35570,17'd29248,17'd33656,17'd30587,17'd52429,17'd29537,17'd28133,17'd27258,17'd25708,17'd26064,17'd52430,17'd52431,17'd33156,17'd32005,17'd30735,17'd26902,17'd35023,17'd29379,17'd28373,17'd36848,17'd29978,17'd29690,17'd49579,17'd33489,17'd31506,17'd33489,17'd31506,17'd30131,17'd30131,17'd29979,17'd29690,17'd32508,17'd29981,17'd31037,17'd29981,17'd31037,17'd32018,17'd35150,17'd52432,17'd52433,17'd52434,17'd49091,17'd49683,17'd51830,17'd52169,17'd52435,17'd52342,17'd50272,17'd49988,17'd49091,17'd52436,17'd40676,17'd46203,17'd43155,17'd32996,17'd28720,17'd28369,17'd24745,17'd29972,17'd23217,17'd31656,17'd22858,17'd39742,17'd39278,17'd31502,17'd23731,17'd31033,17'd32351,17'd22681,17'd46551,17'd22003,17'd31660,17'd49488,17'd31344,17'd32498,17'd52437,17'd52438,17'd52439,17'd51980,17'd51394,17'd42747,17'd34881,17'd42150,17'd52440,17'd32187,17'd48452,17'd46574,17'd52441,17'd52442,17'd52443,17'd51839,17'd37929,17'd19836,17'd52444,17'd52445,17'd8914,17'd52446,17'd52352,17'd5332,17'd50486,17'd50486,17'd6707,17'd5758,17'd5145,17'd52269,17'd5477,17'd33367,17'd5144,17'd5327,17'd30637,17'd31717,17'd9091,17'd7668,17'd6391,17'd6220,17'd6219,17'd6390,17'd28185,17'd30638,17'd25627,17'd25627,17'd25627,17'd31553,17'd28185,17'd28185,17'd6554,17'd6390,17'd6554,17'd6554,17'd6554,17'd6219,17'd8303,17'd8304,17'd7499,17'd32074,17'd32073,17'd6554,17'd30638,17'd5004,17'd30638,17'd30638,17'd50282,17'd5920,17'd5339,17'd52447,17'd51010,17'd52448,17'd52449,17'd52450,17'd52451,17'd52452,17'd52453,17'd52454,17'd52455,17'd52456,17'd52457,17'd52458,17'd52459,17'd52362,17'd52460,17'd52276,17'd41000,17'd5626,17'd45185,17'd41626,17'd10388,17'd5026,17'd52020,17'd11049,17'd5195,17'd1824,17'd1825,17'd1825,17'd1825,17'd1825,17'd1824,17'd1824,17'd1402,17'd796,17'd52461,17'd18144,17'd628,17'd959,17'd235,17'd52462,17'd38332,17'd34510,17'd20562,17'd52463,17'd764,17'd52464,17'd52465,17'd30040,17'd1521,17'd52466
},
'{
17'd35619,17'd3101,17'd2426,17'd17,17'd653,17'd1278,17'd286,17'd286,17'd286,17'd285,17'd1832,17'd1691,17'd1690,17'd1690,17'd8047,17'd7728,17'd7061,17'd7060,17'd7060,17'd27444,17'd4430,17'd4430,17'd4431,17'd4431,17'd3755,17'd3907,17'd11210,17'd5657,17'd5806,17'd5806,17'd5806,17'd4742,17'd5058,17'd4586,17'd30048,17'd5526,17'd28194,17'd6607,17'd52467,17'd50500,17'd24514,17'd20285,17'd12345,17'd20420,17'd17933,17'd16654,17'd17571,17'd15762,17'd12677,17'd12678,17'd13092,17'd13092,17'd12357,17'd12062,17'd50503,17'd50503,17'd13461,17'd13461,17'd13460,17'd14620,17'd14620,17'd13460,17'd13460,17'd52468,17'd11473,17'd50503,17'd13599,17'd19005,17'd13210,17'd13209,17'd19127,17'd12679,17'd12362,17'd19006,17'd19511,17'd17206,17'd16766,17'd17205,17'd18174,17'd16766,17'd15765,17'd15765,17'd46366,17'd9703,17'd52469,17'd52470,17'd52471,17'd52472,17'd4293,17'd52375,17'd7584,17'd7913,17'd7092,17'd6479,17'd52112,17'd52473,17'd52474,17'd52205,17'd51773,17'd52475,17'd39649,17'd48191,17'd42215,17'd52380,17'd41784,17'd50765,17'd52033,17'd51258,17'd52476,17'd52477,17'd37597,17'd50197,17'd52478,17'd27840,17'd9322,17'd9595,17'd52479,17'd52211,17'd10137,17'd52480,17'd21812,17'd16786,17'd52481,17'd16056,17'd51875,17'd27614,17'd27975,17'd10969,17'd10156,17'd11270,17'd11516,17'd52395,17'd52482,17'd27732,17'd17120,17'd12248,17'd52483,17'd22990,17'd52484,17'd52485,17'd33247,17'd30378,17'd14523,17'd14523,17'd14525,17'd21057,17'd15570,17'd15433,17'd15433,17'd15685,17'd12719,17'd12581,17'd15053,17'd18806,17'd19411,17'd19410,17'd20608,17'd23170,17'd26149,17'd28343,17'd34551,17'd30834,17'd34037,17'd50863,17'd52300,17'd51958,17'd52302,17'd52303,17'd51693,17'd51513,17'd35239,17'd33720,17'd31941,17'd31440,17'd28345,17'd28570,17'd24362,17'd16442,17'd22817,17'd19533,17'd11808,17'd14931,17'd24860,17'd17121,17'd14810,17'd10990,17'd14263,17'd14132,17'd10854,17'd12720,17'd12862,17'd14262,17'd12861,17'd14262,17'd48406,17'd14674,17'd8879,17'd8571,17'd8724,17'd24999,17'd9190,17'd9480,17'd18556,17'd11671,17'd20756,17'd13886,17'd11274,17'd11964,17'd11396,17'd11521,17'd11667,17'd11962,17'd16797,17'd29331,17'd29332,17'd25675,17'd52486,17'd9621,17'd8886,17'd16205,17'd11966,17'd30217,17'd8726,17'd29637,17'd28964,17'd28815,17'd19279,17'd16328,17'd9189,17'd9040,17'd22473,17'd15945,17'd15945,17'd25679,17'd17241,17'd16078,17'd52487,17'd52488,17'd52489,17'd52490,17'd52491,17'd20626,17'd52492,17'd20768,17'd20774,17'd52493,17'd52494,17'd52495,17'd21223,17'd52496,17'd52497,17'd21224,17'd20768,17'd52069,17'd131,17'd128,17'd132,17'd5593,17'd52498,17'd52499,17'd52249,17'd52500,17'd52004,17'd52501,17'd52502,17'd52503,17'd49376,17'd49274,17'd52504,17'd48442,17'd52505,17'd49988,17'd50476,17'd52000,17'd51163,17'd42874,17'd52506,17'd50574,17'd50272,17'd51157,17'd52507,17'd48154,17'd51159,17'd44593,17'd37658,17'd28373,17'd28371,17'd30587,17'd28371,17'd52429,17'd28487,17'd26278,17'd28853,17'd38538,17'd28720,17'd52430,17'd52508,17'd40520,17'd36690,17'd26902,17'd28853,17'd26781,17'd28854,17'd29537,17'd31038,17'd29979,17'd29690,17'd30131,17'd31506,17'd31506,17'd33323,17'd34117,17'd30131,17'd49790,17'd29690,17'd29690,17'd34114,17'd29833,17'd29981,17'd32508,17'd33167,17'd37250,17'd40366,17'd52509,17'd52510,17'd52168,17'd43419,17'd50468,17'd51741,17'd52511,17'd52512,17'd52511,17'd50739,17'd49485,17'd48359,17'd52513,17'd46661,17'd48612,17'd43550,17'd28721,17'd28600,17'd25177,17'd29100,17'd29830,17'd32827,17'd36009,17'd39911,17'd33949,17'd29829,17'd29241,17'd24249,17'd30275,17'd46966,17'd33944,17'd32012,17'd33798,17'd31345,17'd49488,17'd31345,17'd32010,17'd51551,17'd52346,17'd52514,17'd51980,17'd46455,17'd52172,17'd22511,17'd22510,17'd50818,17'd52515,17'd48162,17'd23045,17'd52516,17'd52517,17'd50581,17'd52518,17'd52519,17'd25871,17'd52520,17'd12740,17'd52521,17'd9217,17'd5914,17'd5916,17'd8303,17'd8303,17'd6387,17'd5326,17'd33367,17'd52269,17'd4990,17'd33367,17'd5153,17'd28418,17'd30333,17'd6554,17'd9091,17'd7499,17'd6220,17'd6390,17'd6390,17'd6554,17'd28185,17'd30638,17'd5160,17'd5160,17'd30333,17'd30333,17'd30638,17'd31717,17'd6554,17'd6390,17'd6390,17'd6390,17'd6219,17'd6219,17'd8304,17'd8304,17'd7499,17'd32073,17'd6554,17'd6554,17'd30638,17'd5004,17'd30638,17'd37030,17'd52182,17'd36311,17'd5171,17'd52522,17'd38321,17'd52523,17'd52524,17'd52525,17'd52526,17'd52527,17'd52528,17'd52529,17'd52530,17'd52531,17'd52532,17'd2547,17'd52459,17'd52533,17'd41314,17'd50182,17'd52194,17'd4055,17'd41315,17'd48559,17'd18383,17'd18142,17'd52020,17'd5497,17'd3898,17'd3898,17'd3426,17'd1825,17'd1825,17'd1824,17'd2558,17'd2558,17'd4059,17'd960,17'd18144,17'd52462,17'd448,17'd796,17'd235,17'd52462,17'd1665,17'd52534,17'd52535,17'd52536,17'd52537,17'd52538,17'd760,17'd52539,17'd52540,17'd27438
},
'{
17'd15877,17'd3101,17'd2258,17'd17,17'd652,17'd1278,17'd286,17'd286,17'd286,17'd286,17'd285,17'd1691,17'd1690,17'd2937,17'd8988,17'd7728,17'd7061,17'd7060,17'd7060,17'd27444,17'd4430,17'd4430,17'd4431,17'd4431,17'd3907,17'd3907,17'd11210,17'd3756,17'd5658,17'd5806,17'd5806,17'd4742,17'd5058,17'd33052,17'd52541,17'd25502,17'd28661,17'd52542,17'd51021,17'd52543,17'd52544,17'd52545,17'd12665,17'd52546,17'd15894,17'd16762,17'd17571,17'd13598,17'd12678,17'd12678,17'd13092,17'd13092,17'd12357,17'd12062,17'd50503,17'd11084,17'd13461,17'd13461,17'd13460,17'd14620,17'd14620,17'd13460,17'd13460,17'd52468,17'd11473,17'd50503,17'd12954,17'd19005,17'd13210,17'd13209,17'd22802,17'd12527,17'd12815,17'd18884,17'd18655,17'd17206,17'd16766,17'd17205,17'd18174,17'd17205,17'd15765,17'd15765,17'd9702,17'd9300,17'd52547,17'd52548,17'd52549,17'd52373,17'd4770,17'd3784,17'd7090,17'd7913,17'd5839,17'd6319,17'd52550,17'd52551,17'd52474,17'd52552,17'd52473,17'd39815,17'd6486,17'd48304,17'd42506,17'd52380,17'd50394,17'd50765,17'd51421,17'd51258,17'd52553,17'd38742,17'd52554,17'd52555,17'd32428,17'd30662,17'd27841,17'd27724,17'd52479,17'd21811,17'd20443,17'd52556,17'd52557,17'd52558,17'd52559,17'd52560,17'd52561,17'd52562,17'd27731,17'd52563,17'd10317,17'd10156,17'd11128,17'd52564,17'd11124,17'd11124,17'd12248,17'd12248,17'd11265,17'd52483,17'd52565,17'd52566,17'd52567,17'd32604,17'd52568,17'd14523,17'd14930,17'd14525,17'd13517,17'd15570,17'd15433,17'd15433,17'd12106,17'd12719,17'd15053,17'd12582,17'd18806,17'd18806,17'd14258,17'd21363,17'd24992,17'd28105,17'd30071,17'd31439,17'd31127,17'd35644,17'd50952,17'd51958,17'd52401,17'd52302,17'd52303,17'd51602,17'd50952,17'd50111,17'd32592,17'd30834,17'd29067,17'd28227,17'd26149,17'd24995,17'd23169,17'd22817,17'd11808,17'd14931,17'd24860,17'd17121,17'd14810,17'd14931,17'd11131,17'd14263,17'd11131,17'd14931,17'd12720,17'd14262,17'd11963,17'd11667,17'd14806,17'd16680,17'd9621,17'd8409,17'd23517,17'd9046,17'd10336,17'd16328,17'd9479,17'd12116,17'd11528,17'd14518,17'd11274,17'd13762,17'd11396,17'd11807,17'd13135,17'd13135,17'd12113,17'd12112,17'd16797,17'd24860,17'd11528,17'd16793,17'd16681,17'd8570,17'd24547,17'd11967,17'd9887,17'd8730,17'd34039,17'd25814,17'd18556,17'd38236,17'd9346,17'd8873,17'd22473,17'd15945,17'd15945,17'd8415,17'd10608,17'd16918,17'd52569,17'd52570,17'd52571,17'd52572,17'd16578,17'd24056,17'd52492,17'd52573,17'd52574,17'd52575,17'd52576,17'd52577,17'd52578,17'd52579,17'd52580,17'd20770,17'd51987,17'd16090,17'd134,17'd130,17'd5593,17'd11821,17'd51730,17'd20921,17'd52581,17'd52582,17'd42441,17'd52583,17'd51307,17'd52584,17'd52585,17'd49977,17'd52586,17'd48707,17'd45150,17'd50072,17'd52000,17'd52000,17'd50272,17'd50574,17'd50574,17'd50268,17'd50371,17'd50160,17'd49684,17'd49681,17'd46657,17'd43289,17'd32506,17'd32017,17'd28257,17'd28256,17'd28487,17'd52429,17'd28256,17'd26780,17'd28725,17'd28602,17'd28599,17'd52587,17'd33163,17'd46836,17'd36542,17'd27027,17'd27372,17'd31353,17'd28371,17'd29690,17'd29978,17'd29979,17'd49790,17'd30280,17'd31506,17'd33489,17'd33323,17'd34117,17'd30131,17'd49790,17'd29690,17'd29690,17'd34114,17'd29833,17'd32508,17'd32508,17'd33167,17'd28858,17'd41863,17'd42593,17'd49480,17'd48155,17'd49289,17'd51390,17'd52588,17'd52589,17'd52512,17'd52511,17'd50907,17'd52590,17'd49388,17'd52591,17'd46201,17'd42884,17'd44229,17'd25435,17'd28484,17'd28254,17'd24902,17'd29828,17'd23038,17'd40052,17'd39742,17'd32667,17'd29099,17'd32186,17'd30431,17'd23918,17'd40833,17'd33479,17'd44825,17'd33648,17'd31658,17'd21846,17'd31346,17'd22170,17'd51563,17'd52592,17'd52593,17'd52594,17'd51084,17'd35294,17'd42150,17'd32011,17'd52440,17'd33946,17'd46002,17'd52595,17'd52596,17'd52597,17'd52598,17'd52599,17'd52600,17'd21760,17'd52601,17'd47467,17'd52521,17'd52602,17'd6844,17'd5916,17'd26709,17'd6553,17'd26451,17'd5607,17'd5477,17'd33041,17'd5754,17'd4997,17'd5152,17'd30180,17'd31891,17'd6390,17'd7499,17'd7668,17'd7499,17'd6219,17'd6390,17'd6554,17'd27935,17'd28185,17'd5160,17'd5160,17'd30638,17'd30638,17'd31891,17'd31717,17'd6554,17'd6390,17'd6390,17'd6219,17'd6219,17'd6219,17'd8304,17'd8304,17'd7499,17'd32073,17'd6554,17'd31717,17'd30638,17'd5004,17'd30638,17'd36887,17'd52182,17'd36311,17'd52603,17'd52604,17'd52605,17'd52606,17'd52450,17'd52273,17'd52607,17'd52608,17'd52609,17'd2528,17'd52610,17'd52611,17'd52612,17'd2546,17'd52613,17'd52614,17'd52019,17'd52276,17'd41000,17'd4056,17'd41159,17'd48559,17'd18383,17'd5026,17'd52020,17'd5497,17'd3898,17'd1824,17'd52615,17'd3426,17'd1825,17'd1824,17'd2558,17'd2558,17'd4059,17'd960,17'd18144,17'd18144,17'd796,17'd796,17'd235,17'd52462,17'd2738,17'd34930,17'd52535,17'd19362,17'd52537,17'd52616,17'd52617,17'd52618,17'd52619,17'd52620
},
'{
17'd15877,17'd2934,17'd52621,17'd1415,17'd652,17'd1278,17'd286,17'd286,17'd286,17'd285,17'd1832,17'd1691,17'd1690,17'd1690,17'd8047,17'd7728,17'd7061,17'd7060,17'd7060,17'd27444,17'd4430,17'd4430,17'd4431,17'd4431,17'd3907,17'd3907,17'd11210,17'd5657,17'd5806,17'd5806,17'd5806,17'd4742,17'd51415,17'd32088,17'd30048,17'd51862,17'd4099,17'd52542,17'd51021,17'd52622,17'd13194,17'd52545,17'd12515,17'd52546,17'd15894,17'd51499,17'd51418,17'd17444,17'd12678,17'd13092,17'd13092,17'd13092,17'd12357,17'd12062,17'd11084,17'd11084,17'd50503,17'd50503,17'd13460,17'd14620,17'd14620,17'd13460,17'd13460,17'd14620,17'd11473,17'd50503,17'd12954,17'd13210,17'd13463,17'd13598,17'd14469,17'd22802,17'd23154,17'd12531,17'd18774,17'd19007,17'd16766,17'd17205,17'd19891,17'd17205,17'd10943,17'd10944,17'd15517,17'd13845,17'd14100,17'd52548,17'd52623,17'd52624,17'd52625,17'd3784,17'd3949,17'd7913,17'd5839,17'd7257,17'd52626,17'd51868,17'd52627,17'd52628,17'd52286,17'd39057,17'd39505,17'd49716,17'd42506,17'd52629,17'd52630,17'd50847,17'd50765,17'd51257,17'd50766,17'd52631,17'd52632,17'd52633,17'd52634,17'd52119,17'd9025,17'd27842,17'd27469,17'd52635,17'd52636,17'd52637,17'd10303,17'd52039,17'd52638,17'd52214,17'd52639,17'd52640,17'd52641,17'd52642,17'd27617,17'd10970,17'd10156,17'd11269,17'd28100,17'd11954,17'd12248,17'd12248,17'd17228,17'd52643,17'd52644,17'd52645,17'd52646,17'd52647,17'd33098,17'd30231,17'd14930,17'd14930,17'd14525,17'd21207,17'd15433,17'd15433,17'd15685,17'd15685,17'd11958,17'd12581,17'd12582,17'd18806,17'd20609,17'd20450,17'd21505,17'd24538,17'd28943,17'd30072,17'd30973,17'd31943,17'd50863,17'd51512,17'd52401,17'd52401,17'd52648,17'd52402,17'd51881,17'd50951,17'd31590,17'd33568,17'd31440,17'd28461,17'd26873,17'd28231,17'd21362,17'd18681,17'd13645,17'd10853,17'd10604,17'd24860,17'd12720,17'd14810,17'd10990,17'd11131,17'd14263,17'd10854,17'd24860,17'd11519,17'd13362,17'd13253,17'd24034,17'd52649,17'd10174,17'd15178,17'd30672,17'd22473,17'd29920,17'd17480,17'd16328,17'd10742,17'd17839,17'd10606,17'd10990,17'd16068,17'd11807,17'd11667,17'd13135,17'd12858,17'd12259,17'd15809,17'd21204,17'd18805,17'd51273,17'd9883,17'd20757,17'd52650,17'd24368,17'd8576,17'd25148,17'd13257,17'd52651,17'd28237,17'd18556,17'd9884,17'd10992,17'd9347,17'd12722,17'd37334,17'd25679,17'd8418,17'd18686,17'd12120,17'd14390,17'd52225,17'd52652,17'd52653,17'd15069,17'd52654,17'd52655,17'd52656,17'd52657,17'd52658,17'd52659,17'd52660,17'd52661,17'd52662,17'd52663,17'd51987,17'd11683,17'd131,17'd3025,17'd133,17'd131,17'd52664,17'd52665,17'd52666,17'd52667,17'd52160,17'd31030,17'd52668,17'd49976,17'd52669,17'd52670,17'd46662,17'd47535,17'd48049,17'd49988,17'd52000,17'd52671,17'd51741,17'd50272,17'd50072,17'd50736,17'd51157,17'd50160,17'd49787,17'd40952,17'd39580,17'd44476,17'd32004,17'd28370,17'd29380,17'd28256,17'd52672,17'd40050,17'd49179,17'd30279,17'd28726,17'd27883,17'd40828,17'd48043,17'd33815,17'd35854,17'd31503,17'd26901,17'd26902,17'd26055,17'd49086,17'd29831,17'd49790,17'd29979,17'd29979,17'd30131,17'd30280,17'd30736,17'd30280,17'd49790,17'd49790,17'd29979,17'd29690,17'd29536,17'd29536,17'd34114,17'd34114,17'd32508,17'd32508,17'd32508,17'd50369,17'd47333,17'd48041,17'd48259,17'd49082,17'd49390,17'd51995,17'd52673,17'd52674,17'd52589,17'd52675,17'd50163,17'd52676,17'd47536,17'd52677,17'd52678,17'd45036,17'd42749,17'd42749,17'd28850,17'd24742,17'd23566,17'd23389,17'd22857,17'd51747,17'd33949,17'd29828,17'd23920,17'd30431,17'd29534,17'd23918,17'd32015,17'd40679,17'd40369,17'd31346,17'd31830,17'd21846,17'd31660,17'd51302,17'd52174,17'd52679,17'd52680,17'd52681,17'd51226,17'd34280,17'd42150,17'd47948,17'd52515,17'd52682,17'd35155,17'd52683,17'd47155,17'd52087,17'd52684,17'd52685,17'd20502,17'd21919,17'd50584,17'd27080,17'd10627,17'd52686,17'd6844,17'd5916,17'd6218,17'd6707,17'd5758,17'd5322,17'd4521,17'd4521,17'd5754,17'd5144,17'd5327,17'd30637,17'd31717,17'd9091,17'd7499,17'd7668,17'd7668,17'd9091,17'd6390,17'd6390,17'd27935,17'd27935,17'd28185,17'd28185,17'd28185,17'd28185,17'd31717,17'd6554,17'd32073,17'd9091,17'd9091,17'd9091,17'd9091,17'd9091,17'd6220,17'd6220,17'd7499,17'd9091,17'd6554,17'd28185,17'd5160,17'd5004,17'd36887,17'd36887,17'd35760,17'd52687,17'd36032,17'd52688,17'd52689,17'd49104,17'd52690,17'd52451,17'd52691,17'd52692,17'd52693,17'd52694,17'd52695,17'd23127,17'd52018,17'd52696,17'd51938,17'd52193,17'd50182,17'd50001,17'd52697,17'd40411,17'd41159,17'd48559,17'd18383,17'd5026,17'd4557,17'd11049,17'd1824,17'd1825,17'd52615,17'd3426,17'd1402,17'd3072,17'd2558,17'd4398,17'd52698,17'd1265,17'd18144,17'd52363,17'd448,17'd796,17'd1943,17'd52462,17'd36181,17'd20710,17'd763,17'd52699,17'd52616,17'd52367,17'd52700,17'd52701,17'd52702,17'd52703
},
'{
17'd52704,17'd3901,17'd10669,17'd1415,17'd652,17'd1278,17'd286,17'd286,17'd286,17'd286,17'd285,17'd1691,17'd1690,17'd2937,17'd8988,17'd7728,17'd7061,17'd7060,17'd7060,17'd27444,17'd4430,17'd4430,17'd4431,17'd4431,17'd3907,17'd3907,17'd11210,17'd3756,17'd5658,17'd5806,17'd5806,17'd4742,17'd51415,17'd33052,17'd52541,17'd29176,17'd3924,17'd52542,17'd51021,17'd52705,17'd52706,17'd24338,17'd52707,17'd12942,17'd19749,17'd52708,17'd52709,17'd32896,17'd12678,17'd13092,17'd13092,17'd13092,17'd12357,17'd12062,17'd50503,17'd50503,17'd11084,17'd50503,17'd13460,17'd14620,17'd14620,17'd13460,17'd13460,17'd14620,17'd11473,17'd50503,17'd12954,17'd13599,17'd13463,17'd13462,17'd14468,17'd22802,17'd23154,17'd20424,17'd17689,17'd19007,17'd19754,17'd17205,17'd18174,17'd17205,17'd11088,17'd10944,17'd10429,17'd13845,17'd14099,17'd47866,17'd52710,17'd52471,17'd52625,17'd3629,17'd3628,17'd3626,17'd5839,17'd6472,17'd43887,17'd52550,17'd52627,17'd52474,17'd52285,17'd39814,17'd40426,17'd50095,17'd52711,17'd52629,17'd52630,17'd51104,17'd50765,17'd51257,17'd50766,17'd52712,17'd52713,17'd52714,17'd50197,17'd8393,17'd28443,17'd27607,17'd27468,17'd52715,17'd52636,17'd10137,17'd52480,17'd17222,17'd10447,17'd52716,17'd51508,17'd15037,17'd52717,17'd52718,17'd27476,17'd28095,17'd10970,17'd10465,17'd52719,17'd24853,17'd12248,17'd17228,17'd52720,17'd52721,17'd52722,17'd52723,17'd52724,17'd20172,17'd52725,17'd29205,17'd14523,17'd14930,17'd14930,17'd21057,17'd15570,17'd15433,17'd15685,17'd13252,17'd11958,17'd12719,17'd18917,17'd12582,17'd20609,17'd20609,17'd20608,17'd23170,17'd29778,17'd29329,17'd31765,17'd32920,17'd50863,17'd51692,17'd52401,17'd52401,17'd52648,17'd52648,17'd51959,17'd51958,17'd35239,17'd34037,17'd31941,17'd29330,17'd28573,17'd31443,17'd24705,17'd14258,17'd19643,17'd11129,17'd10990,17'd14931,17'd12720,17'd12720,17'd14810,17'd10854,17'd14263,17'd14263,17'd16320,17'd12720,17'd11667,17'd15185,17'd11521,17'd52726,17'd15048,17'd16794,17'd32921,17'd8573,17'd33404,17'd39660,17'd10173,17'd10742,17'd17839,17'd17720,17'd10476,17'd14673,17'd13253,17'd13253,17'd11806,17'd12858,17'd11958,17'd13365,17'd13763,17'd12718,17'd11667,17'd12862,17'd11276,17'd52727,17'd10338,17'd24546,17'd50523,17'd13257,17'd52728,17'd38904,17'd14674,17'd15048,17'd9741,17'd9339,17'd8567,17'd44981,17'd9196,17'd10028,17'd18686,17'd14676,17'd10180,17'd12591,17'd17133,17'd52729,17'd52730,17'd52731,17'd52732,17'd52733,17'd52734,17'd52735,17'd52736,17'd52737,17'd52409,17'd52738,17'd20623,17'd20465,17'd52245,17'd131,17'd11413,17'd1045,17'd5593,17'd20768,17'd52739,17'd52740,17'd52741,17'd35293,17'd40521,17'd51735,17'd52742,17'd52743,17'd50566,17'd48443,17'd49889,17'd48909,17'd50365,17'd51652,17'd52671,17'd50371,17'd50476,17'd50736,17'd50268,17'd50160,17'd49788,17'd49382,17'd52340,17'd46657,17'd43560,17'd32356,17'd29380,17'd29106,17'd28256,17'd49179,17'd28487,17'd28256,17'd33952,17'd46431,17'd52744,17'd52745,17'd35578,17'd32016,17'd39743,17'd38537,17'd34767,17'd33963,17'd25696,17'd49284,17'd29979,17'd33489,17'd49579,17'd29979,17'd30280,17'd30280,17'd30280,17'd30131,17'd49790,17'd49790,17'd29690,17'd29690,17'd28857,17'd29536,17'd34285,17'd34114,17'd32508,17'd34285,17'd36989,17'd37248,17'd52746,17'd39580,17'd48616,17'd47641,17'd49485,17'd52747,17'd52748,17'd52674,17'd52749,17'd50371,17'd50822,17'd52750,17'd47340,17'd52751,17'd42742,17'd37778,17'd42749,17'd29825,17'd25179,17'd29100,17'd29374,17'd22679,17'd36009,17'd52752,17'd32830,17'd23566,17'd24249,17'd32659,17'd29534,17'd29376,17'd45754,17'd50826,17'd38041,17'd31658,17'd23220,17'd49488,17'd22864,17'd42440,17'd52753,17'd21387,17'd52754,17'd51654,17'd35293,17'd51912,17'd34280,17'd41728,17'd52515,17'd41728,17'd52755,17'd52756,17'd52757,17'd52758,17'd52759,17'd52760,17'd20220,17'd24138,17'd25482,17'd26826,17'd10359,17'd52686,17'd6844,17'd5916,17'd6218,17'd6706,17'd5326,17'd52761,17'd33041,17'd4521,17'd5754,17'd5153,17'd28536,17'd31553,17'd6554,17'd9091,17'd7499,17'd7668,17'd27696,17'd29740,17'd32073,17'd6390,17'd27935,17'd27935,17'd28185,17'd28185,17'd28185,17'd31717,17'd6554,17'd6554,17'd32073,17'd9091,17'd9091,17'd9091,17'd9091,17'd7499,17'd6220,17'd6220,17'd7499,17'd9091,17'd6554,17'd28185,17'd25627,17'd5004,17'd36887,17'd37434,17'd35760,17'd52762,17'd52763,17'd38322,17'd52764,17'd52765,17'd52766,17'd52451,17'd52767,17'd35902,17'd52768,17'd52769,17'd52695,17'd52770,17'd52771,17'd37571,17'd51938,17'd50384,17'd52772,17'd51412,17'd9530,17'd43742,17'd41159,17'd48559,17'd18383,17'd5026,17'd4557,17'd11049,17'd1825,17'd52615,17'd52615,17'd3426,17'd3072,17'd3072,17'd2558,17'd4398,17'd52698,17'd960,17'd1943,17'd1943,17'd796,17'd796,17'd1943,17'd8164,17'd36322,17'd52773,17'd18983,17'd26122,17'd51859,17'd52774,17'd25782,17'd52775,17'd52776,17'd52777
},
'{
17'd52778,17'd3592,17'd10802,17'd2596,17'd289,17'd653,17'd287,17'd28,17'd286,17'd285,17'd1832,17'd1691,17'd1690,17'd1690,17'd8047,17'd7728,17'd7061,17'd7061,17'd7060,17'd7060,17'd4430,17'd4430,17'd4431,17'd4431,17'd3907,17'd3907,17'd11210,17'd5657,17'd5806,17'd5806,17'd5806,17'd4742,17'd51415,17'd32088,17'd30048,17'd51862,17'd28433,17'd6447,17'd52779,17'd52705,17'd52706,17'd13195,17'd12344,17'd12800,17'd52780,17'd18406,17'd16162,17'd32896,17'd12678,17'd12678,17'd14469,17'd14469,17'd12357,17'd12357,17'd12062,17'd12062,17'd11084,17'd50503,17'd13461,17'd12355,17'd14620,17'd13460,17'd13460,17'd14620,17'd11473,17'd50503,17'd13092,17'd13599,17'd13463,17'd13462,17'd14468,17'd14469,17'd17096,17'd20885,17'd19382,17'd18774,17'd19754,17'd16766,17'd18174,17'd17205,17'd10943,17'd10944,17'd10429,17'd15898,17'd15009,17'd15384,17'd48387,17'd52781,17'd52782,17'd52783,17'd3948,17'd3626,17'd3470,17'd6631,17'd43470,17'd52784,17'd52474,17'd52785,17'd52286,17'd39504,17'd39816,17'd48304,17'd42505,17'd42666,17'd52630,17'd51022,17'd41333,17'd50934,17'd50935,17'd52786,17'd52787,17'd52632,17'd50297,17'd52788,17'd29909,17'd27607,17'd27724,17'd26860,17'd22123,17'd52385,17'd52556,17'd18072,17'd16424,17'd10582,17'd26618,17'd26361,17'd15416,17'd26489,17'd52789,17'd27476,17'd52790,17'd52791,17'd26867,17'd26031,17'd27341,17'd15293,17'd11392,17'd52792,17'd52793,17'd13756,17'd52794,17'd52795,17'd18914,17'd52796,17'd14523,17'd14930,17'd14930,17'd14525,17'd52797,17'd51039,17'd15685,17'd13252,17'd11958,17'd12719,17'd12996,17'd16204,17'd18681,17'd19921,17'd25143,17'd25926,17'd24537,17'd28943,17'd31440,17'd31127,17'd51118,17'd52798,17'd51692,17'd51881,17'd52402,17'd52799,17'd52800,17'd52132,17'd50952,17'd35644,17'd31287,17'd30676,17'd29924,17'd28227,17'd24857,17'd26035,17'd18681,17'd14671,17'd11275,17'd10990,17'd14810,17'd12720,17'd14673,17'd11808,17'd14263,17'd14263,17'd10739,17'd14810,17'd14133,17'd19158,17'd15185,17'd16069,17'd45549,17'd18324,17'd52801,17'd12866,17'd24711,17'd33404,17'd15944,17'd10742,17'd11134,17'd11133,17'd14518,17'd17236,17'd16069,17'd11667,17'd12861,17'd12113,17'd11958,17'd12419,17'd12419,17'd12110,17'd12857,17'd13253,17'd13001,17'd11277,17'd9042,17'd30969,17'd9887,17'd23173,17'd52802,17'd47292,17'd29920,17'd50609,17'd16549,17'd9480,17'd16067,17'd8731,17'd52803,17'd9887,17'd10028,17'd12120,17'd11534,17'd25155,17'd16920,17'd52804,17'd52805,17'd52806,17'd52807,17'd52808,17'd52809,17'd52311,17'd52810,17'd52811,17'd21067,17'd15823,17'd131,17'd11541,17'd131,17'd131,17'd1045,17'd133,17'd20623,17'd52812,17'd52813,17'd52814,17'd51563,17'd31660,17'd52815,17'd52816,17'd46548,17'd52817,17'd52818,17'd52255,17'd44929,17'd49582,17'd51830,17'd52001,17'd51741,17'd50476,17'd50476,17'd50272,17'd50268,17'd51390,17'd50467,17'd48446,17'd43150,17'd44698,17'd34104,17'd33485,17'd28372,17'd31196,17'd28372,17'd28487,17'd28371,17'd28854,17'd37513,17'd46431,17'd52819,17'd35023,17'd31503,17'd39910,17'd31503,17'd38537,17'd28979,17'd44703,17'd27768,17'd49578,17'd29979,17'd30280,17'd32508,17'd29981,17'd30130,17'd30130,17'd49790,17'd49579,17'd29690,17'd29690,17'd29536,17'd28857,17'd28857,17'd28857,17'd29690,17'd29690,17'd32833,17'd36989,17'd38154,17'd43547,17'd49282,17'd43148,17'd46847,17'd47737,17'd49692,17'd52820,17'd52748,17'd52821,17'd52001,17'd50365,17'd49091,17'd52822,17'd48254,17'd52823,17'd44230,17'd32996,17'd43977,17'd38406,17'd28977,17'd23564,17'd23216,17'd34458,17'd30427,17'd52824,17'd37117,17'd23918,17'd23916,17'd35159,17'd30424,17'd29829,17'd35158,17'd50826,17'd48911,17'd33312,17'd32829,17'd49488,17'd34617,17'd51921,17'd52825,17'd21538,17'd52594,17'd52345,17'd34880,17'd34617,17'd33946,17'd35710,17'd35155,17'd42441,17'd46574,17'd52826,17'd52827,17'd52828,17'd52829,17'd52830,17'd21130,17'd52831,17'd11985,17'd26448,17'd52832,17'd7165,17'd6382,17'd5916,17'd6388,17'd24800,17'd5325,17'd33365,17'd43584,17'd4520,17'd4188,17'd42910,17'd4842,17'd30333,17'd6554,17'd6219,17'd7499,17'd7668,17'd29740,17'd32074,17'd36586,17'd6554,17'd6554,17'd31717,17'd28185,17'd28185,17'd31717,17'd6554,17'd6554,17'd32073,17'd9091,17'd9091,17'd9091,17'd9091,17'd7499,17'd7499,17'd6220,17'd6220,17'd6220,17'd6219,17'd27935,17'd30638,17'd25627,17'd25627,17'd37030,17'd5338,17'd34336,17'd52833,17'd52834,17'd52835,17'd52836,17'd52525,17'd52273,17'd52014,17'd52837,17'd52838,17'd2214,17'd52839,17'd36320,17'd52840,17'd52841,17'd37571,17'd3061,17'd52460,17'd50290,17'd50001,17'd4054,17'd40411,17'd41159,17'd48559,17'd18383,17'd5026,17'd4557,17'd5497,17'd1825,17'd52615,17'd52615,17'd1825,17'd2558,17'd2558,17'd4398,17'd38071,17'd796,17'd960,17'd1943,17'd1943,17'd628,17'd628,17'd1943,17'd8164,17'd36322,17'd52773,17'd18983,17'd34164,17'd52842,17'd52198,17'd25494,17'd52843,17'd52844,17'd52845
},
'{
17'd52778,17'd5204,17'd3251,17'd2596,17'd289,17'd653,17'd28,17'd28,17'd286,17'd286,17'd285,17'd1691,17'd1690,17'd2937,17'd8988,17'd7728,17'd7061,17'd7061,17'd7060,17'd7060,17'd4430,17'd4430,17'd4431,17'd4431,17'd3907,17'd3907,17'd11210,17'd3756,17'd5210,17'd5806,17'd5806,17'd4742,17'd51415,17'd33052,17'd52541,17'd29176,17'd4902,17'd27323,17'd52779,17'd52846,17'd52706,17'd13195,17'd12514,17'd12800,17'd52847,17'd18406,17'd18057,17'd52848,17'd16407,17'd12678,17'd14469,17'd14469,17'd12357,17'd12357,17'd12357,17'd12357,17'd11084,17'd50503,17'd13461,17'd12355,17'd14620,17'd14620,17'd14620,17'd14620,17'd11473,17'd50503,17'd13092,17'd13599,17'd13463,17'd13462,17'd14468,17'd22802,17'd23154,17'd20424,17'd17204,17'd17689,17'd19754,17'd19754,17'd17205,17'd17205,17'd10943,17'd10944,17'd10429,17'd13972,17'd52849,17'd47971,17'd52850,17'd52851,17'd3632,17'd4612,17'd3948,17'd3626,17'd3470,17'd6309,17'd52852,17'd6320,17'd52853,17'd52552,17'd52473,17'd39814,17'd40583,17'd40584,17'd48564,17'd42666,17'd6648,17'd51022,17'd41333,17'd50934,17'd50935,17'd52854,17'd49415,17'd50507,17'd35362,17'd8553,17'd52855,17'd52856,17'd27332,17'd52479,17'd26027,17'd20895,17'd52212,17'd52038,17'd18433,17'd16786,17'd52481,17'd52857,17'd26619,17'd52858,17'd52859,17'd52860,17'd52861,17'd27230,17'd52862,17'd26867,17'd24989,17'd26751,17'd52792,17'd52863,17'd26364,17'd52864,17'd52865,17'd52866,17'd52646,17'd52725,17'd29205,17'd14672,17'd14672,17'd14930,17'd21057,17'd52797,17'd15570,17'd13252,17'd11958,17'd12719,17'd12996,17'd12996,17'd18443,17'd18681,17'd25143,17'd33084,17'd24705,17'd29778,17'd28686,17'd31941,17'd32920,17'd51272,17'd52867,17'd51959,17'd52868,17'd52869,17'd52870,17'd52871,17'd51881,17'd50863,17'd32920,17'd31941,17'd37065,17'd30071,17'd29327,17'd24031,17'd22472,17'd18444,17'd19533,17'd11808,17'd11274,17'd14673,17'd14673,17'd11274,17'd11275,17'd11131,17'd10739,17'd14931,17'd11396,17'd14379,17'd11961,17'd11963,17'd52872,17'd18196,17'd52873,17'd52874,17'd12119,17'd52803,17'd17123,17'd10743,17'd17719,17'd11133,17'd11527,17'd10476,17'd11274,17'd13762,17'd11962,17'd12861,17'd11961,17'd12419,17'd12110,17'd12109,17'd12580,17'd11961,17'd11666,17'd31130,17'd11809,17'd29333,17'd30523,17'd9887,17'd13257,17'd11967,17'd8413,17'd8723,17'd17716,17'd51696,17'd16071,17'd8724,17'd26154,17'd52222,17'd19923,17'd17850,17'd15441,17'd52875,17'd15573,17'd52876,17'd52877,17'd52878,17'd52879,17'd52880,17'd52881,17'd52882,17'd52883,17'd52884,17'd15823,17'd133,17'd128,17'd132,17'd131,17'd11541,17'd133,17'd15823,17'd20625,17'd52578,17'd52885,17'd52886,17'd35293,17'd34279,17'd52887,17'd52888,17'd46548,17'd48037,17'd46757,17'd52256,17'd52590,17'd50574,17'd52671,17'd51741,17'd50272,17'd50907,17'd50476,17'd51830,17'd50268,17'd49683,17'd48904,17'd43542,17'd45264,17'd46094,17'd36127,17'd32355,17'd30587,17'd52889,17'd29106,17'd28857,17'd29380,17'd28854,17'd33952,17'd44703,17'd34767,17'd31354,17'd38026,17'd37250,17'd29245,17'd28727,17'd29246,17'd44826,17'd51918,17'd50906,17'd29979,17'd49790,17'd29981,17'd31037,17'd30130,17'd29979,17'd49579,17'd49579,17'd29690,17'd29690,17'd28857,17'd28857,17'd28857,17'd28857,17'd29690,17'd29690,17'd32833,17'd36989,17'd48042,17'd51651,17'd52890,17'd46666,17'd47054,17'd48909,17'd50164,17'd52891,17'd52674,17'd52892,17'd51830,17'd49582,17'd51557,17'd47934,17'd52893,17'd52894,17'd43978,17'd33643,17'd43977,17'd38667,17'd34467,17'd23386,17'd30425,17'd22857,17'd31343,17'd31656,17'd23923,17'd30879,17'd28851,17'd30126,17'd33801,17'd23388,17'd34638,17'd31499,17'd23393,17'd39745,17'd49094,17'd49488,17'd51302,17'd52895,17'd52896,17'd52680,17'd51382,17'd46455,17'd51302,17'd42150,17'd35710,17'd41275,17'd35710,17'd52897,17'd46765,17'd46963,17'd52898,17'd52899,17'd52900,17'd52901,17'd52902,17'd52903,17'd52904,17'd52905,17'd9907,17'd6212,17'd5914,17'd5916,17'd26451,17'd5482,17'd24798,17'd52906,17'd33041,17'd4522,17'd4838,17'd4995,17'd30637,17'd30638,17'd6390,17'd6219,17'd7499,17'd27696,17'd35052,17'd32074,17'd37152,17'd6554,17'd6554,17'd31717,17'd28185,17'd30638,17'd31717,17'd6554,17'd36586,17'd32073,17'd9091,17'd7499,17'd7499,17'd7499,17'd7499,17'd7499,17'd6220,17'd6220,17'd6219,17'd6390,17'd28185,17'd30333,17'd25627,17'd5160,17'd37030,17'd5338,17'd34336,17'd37698,17'd52907,17'd52908,17'd52909,17'd52525,17'd51847,17'd52910,17'd52911,17'd23124,17'd52912,17'd52913,17'd23298,17'd52914,17'd52915,17'd37571,17'd3061,17'd52916,17'd52917,17'd51855,17'd6081,17'd40411,17'd41159,17'd48559,17'd10906,17'd5026,17'd52020,17'd52918,17'd3426,17'd52615,17'd52615,17'd1825,17'd2391,17'd2558,17'd4398,17'd38071,17'd796,17'd1121,17'd18144,17'd235,17'd447,17'd447,17'd1121,17'd8164,17'd36322,17'd52919,17'd52920,17'd52921,17'd52922,17'd52923,17'd52924,17'd52925,17'd52926,17'd52927
},
'{
17'd52928,17'd5204,17'd3251,17'd2596,17'd809,17'd289,17'd287,17'd28,17'd286,17'd285,17'd1832,17'd1691,17'd52025,17'd8047,17'd8988,17'd9275,17'd7061,17'd7061,17'd7060,17'd7060,17'd4430,17'd4430,17'd4431,17'd4431,17'd3907,17'd3907,17'd11210,17'd5379,17'd5055,17'd5806,17'd5806,17'd4742,17'd51861,17'd4437,17'd52541,17'd29176,17'd4902,17'd4100,17'd52779,17'd52929,17'd52930,17'd13312,17'd12514,17'd12800,17'd52847,17'd52931,17'd18057,17'd52848,17'd15762,17'd13597,17'd14469,17'd14469,17'd12357,17'd12357,17'd12062,17'd12357,17'd50503,17'd14763,17'd50503,17'd11084,17'd14620,17'd14620,17'd14620,17'd14620,17'd11473,17'd50503,17'd13598,17'd13463,17'd13968,17'd13462,17'd14468,17'd14469,17'd17096,17'd30058,17'd19006,17'd17689,17'd19754,17'd19754,17'd17205,17'd18174,17'd16766,17'd10943,17'd10429,17'd15766,17'd15009,17'd15641,17'd33857,17'd52932,17'd52933,17'd4612,17'd3948,17'd3781,17'd3469,17'd5842,17'd52934,17'd6311,17'd46367,17'd50006,17'd52113,17'd39504,17'd40582,17'd40427,17'd42063,17'd42666,17'd6648,17'd52630,17'd51104,17'd50934,17'd52935,17'd52936,17'd49415,17'd52631,17'd50681,17'd52937,17'd52938,17'd27723,17'd51782,17'd23158,17'd52939,17'd24527,17'd52940,17'd52941,17'd20896,17'd52942,17'd52559,17'd26618,17'd15038,17'd52943,17'd52944,17'd52945,17'd52946,17'd52947,17'd52862,17'd26257,17'd11952,17'd11392,17'd52948,17'd52949,17'd26366,17'd24986,17'd52950,17'd52643,17'd52484,17'd52647,17'd29205,17'd13642,17'd14672,17'd14672,17'd14525,17'd21057,17'd15942,17'd21506,17'd13136,17'd11958,17'd13135,17'd12996,17'd16442,17'd18681,17'd44982,17'd20450,17'd28459,17'd27347,17'd30831,17'd39211,17'd32592,17'd52951,17'd52867,17'd52867,17'd52401,17'd52869,17'd52870,17'd52870,17'd51959,17'd51512,17'd35093,17'd31127,17'd32761,17'd30832,17'd29328,17'd25927,17'd24362,17'd18443,17'd24029,17'd11275,17'd11274,17'd11274,17'd14673,17'd14673,17'd11274,17'd10854,17'd10475,17'd10854,17'd18326,17'd23171,17'd13363,17'd11957,17'd29477,17'd16908,17'd9041,17'd33570,17'd33405,17'd9196,17'd24999,17'd23679,17'd23339,17'd19532,17'd20756,17'd10991,17'd11965,17'd12262,17'd11666,17'd13764,17'd13764,17'd13363,17'd13882,17'd18450,17'd12580,17'd12580,17'd11961,17'd12862,17'd15943,17'd18080,17'd12118,17'd52952,17'd17126,17'd8418,17'd52953,17'd12865,17'd9046,17'd34039,17'd23860,17'd17607,17'd32924,17'd33879,17'd11967,17'd13375,17'd22133,17'd23175,17'd52954,17'd52955,17'd52956,17'd52957,17'd52958,17'd52959,17'd20058,17'd52960,17'd52961,17'd20464,17'd7980,17'd133,17'd128,17'd129,17'd135,17'd132,17'd1481,17'd13777,17'd23360,17'd52962,17'd52963,17'd52964,17'd22012,17'd52965,17'd52966,17'd52967,17'd52968,17'd52969,17'd52970,17'd52971,17'd52972,17'd51744,17'd52973,17'd52974,17'd50476,17'd50907,17'd50272,17'd51830,17'd50072,17'd49485,17'd49279,17'd52975,17'd44933,17'd34105,17'd27885,17'd32355,17'd29104,17'd28856,17'd30884,17'd30884,17'd32193,17'd28134,17'd29977,17'd37513,17'd32356,17'd52976,17'd29981,17'd33321,17'd31035,17'd34637,17'd27642,17'd32192,17'd29537,17'd31038,17'd29690,17'd29690,17'd31037,17'd30434,17'd29981,17'd32833,17'd29691,17'd30884,17'd29690,17'd29690,17'd28857,17'd28857,17'd28857,17'd28857,17'd29690,17'd29690,17'd49579,17'd52429,17'd39584,17'd52977,17'd52978,17'd46666,17'd48709,17'd48263,17'd51157,17'd52979,17'd52821,17'd52675,17'd50268,17'd49288,17'd52822,17'd52980,17'd52981,17'd52982,17'd32996,17'd28721,17'd39591,17'd32007,17'd23732,17'd29374,17'd30129,17'd39911,17'd31343,17'd39131,17'd29099,17'd24415,17'd25032,17'd30126,17'd29528,17'd23215,17'd33479,17'd36427,17'd23926,17'd46958,17'd48911,17'd41726,17'd35293,17'd52983,17'd52984,17'd52680,17'd51922,17'd52985,17'd34881,17'd22511,17'd42441,17'd34880,17'd48366,17'd52986,17'd52987,17'd52988,17'd52989,17'd52990,17'd52991,17'd21738,17'd21447,17'd52992,17'd52993,17'd52994,17'd7007,17'd6382,17'd5914,17'd5916,17'd5760,17'd5478,17'd52995,17'd52906,17'd4521,17'd4523,17'd5145,17'd4841,17'd5004,17'd28185,17'd5615,17'd6220,17'd7499,17'd27696,17'd35052,17'd52996,17'd37152,17'd6554,17'd6554,17'd6554,17'd28185,17'd28185,17'd6554,17'd6390,17'd32073,17'd32073,17'd32074,17'd29740,17'd29740,17'd29740,17'd7499,17'd7499,17'd6220,17'd6220,17'd6219,17'd6390,17'd28185,17'd30333,17'd25627,17'd5160,17'd36887,17'd5616,17'd34336,17'd37436,17'd52997,17'd52998,17'd52999,17'd53000,17'd53001,17'd52187,17'd47378,17'd53002,17'd53003,17'd36452,17'd36042,17'd2380,17'd53004,17'd37571,17'd3061,17'd52460,17'd53005,17'd40861,17'd53006,17'd4056,17'd48812,17'd5354,17'd18142,17'd52020,17'd52918,17'd4399,17'd3426,17'd52615,17'd3426,17'd1824,17'd2391,17'd2558,17'd38071,17'd4059,17'd628,17'd796,17'd630,17'd235,17'd959,17'd447,17'd1121,17'd3071,17'd36322,17'd53007,17'd19100,17'd52921,17'd53008,17'd53009,17'd52619,17'd53010,17'd53011,17'd53012
},
'{
17'd52928,17'd3902,17'd2934,17'd2596,17'd17187,17'd289,17'd287,17'd287,17'd286,17'd285,17'd285,17'd1691,17'd52025,17'd8047,17'd8988,17'd7728,17'd7061,17'd7061,17'd7060,17'd7060,17'd6744,17'd4430,17'd4431,17'd3907,17'd3907,17'd9816,17'd3756,17'd3434,17'd5210,17'd5806,17'd5806,17'd4742,17'd4897,17'd53013,17'd52541,17'd29176,17'd28661,17'd53014,17'd4440,17'd53015,17'd53016,17'd13444,17'd53017,17'd12516,17'd15128,17'd18772,17'd18295,17'd19125,17'd15762,17'd14469,17'd14469,17'd14469,17'd12357,17'd12062,17'd12062,17'd12062,17'd50503,17'd14763,17'd50503,17'd11084,17'd14620,17'd14620,17'd14620,17'd14620,17'd11473,17'd50503,17'd13598,17'd13463,17'd13463,17'd16284,17'd14468,17'd22802,17'd13093,17'd12815,17'd18884,17'd17689,17'd19893,17'd19754,17'd18174,17'd18174,17'd16766,17'd19754,17'd11231,17'd13470,17'd14099,17'd47973,17'd49200,17'd49200,17'd53018,17'd53019,17'd4289,17'd3781,17'd3469,17'd6007,17'd6310,17'd53020,17'd45667,17'd47094,17'd53021,17'd51868,17'd41498,17'd53022,17'd49016,17'd42937,17'd6648,17'd51022,17'd51104,17'd50296,17'd45198,17'd42065,17'd50680,17'd50598,17'd53023,17'd53024,17'd52788,17'd28672,17'd50401,17'd23158,17'd20598,17'd53025,17'd17112,17'd52212,17'd10303,17'd53026,17'd16541,17'd16900,17'd25668,17'd10714,17'd26489,17'd53027,17'd26621,17'd52947,17'd52861,17'd53028,17'd27479,17'd11514,17'd53029,17'd26364,17'd11659,17'd22470,17'd19915,17'd53030,17'd52644,17'd53031,17'd13641,17'd44647,17'd16686,17'd15571,17'd15687,17'd14525,17'd14526,17'd21506,17'd12995,17'd13519,17'd12719,17'd15053,17'd18917,17'd18443,17'd23169,17'd20609,17'd20608,17'd23682,17'd30218,17'd30527,17'd32283,17'd35093,17'd52867,17'd52133,17'd52301,17'd52869,17'd53032,17'd53032,17'd52800,17'd51692,17'd34828,17'd31442,17'd31287,17'd32761,17'd29924,17'd28227,17'd24538,17'd22472,17'd22817,17'd19533,17'd11808,17'd11808,17'd11274,17'd16068,17'd16068,17'd11808,17'd11131,17'd11131,17'd25280,17'd14133,17'd13135,17'd12857,17'd12112,17'd51273,17'd29090,17'd30969,17'd53033,17'd19923,17'd9046,17'd9481,17'd20755,17'd10329,17'd20756,17'd10606,17'd14931,17'd11395,17'd11666,17'd13885,17'd15175,17'd15299,17'd13882,17'd18450,17'd12579,17'd12580,17'd11960,17'd13253,17'd52872,17'd25676,17'd9337,17'd53034,17'd8098,17'd9484,17'd53035,17'd8249,17'd21987,17'd53036,17'd50522,17'd28353,17'd22645,17'd9042,17'd9744,17'd8579,17'd17127,17'd53037,17'd53038,17'd53039,17'd53040,17'd53041,17'd23006,17'd15068,17'd10873,17'd16220,17'd14017,17'd16090,17'd17363,17'd133,17'd130,17'd130,17'd132,17'd132,17'd128,17'd20622,17'd21835,17'd51458,17'd53042,17'd51066,17'd23742,17'd51074,17'd50362,17'd52743,17'd53043,17'd53044,17'd40517,17'd53045,17'd50907,17'd51920,17'd52973,17'd52974,17'd50736,17'd50907,17'd52000,17'd51830,17'd49890,17'd48264,17'd46667,17'd45621,17'd39585,17'd35570,17'd28134,17'd32355,17'd29247,17'd30587,17'd30884,17'd29691,17'd36988,17'd32507,17'd33164,17'd33319,17'd52976,17'd53046,17'd32833,17'd53047,17'd28980,17'd31352,17'd28134,17'd32018,17'd29979,17'd29979,17'd29978,17'd30130,17'd30885,17'd30739,17'd29833,17'd29249,17'd31196,17'd29691,17'd29690,17'd29690,17'd28857,17'd28857,17'd28857,17'd28857,17'd29690,17'd29690,17'd29536,17'd38154,17'd46837,17'd41412,17'd47938,17'd47054,17'd47737,17'd51648,17'd53048,17'd52979,17'd52749,17'd52000,17'd51390,17'd48360,17'd47443,17'd53049,17'd53050,17'd53051,17'd25566,17'd25435,17'd41730,17'd29688,17'd29376,17'd23217,17'd34458,17'd51314,17'd45037,17'd23217,17'd31033,17'd24742,17'd25180,17'd30126,17'd23733,17'd30425,17'd36566,17'd30728,17'd39441,17'd36566,17'd32666,17'd31831,17'd51543,17'd53052,17'd21538,17'd52680,17'd52347,17'd42888,17'd43841,17'd33946,17'd50740,17'd35014,17'd53053,17'd48159,17'd47150,17'd51482,17'd53054,17'd53055,17'd35882,17'd19695,17'd21918,17'd24299,17'd29157,17'd52994,17'd7007,17'd25225,17'd5914,17'd5916,17'd5759,17'd4993,17'd53056,17'd52906,17'd5477,17'd4676,17'd4682,17'd4686,17'd25627,17'd27935,17'd6219,17'd6220,17'd7499,17'd27696,17'd35052,17'd32074,17'd37152,17'd6554,17'd6554,17'd6554,17'd28185,17'd28185,17'd6554,17'd6390,17'd32073,17'd9091,17'd32074,17'd29740,17'd29740,17'd29740,17'd7499,17'd7499,17'd7668,17'd9091,17'd6390,17'd27935,17'd30638,17'd5004,17'd25627,17'd5335,17'd37434,17'd5616,17'd35197,17'd52763,17'd50836,17'd53057,17'd47081,17'd53058,17'd53059,17'd36742,17'd53060,17'd29744,17'd53061,17'd53062,17'd53063,17'd53064,17'd53065,17'd53066,17'd3061,17'd52772,17'd53067,17'd4053,17'd3707,17'd4056,17'd48812,17'd5354,17'd5026,17'd5026,17'd5496,17'd53068,17'd53068,17'd3426,17'd3426,17'd1824,17'd2391,17'd2558,17'd38071,17'd4059,17'd628,17'd628,17'd630,17'd960,17'd52698,17'd4059,17'd1121,17'd3071,17'd36322,17'd52919,17'd53069,17'd52921,17'd53070,17'd53071,17'd53072,17'd53073,17'd53011,17'd53074
},
'{
17'd53075,17'd5204,17'd11609,17'd3752,17'd17187,17'd17,17'd652,17'd27,17'd285,17'd285,17'd285,17'd467,17'd467,17'd467,17'd467,17'd467,17'd7385,17'd7385,17'd7060,17'd7060,17'd4430,17'd4430,17'd4431,17'd3907,17'd3907,17'd9816,17'd3756,17'd3435,17'd4250,17'd5210,17'd5806,17'd32729,17'd5381,17'd4586,17'd12658,17'd53076,17'd29043,17'd53077,17'd5066,17'd26130,17'd53016,17'd23320,17'd12046,17'd12345,17'd15508,17'd16403,17'd53078,17'd18532,17'd12954,17'd12678,17'd12678,17'd13092,17'd13598,17'd15762,17'd12356,17'd13597,17'd12357,17'd14469,17'd14763,17'd50503,17'd14620,17'd14620,17'd14620,17'd52468,17'd12675,17'd13460,17'd12357,17'd13209,17'd21184,17'd13092,17'd12678,17'd12527,17'd12527,17'd13094,17'd22630,17'd19382,17'd53079,17'd23155,17'd18533,17'd18174,17'd18774,17'd21649,17'd16410,17'd13469,17'd14623,17'd47973,17'd49200,17'd53080,17'd53081,17'd53082,17'd3633,17'd4288,17'd3138,17'd3468,17'd5844,17'd53083,17'd53084,17'd53085,17'd53086,17'd53087,17'd52550,17'd53088,17'd53089,17'd43891,17'd41925,17'd51022,17'd53090,17'd6649,17'd53091,17'd43075,17'd52936,17'd53092,17'd52477,17'd53093,17'd52118,17'd30061,17'd27841,17'd27724,17'd53094,17'd26027,17'd22123,17'd52291,17'd17956,17'd10446,17'd16674,17'd52716,17'd26252,17'd53095,17'd15165,17'd53096,17'd53097,17'd11381,17'd11381,17'd11382,17'd27116,17'd53098,17'd52863,17'd11511,17'd18438,17'd11796,17'd11796,17'd15561,17'd13756,17'd53099,17'd53100,17'd53101,17'd17349,17'd53102,17'd18563,17'd19413,17'd14809,17'd13518,17'd13518,17'd13252,17'd15685,17'd17603,17'd18917,17'd12996,17'd19158,17'd18443,17'd20609,17'd21505,17'd24857,17'd30831,17'd31941,17'd31589,17'd50951,17'd52133,17'd52869,17'd52868,17'd52869,17'd52799,17'd53103,17'd52133,17'd51881,17'd50952,17'd31590,17'd32283,17'd31439,17'd28461,17'd26370,17'd24209,17'd25143,17'd30532,17'd24029,17'd11274,17'd11274,17'd11274,17'd11274,17'd11808,17'd11129,17'd22647,17'd17236,17'd16068,17'd11806,17'd12419,17'd12419,17'd13764,17'd31130,17'd33083,17'd53104,17'd53105,17'd8724,17'd23860,17'd10173,17'd16549,17'd12116,17'd10479,17'd11132,17'd14810,17'd16069,17'd11666,17'd13764,17'd13363,17'd12109,17'd12579,17'd12417,17'd12856,17'd12110,17'd18679,17'd16064,17'd18915,17'd10163,17'd24038,17'd53106,17'd16072,17'd8252,17'd19780,17'd53107,17'd35514,17'd33404,17'd16071,17'd9040,17'd9040,17'd12264,17'd8100,17'd8580,17'd17127,17'd53108,17'd53109,17'd53110,17'd53111,17'd12870,17'd53112,17'd10874,17'd140,17'd132,17'd11541,17'd133,17'd542,17'd1197,17'd132,17'd5593,17'd131,17'd133,17'd23537,17'd53113,17'd53114,17'd53115,17'd22864,17'd45746,17'd50156,17'd46548,17'd53116,17'd53117,17'd49572,17'd53118,17'd41858,17'd50268,17'd51741,17'd50476,17'd50736,17'd50476,17'd50476,17'd51741,17'd50268,17'd41721,17'd41579,17'd38971,17'd42298,17'd35152,17'd32832,17'd28134,17'd32017,17'd32507,17'd32193,17'd33656,17'd33486,17'd37118,17'd36988,17'd32193,17'd36989,17'd53119,17'd50906,17'd29106,17'd53120,17'd53121,17'd29247,17'd29537,17'd29979,17'd29690,17'd49790,17'd30280,17'd30736,17'd31036,17'd29831,17'd28371,17'd28256,17'd29380,17'd28857,17'd49579,17'd53122,17'd28372,17'd28372,17'd29380,17'd28857,17'd32833,17'd33486,17'd33320,17'd53123,17'd53124,17'd53125,17'd43148,17'd47344,17'd49484,17'd50568,17'd52675,17'd52821,17'd52891,17'd51995,17'd41721,17'd41105,17'd53126,17'd53127,17'd52343,17'd32996,17'd25566,17'd43022,17'd30432,17'd31033,17'd30128,17'd39131,17'd36009,17'd35018,17'd39132,17'd23566,17'd24743,17'd24745,17'd32007,17'd34883,17'd29530,17'd39131,17'd34638,17'd53128,17'd35157,17'd32666,17'd49096,17'd21697,17'd53129,17'd53130,17'd21383,17'd53131,17'd46775,17'd21530,17'd52344,17'd50740,17'd35154,17'd42602,17'd50999,17'd53132,17'd53133,17'd53134,17'd53135,17'd53136,17'd23432,17'd21446,17'd53137,17'd23968,17'd53138,17'd26215,17'd24480,17'd6382,17'd6845,17'd6846,17'd6382,17'd6381,17'd33365,17'd52906,17'd6210,17'd6381,17'd4840,17'd5005,17'd28185,17'd6554,17'd32073,17'd9091,17'd29740,17'd27696,17'd7499,17'd32073,17'd31717,17'd27935,17'd5614,17'd27935,17'd31717,17'd31717,17'd6554,17'd6390,17'd6390,17'd6219,17'd7499,17'd7499,17'd7499,17'd9091,17'd29740,17'd27696,17'd29740,17'd7499,17'd6219,17'd27935,17'd25627,17'd30637,17'd30333,17'd30333,17'd6853,17'd35197,17'd53139,17'd53140,17'd53141,17'd52355,17'd47081,17'd53000,17'd53142,17'd52911,17'd2879,17'd35484,17'd53143,17'd53144,17'd53145,17'd53146,17'd53147,17'd2545,17'd53148,17'd52460,17'd51252,17'd49712,17'd53006,17'd40099,17'd4709,17'd4865,17'd18142,17'd18142,17'd4557,17'd4399,17'd53149,17'd53150,17'd1825,17'd1825,17'd2391,17'd2558,17'd628,17'd628,17'd3874,17'd53151,17'd630,17'd630,17'd796,17'd6239,17'd3711,17'd6084,17'd53152,17'd53007,17'd53153,17'd53154,17'd53155,17'd53156,17'd53157,17'd53158,17'd53011,17'd53159
},
'{
17'd53075,17'd15496,17'd11609,17'd3752,17'd17187,17'd17,17'd652,17'd27,17'd285,17'd285,17'd467,17'd467,17'd467,17'd467,17'd467,17'd467,17'd7385,17'd7385,17'd7060,17'd7060,17'd4430,17'd4430,17'd4431,17'd3907,17'd9816,17'd9816,17'd12335,17'd3435,17'd4250,17'd5210,17'd5806,17'd32729,17'd5381,17'd4897,17'd12509,17'd30503,17'd50758,17'd27828,17'd27100,17'd26349,17'd53160,17'd23146,17'd52545,17'd12665,17'd53161,17'd16510,17'd53162,17'd18532,17'd13599,17'd12527,17'd12678,17'd13092,17'd13598,17'd15762,17'd13597,17'd13597,17'd12357,17'd14469,17'd14763,17'd50503,17'd14620,17'd14620,17'd14620,17'd52468,17'd12675,17'd13460,17'd12357,17'd13209,17'd13210,17'd13599,17'd12527,17'd12527,17'd12527,17'd12955,17'd14471,17'd28438,17'd53079,17'd23155,17'd18533,17'd18174,17'd27461,17'd21649,17'd16410,17'd13470,17'd13468,17'd48081,17'd49200,17'd53080,17'd53163,17'd53164,17'd3634,17'd53165,17'd3139,17'd3468,17'd2655,17'd53166,17'd53167,17'd41329,17'd53168,17'd53169,17'd52031,17'd44154,17'd53170,17'd43608,17'd53171,17'd51022,17'd53172,17'd6649,17'd53091,17'd53173,17'd49304,17'd53092,17'd50507,17'd53174,17'd53175,17'd53176,17'd28557,17'd27842,17'd9595,17'd20598,17'd52122,17'd53177,17'd10302,17'd53178,17'd52558,17'd16541,17'd16900,17'd52857,17'd15668,17'd53179,17'd53180,17'd52859,17'd53181,17'd16547,17'd16547,17'd11384,17'd11951,17'd52863,17'd18438,17'd13998,17'd11798,17'd11796,17'd53182,17'd53183,17'd53184,17'd53185,17'd40744,17'd40284,17'd53102,17'd16914,17'd13643,17'd13760,17'd14809,17'd14526,17'd15433,17'd17603,17'd15053,17'd12996,17'd15185,17'd18443,17'd18443,17'd22992,17'd24031,17'd53186,17'd32919,17'd32592,17'd50111,17'd51959,17'd52869,17'd52869,17'd52402,17'd52648,17'd53103,17'd53187,17'd52132,17'd51958,17'd35239,17'd33720,17'd30834,17'd31587,17'd28943,17'd24537,17'd21363,17'd24994,17'd19533,17'd11808,17'd10990,17'd14931,17'd14673,17'd11274,17'd13645,17'd11275,17'd10476,17'd14931,17'd15185,17'd11959,17'd12580,17'd13882,17'd15182,17'd20756,17'd17600,17'd53188,17'd8410,17'd23861,17'd9194,17'd10173,17'd9619,17'd10479,17'd11133,17'd13886,17'd12720,17'd13000,17'd13764,17'd13882,17'd12109,17'd12579,17'd12417,17'd12856,17'd12110,17'd12111,17'd18679,17'd18805,17'd10736,17'd10856,17'd14675,17'd8419,17'd25680,17'd15301,17'd53189,17'd12119,17'd8730,17'd50864,17'd8877,17'd8567,17'd8728,17'd17481,17'd8580,17'd17240,17'd23687,17'd53190,17'd16448,17'd53191,17'd26042,17'd16925,17'd13533,17'd132,17'd132,17'd132,17'd133,17'd542,17'd133,17'd131,17'd11683,17'd5593,17'd131,17'd24056,17'd23538,17'd52963,17'd46678,17'd33312,17'd53192,17'd53193,17'd43285,17'd50068,17'd53194,17'd53195,17'd53196,17'd42432,17'd53197,17'd50371,17'd50273,17'd50273,17'd50273,17'd50272,17'd50476,17'd49794,17'd53198,17'd47930,17'd44933,17'd34275,17'd32832,17'd28134,17'd28134,17'd32017,17'd32017,17'd32193,17'd32507,17'd33486,17'd37118,17'd53199,17'd36847,17'd29833,17'd50570,17'd49686,17'd29380,17'd53200,17'd53201,17'd29691,17'd29979,17'd29979,17'd49790,17'd30131,17'd30280,17'd30736,17'd30736,17'd28857,17'd28133,17'd28255,17'd28257,17'd28857,17'd49579,17'd53122,17'd28372,17'd28257,17'd29380,17'd28857,17'd33166,17'd29248,17'd35990,17'd45612,17'd53202,17'd47938,17'd46761,17'd48264,17'd49891,17'd52000,17'd52169,17'd52749,17'd52820,17'd51916,17'd39423,17'd47529,17'd50821,17'd53203,17'd43285,17'd28721,17'd28721,17'd28484,17'd32007,17'd23918,17'd22501,17'd22332,17'd36009,17'd33949,17'd42744,17'd23384,17'd28718,17'd24898,17'd32007,17'd30431,17'd23388,17'd39131,17'd33645,17'd48367,17'd30728,17'd32009,17'd44824,17'd53204,17'd53205,17'd53206,17'd53207,17'd53131,17'd51303,17'd21531,17'd51464,17'd35293,17'd42602,17'd42747,17'd53208,17'd53209,17'd53210,17'd53211,17'd53212,17'd53213,17'd20091,17'd21916,17'd22735,17'd24301,17'd24942,17'd26215,17'd24480,17'd6382,17'd6845,17'd7661,17'd23975,17'd24795,17'd52906,17'd33365,17'd52995,17'd5323,17'd4686,17'd5002,17'd28185,17'd32073,17'd32074,17'd32074,17'd29740,17'd7668,17'd6219,17'd6390,17'd28185,17'd27935,17'd5614,17'd27935,17'd31717,17'd31717,17'd6554,17'd6390,17'd6390,17'd6219,17'd7499,17'd7499,17'd7499,17'd9091,17'd29740,17'd27696,17'd31888,17'd32074,17'd6219,17'd5336,17'd5002,17'd30637,17'd30638,17'd31891,17'd53214,17'd35197,17'd53215,17'd4374,17'd39618,17'd51846,17'd53216,17'd53058,17'd52607,17'd47378,17'd53217,17'd53218,17'd53219,17'd53144,17'd53220,17'd53221,17'd40096,17'd51182,17'd41622,17'd52772,17'd51412,17'd49712,17'd53006,17'd3871,17'd4709,17'd4865,17'd5026,17'd18142,17'd52020,17'd38718,17'd53222,17'd53068,17'd1825,17'd1825,17'd2558,17'd4398,17'd628,17'd628,17'd3874,17'd3222,17'd630,17'd1121,17'd3390,17'd6239,17'd10072,17'd2557,17'd53152,17'd52773,17'd53153,17'd53223,17'd53224,17'd53225,17'd53157,17'd53226,17'd53227,17'd53159
},
'{
17'd53228,17'd15496,17'd11609,17'd3752,17'd9969,17'd17,17'd652,17'd27,17'd285,17'd285,17'd467,17'd467,17'd467,17'd467,17'd467,17'd467,17'd7385,17'd7385,17'd7060,17'd7060,17'd4430,17'd4430,17'd4431,17'd4431,17'd3907,17'd3907,17'd3756,17'd3434,17'd5210,17'd5658,17'd5806,17'd32729,17'd5381,17'd53229,17'd12658,17'd30503,17'd50758,17'd12340,17'd26980,17'd26349,17'd49409,17'd53230,17'd52545,17'd12665,17'd52546,17'd52847,17'd19381,17'd18172,17'd13210,17'd12527,17'd12677,17'd12678,17'd13092,17'd12678,17'd12357,17'd12357,17'd12062,17'd12357,17'd14763,17'd50503,17'd14620,17'd14620,17'd14620,17'd52468,17'd14620,17'd12214,17'd12062,17'd13209,17'd13210,17'd13599,17'd12527,17'd12527,17'd12527,17'd12955,17'd14471,17'd28554,17'd18884,17'd28205,17'd19753,17'd53231,17'd18655,17'd21649,17'd16410,17'd16880,17'd13721,17'd47974,17'd52850,17'd53080,17'd53232,17'd53081,17'd53233,17'd53234,17'd3139,17'd2984,17'd2655,17'd53235,17'd53236,17'd6324,17'd51771,17'd53168,17'd52031,17'd44154,17'd53170,17'd43206,17'd43891,17'd41925,17'd53172,17'd6649,17'd53091,17'd53173,17'd49304,17'd53237,17'd53238,17'd38227,17'd49719,17'd53239,17'd30061,17'd50401,17'd27223,17'd22289,17'd19910,17'd22123,17'd10137,17'd52213,17'd52039,17'd20600,17'd52716,17'd15932,17'd52639,17'd27115,17'd53240,17'd53241,17'd53242,17'd53242,17'd16547,17'd11384,17'd53243,17'd11951,17'd13998,17'd11799,17'd18912,17'd22470,17'd53244,17'd53245,17'd53246,17'd53247,17'd46154,17'd17233,17'd17013,17'd16560,17'd14523,17'd13643,17'd13643,17'd14809,17'd15570,17'd15685,17'd12719,17'd13135,17'd16442,17'd16442,17'd18443,17'd21361,17'd53248,17'd37341,17'd30527,17'd31762,17'd34545,17'd51512,17'd53187,17'd52800,17'd52869,17'd52799,17'd53249,17'd53249,17'd52800,17'd51881,17'd51694,17'd53250,17'd33568,17'd30972,17'd30673,17'd28570,17'd24992,17'd22472,17'd30532,17'd11275,17'd10990,17'd14931,17'd14810,17'd14810,17'd10989,17'd10989,17'd10475,17'd10854,17'd13762,17'd13883,17'd12580,17'd14131,17'd28108,17'd31130,17'd16065,17'd16681,17'd31444,17'd8886,17'd9041,17'd9743,17'd17011,17'd11134,17'd10165,17'd10476,17'd14810,17'd11520,17'd12861,17'd13882,17'd12414,17'd12109,17'd12417,17'd12856,17'd12110,17'd12111,17'd18679,17'd53251,17'd15047,17'd25928,17'd9039,17'd8247,17'd53252,17'd33716,17'd17128,17'd13648,17'd19923,17'd53253,17'd29637,17'd9348,17'd22473,17'd8574,17'd10028,17'd13258,17'd23519,17'd22133,17'd53254,17'd53255,17'd17610,17'd53256,17'd53257,17'd53258,17'd13777,17'd133,17'd542,17'd542,17'd133,17'd132,17'd5593,17'd5593,17'd131,17'd53259,17'd53260,17'd51222,17'd35015,17'd53261,17'd51735,17'd52888,17'd53262,17'd53263,17'd53264,17'd53265,17'd49484,17'd50160,17'd51830,17'd50661,17'd42875,17'd42875,17'd51163,17'd51830,17'd50996,17'd41410,17'd49276,17'd48894,17'd43980,17'd35707,17'd27885,17'd28134,17'd28134,17'd28373,17'd28134,17'd33654,17'd32507,17'd29249,17'd29691,17'd49687,17'd29979,17'd49789,17'd49789,17'd29831,17'd31196,17'd53266,17'd29106,17'd29690,17'd29978,17'd30131,17'd49790,17'd30280,17'd30736,17'd31036,17'd29978,17'd30587,17'd26522,17'd28370,17'd28372,17'd29536,17'd28857,17'd29380,17'd28256,17'd28256,17'd29380,17'd29106,17'd33486,17'd33165,17'd38974,17'd53267,17'd53268,17'd43282,17'd48709,17'd48263,17'd50365,17'd52671,17'd52749,17'd52675,17'd53197,17'd51648,17'd53269,17'd47338,17'd50651,17'd50361,17'd43835,17'd28721,17'd28721,17'd29103,17'd23916,17'd23566,17'd23389,17'd22857,17'd36009,17'd41419,17'd23923,17'd24902,17'd24417,17'd25180,17'd28368,17'd31033,17'd29374,17'd30425,17'd34278,17'd39281,17'd32503,17'd32009,17'd21849,17'd47359,17'd53270,17'd53271,17'd52593,17'd21705,17'd51551,17'd51230,17'd42153,17'd52086,17'd53272,17'd42305,17'd53273,17'd22869,17'd53274,17'd53275,17'd53276,17'd53277,17'd23778,17'd22235,17'd22408,17'd22584,17'd25877,17'd11158,17'd24480,17'd5610,17'd5914,17'd6383,17'd24647,17'd53278,17'd53279,17'd53280,17'd24795,17'd5323,17'd4845,17'd5160,17'd27935,17'd6390,17'd9091,17'd32074,17'd7499,17'd7499,17'd6219,17'd6554,17'd6554,17'd6390,17'd6390,17'd6554,17'd31717,17'd31717,17'd6554,17'd6390,17'd32073,17'd9091,17'd7499,17'd7499,17'd9091,17'd9091,17'd29740,17'd27696,17'd9933,17'd9091,17'd5615,17'd5336,17'd4842,17'd30180,17'd30638,17'd52270,17'd5338,17'd5013,17'd53281,17'd53282,17'd51094,17'd53283,17'd47082,17'd53284,17'd36742,17'd53285,17'd53286,17'd53287,17'd53288,17'd53289,17'd53220,17'd53290,17'd40096,17'd53291,17'd41477,17'd52772,17'd51855,17'd53292,17'd50089,17'd3871,17'd4709,17'd10906,17'd5026,17'd18142,17'd5496,17'd53293,17'd53222,17'd4399,17'd1824,17'd1824,17'd2558,17'd38071,17'd628,17'd1120,17'd3711,17'd53294,17'd235,17'd448,17'd3874,17'd4228,17'd10072,17'd2557,17'd53152,17'd18758,17'd53295,17'd53223,17'd53296,17'd53225,17'd53157,17'd53158,17'd53297,17'd53012
},
'{
17'd53228,17'd3592,17'd11609,17'd3752,17'd9969,17'd17,17'd652,17'd27,17'd285,17'd285,17'd467,17'd467,17'd467,17'd467,17'd467,17'd467,17'd7385,17'd7385,17'd7060,17'd7060,17'd4430,17'd4430,17'd4431,17'd4431,17'd3907,17'd3907,17'd3756,17'd3434,17'd5210,17'd5658,17'd5806,17'd32729,17'd5381,17'd4898,17'd12509,17'd30503,17'd3270,17'd3764,17'd27100,17'd48472,17'd21337,17'd53298,17'd24338,17'd12665,17'd21179,17'd14760,17'd53299,17'd53300,17'd19890,17'd12679,17'd12677,17'd12677,17'd12678,17'd13092,17'd14469,17'd12357,17'd12062,17'd12357,17'd14763,17'd50503,17'd13460,17'd13460,17'd14620,17'd14620,17'd14620,17'd12214,17'd12062,17'd13209,17'd13210,17'd13599,17'd12527,17'd12527,17'd12527,17'd12955,17'd13969,17'd28438,17'd28205,17'd28205,17'd19753,17'd53231,17'd18655,17'd16986,17'd16410,17'd16880,17'd13721,17'd14625,17'd48298,17'd53080,17'd53301,17'd53163,17'd53302,17'd3957,17'd53303,17'd2984,17'd2655,17'd53304,17'd53305,17'd6155,17'd52204,17'd53168,17'd52031,17'd44154,17'd42352,17'd44283,17'd44522,17'd41925,17'd53306,17'd53090,17'd53307,17'd43075,17'd42354,17'd46900,17'd53308,17'd53309,17'd52633,17'd52118,17'd53310,17'd53311,17'd27223,17'd52121,17'd53312,17'd53313,17'd18905,17'd18432,17'd20896,17'd10581,17'd16541,17'd17004,17'd51686,17'd53314,17'd52717,17'd53240,17'd11380,17'd26490,17'd17713,17'd26997,17'd26624,17'd26624,17'd11794,17'd11947,17'd12246,17'd11945,17'd53315,17'd53316,17'd53317,17'd53318,17'd53319,17'd32445,17'd17014,17'd17014,17'd14672,17'd14523,17'd13643,17'd14809,17'd13517,17'd13252,17'd11958,17'd15053,17'd22472,17'd22472,17'd22472,17'd22472,17'd26035,17'd46382,17'd30831,17'd30833,17'd32592,17'd50863,17'd53187,17'd53320,17'd52799,17'd53321,17'd53322,17'd53323,17'd53320,17'd53324,17'd51602,17'd34705,17'd33720,17'd30677,17'd29779,17'd29475,17'd28110,17'd21505,17'd24994,17'd24029,17'd11275,17'd10990,17'd14810,17'd14810,17'd10989,17'd14931,17'd10476,17'd10990,17'd11964,17'd13135,17'd12420,17'd14131,17'd16323,17'd52726,17'd15681,17'd10335,17'd16681,17'd9621,17'd10174,17'd10335,17'd9479,17'd12116,17'd17719,17'd10326,17'd13886,17'd16068,17'd11667,17'd13364,17'd16443,17'd12580,17'd12253,17'd12417,17'd12580,17'd12419,17'd13363,17'd16322,17'd28108,17'd17121,17'd16070,17'd9045,17'd33570,17'd35089,17'd9889,17'd53325,17'd8419,17'd8575,17'd24999,17'd9348,17'd12425,17'd24710,17'd8733,17'd17352,17'd17128,17'd9197,17'd22996,17'd21828,17'd20181,17'd53326,17'd53327,17'd22487,17'd20188,17'd1045,17'd542,17'd542,17'd1481,17'd132,17'd11683,17'd5593,17'd53328,17'd51623,17'd53329,17'd51654,17'd31658,17'd53330,17'd53331,17'd53332,17'd53333,17'd46434,17'd53334,17'd53335,17'd49683,17'd51830,17'd52000,17'd43012,17'd50660,17'd43146,17'd51652,17'd50272,17'd51078,17'd39122,17'd47930,17'd53336,17'd33476,17'd32832,17'd32192,17'd33654,17'd28258,17'd32832,17'd27885,17'd32354,17'd32507,17'd33166,17'd49579,17'd30131,17'd30736,17'd30738,17'd30130,17'd29536,17'd29106,17'd53337,17'd29979,17'd29978,17'd30131,17'd30131,17'd30131,17'd30736,17'd30736,17'd30738,17'd28857,17'd53338,17'd53339,17'd28257,17'd28857,17'd28857,17'd28372,17'd28257,17'd28255,17'd28255,17'd29380,17'd29106,17'd32507,17'd40219,17'd43700,17'd53340,17'd48147,17'd48616,17'd49586,17'd49478,17'd51157,17'd53341,17'd52749,17'd52671,17'd50468,17'd43541,17'd53342,17'd53126,17'd50157,17'd53333,17'd43550,17'd44229,17'd43022,17'd29976,17'd30879,17'd29686,17'd39131,17'd22858,17'd31656,17'd29973,17'd23565,17'd29100,17'd24896,17'd29976,17'd28977,17'd30275,17'd29975,17'd41273,17'd45754,17'd39441,17'd32503,17'd47834,17'd36129,17'd53343,17'd51982,17'd53271,17'd53344,17'd51304,17'd21529,17'd51464,17'd42602,17'd52086,17'd53345,17'd42439,17'd53346,17'd47154,17'd53347,17'd53348,17'd53349,17'd53350,17'd43314,17'd53351,17'd23787,17'd24303,17'd25221,17'd10196,17'd6211,17'd5610,17'd5913,17'd6212,17'd5322,17'd52906,17'd52906,17'd52995,17'd53352,17'd5325,17'd5330,17'd5335,17'd6390,17'd9091,17'd32074,17'd32074,17'd9091,17'd9091,17'd6390,17'd6554,17'd6390,17'd6390,17'd6390,17'd6554,17'd31717,17'd31717,17'd6390,17'd6390,17'd9091,17'd9091,17'd7499,17'd7499,17'd9091,17'd9091,17'd29740,17'd27696,17'd9933,17'd32073,17'd5615,17'd5160,17'd28536,17'd30180,17'd30638,17'd52270,17'd5338,17'd53353,17'd53354,17'd49706,17'd53355,17'd53356,17'd53357,17'd53358,17'd48182,17'd43737,17'd53359,17'd53360,17'd53361,17'd53362,17'd53363,17'd53290,17'd40096,17'd51182,17'd41622,17'd52772,17'd41158,17'd42043,17'd4055,17'd48812,17'd18512,17'd10906,17'd5026,17'd5495,17'd38718,17'd53293,17'd53150,17'd52918,17'd1824,17'd1824,17'd4398,17'd4059,17'd628,17'd1120,17'd3711,17'd53364,17'd235,17'd796,17'd6239,17'd4228,17'd10072,17'd2557,17'd53152,17'd52773,17'd33846,17'd53070,17'd53365,17'd53225,17'd53157,17'd53226,17'd53366,17'd53012
},
'{
17'd53228,17'd3592,17'd11609,17'd3752,17'd9969,17'd17,17'd652,17'd27,17'd285,17'd285,17'd467,17'd467,17'd467,17'd467,17'd467,17'd467,17'd7385,17'd7385,17'd7060,17'd7060,17'd4430,17'd4430,17'd4431,17'd4431,17'd3907,17'd3907,17'd11210,17'd3434,17'd5379,17'd5657,17'd5806,17'd32729,17'd5381,17'd53229,17'd4261,17'd32410,17'd50389,17'd3272,17'd3608,17'd48472,17'd53367,17'd13699,17'd24338,17'd52109,17'd53368,17'd53369,17'd16511,17'd53300,17'd18411,17'd12955,17'd35352,17'd11625,17'd12678,17'd14469,17'd14469,17'd12357,17'd12357,17'd14469,17'd14763,17'd50503,17'd11084,17'd11084,17'd13460,17'd14620,17'd14620,17'd12214,17'd12062,17'd13209,17'd12955,17'd12955,17'd12679,17'd12527,17'd12813,17'd13211,17'd13969,17'd22630,17'd18884,17'd28205,17'd17941,17'd19753,17'd18655,17'd18774,17'd16986,17'd20585,17'd13721,17'd48474,17'd47972,17'd34178,17'd50094,17'd53370,17'd53302,17'd3477,17'd3302,17'd3467,17'd53371,17'd53372,17'd53373,17'd53374,17'd53375,17'd53376,17'd52031,17'd44154,17'd53377,17'd42800,17'd42936,17'd6648,17'd51022,17'd41333,17'd50096,17'd43075,17'd42354,17'd45669,17'd53378,17'd50507,17'd37597,17'd53379,17'd53380,17'd51781,17'd27222,17'd22805,17'd20302,17'd53381,17'd19147,17'd10137,17'd52038,17'd18186,17'd53382,17'd53383,17'd52560,17'd26619,17'd10963,17'd53384,17'd53385,17'd26490,17'd17713,17'd16547,17'd11383,17'd18075,17'd12851,17'd12099,17'd23335,17'd11946,17'd53386,17'd52864,17'd53387,17'd53388,17'd53389,17'd53390,17'd53391,17'd17234,17'd13642,17'd32138,17'd14930,17'd13643,17'd13517,17'd13252,17'd11958,17'd12719,17'd18197,17'd18197,17'd22472,17'd22472,17'd53392,17'd41187,17'd30218,17'd35931,17'd30834,17'd35093,17'd52867,17'd52800,17'd53321,17'd53321,17'd53322,17'd53393,17'd53322,17'd52799,17'd52302,17'd53394,17'd34545,17'd33568,17'd30972,17'd30829,17'd33726,17'd28111,17'd23167,17'd21985,17'd11275,17'd11808,17'd14931,17'd14931,17'd14931,17'd14931,17'd10605,17'd10990,17'd10989,17'd11963,17'd11958,17'd12110,17'd14808,17'd53395,17'd26630,17'd26759,17'd20757,17'd17471,17'd15944,17'd15807,17'd9620,17'd9741,17'd16796,17'd10166,17'd11132,17'd14931,17'd11520,17'd13363,17'd14131,17'd12109,17'd12579,17'd14807,17'd12580,17'd12419,17'd13761,17'd14808,17'd15564,17'd11666,17'd10605,17'd9479,17'd11404,17'd53396,17'd15694,17'd17129,17'd14527,17'd12867,17'd9046,17'd9195,17'd36205,17'd53397,17'd53398,17'd24044,17'd19418,17'd14005,17'd53399,17'd14010,17'd14266,17'd20183,17'd53400,17'd53401,17'd53402,17'd17363,17'd717,17'd542,17'd130,17'd132,17'd5593,17'd11683,17'd52810,17'd53403,17'd53404,17'd35709,17'd45874,17'd53405,17'd52888,17'd52967,17'd52426,17'd51234,17'd53406,17'd53407,17'd50568,17'd52000,17'd43146,17'd53408,17'd43012,17'd51236,17'd53409,17'd53410,17'd41097,17'd53411,17'd44226,17'd39740,17'd32356,17'd33164,17'd33654,17'd32017,17'd28258,17'd31354,17'd31503,17'd32354,17'd29380,17'd30884,17'd30131,17'd30280,17'd31036,17'd30738,17'd29979,17'd30884,17'd30884,17'd29690,17'd30130,17'd30280,17'd30131,17'd30131,17'd30280,17'd30736,17'd30736,17'd29978,17'd33321,17'd53412,17'd28981,17'd28372,17'd28857,17'd31196,17'd28257,17'd28255,17'd53413,17'd27884,17'd32507,17'd33656,17'd32355,17'd34450,17'd45481,17'd43421,17'd43282,17'd48709,17'd48536,17'd49788,17'd51830,17'd52749,17'd52749,17'd51830,17'd49691,17'd45368,17'd49271,17'd50821,17'd53414,17'd50153,17'd43694,17'd43550,17'd43553,17'd24745,17'd23384,17'd29828,17'd41419,17'd35018,17'd30129,17'd32191,17'd24086,17'd28601,17'd24745,17'd25031,17'd35159,17'd34137,17'd29828,17'd23389,17'd22680,17'd22333,17'd22159,17'd44701,17'd35855,17'd53415,17'd53131,17'd51991,17'd51225,17'd51563,17'd42153,17'd51230,17'd53416,17'd53417,17'd51633,17'd51066,17'd53418,17'd46851,17'd53419,17'd53420,17'd53421,17'd53422,17'd53423,17'd29021,17'd22583,17'd53424,17'd12443,17'd26449,17'd6549,17'd5611,17'd5609,17'd4994,17'd24148,17'd53425,17'd33365,17'd24796,17'd6067,17'd4840,17'd5330,17'd5336,17'd6219,17'd9091,17'd29740,17'd29740,17'd9091,17'd32073,17'd6554,17'd6554,17'd6219,17'd6390,17'd6390,17'd6554,17'd36586,17'd36586,17'd32073,17'd9091,17'd9091,17'd7499,17'd7499,17'd7499,17'd9091,17'd9091,17'd29740,17'd27696,17'd8780,17'd6390,17'd5615,17'd5004,17'd31716,17'd30637,17'd37030,17'd50282,17'd5616,17'd53426,17'd53427,17'd53428,17'd50837,17'd51095,17'd47082,17'd53429,17'd53430,17'd53431,17'd53432,17'd23472,17'd53433,17'd53434,17'd53435,17'd2225,17'd41312,17'd20559,17'd41477,17'd52019,17'd3866,17'd53292,17'd50185,17'd3709,17'd4553,17'd18142,17'd52020,17'd38857,17'd53068,17'd53222,17'd53068,17'd5497,17'd2558,17'd2558,17'd4398,17'd4059,17'd3874,17'd3874,17'd18144,17'd52461,17'd235,17'd796,17'd4059,17'd38071,17'd3874,17'd2557,17'd53152,17'd18758,17'd53436,17'd53437,17'd53365,17'd53438,17'd53439,17'd53226,17'd53366,17'd53440
},
'{
17'd53228,17'd3592,17'd11609,17'd3752,17'd9969,17'd1416,17'd652,17'd27,17'd285,17'd285,17'd467,17'd467,17'd467,17'd467,17'd467,17'd467,17'd7385,17'd7385,17'd7060,17'd7060,17'd4430,17'd4430,17'd4431,17'd4431,17'd3907,17'd3907,17'd11210,17'd3434,17'd5379,17'd5657,17'd5806,17'd32729,17'd5381,17'd4897,17'd33053,17'd30812,17'd29449,17'd49010,17'd27325,17'd14876,17'd53441,17'd53442,17'd53443,17'd19748,17'd53368,17'd53444,17'd53445,17'd20734,17'd53446,17'd14890,17'd12813,17'd35352,17'd12678,17'd14469,17'd14469,17'd12357,17'd12357,17'd14469,17'd14468,17'd50503,17'd11084,17'd11084,17'd13460,17'd14620,17'd14620,17'd12214,17'd12062,17'd13209,17'd14890,17'd12955,17'd12679,17'd12527,17'd13093,17'd13211,17'd13969,17'd20292,17'd28205,17'd28205,17'd17941,17'd19753,17'd18655,17'd16766,17'd16410,17'd20585,17'd13721,17'd14624,17'd47971,17'd34178,17'd50094,17'd53447,17'd53448,17'd53449,17'd3302,17'd3467,17'd3134,17'd2652,17'd53450,17'd6009,17'd43602,17'd53451,17'd45528,17'd6324,17'd6157,17'd43203,17'd53452,17'd43074,17'd51022,17'd50765,17'd50934,17'd43892,17'd53453,17'd48192,17'd40124,17'd53308,17'd53454,17'd53379,17'd8393,17'd28672,17'd27110,17'd26990,17'd53455,17'd25917,17'd53456,17'd18905,17'd53457,17'd53458,17'd53459,17'd53460,17'd53461,17'd26361,17'd53462,17'd53463,17'd53464,17'd53385,17'd26490,17'd17713,17'd26997,17'd15043,17'd11652,17'd12099,17'd13248,17'd12246,17'd25271,17'd53465,17'd53466,17'd53467,17'd53468,17'd53469,17'd53470,17'd17234,17'd16686,17'd13642,17'd14930,17'd14525,17'd12417,17'd12995,17'd12420,17'd12106,17'd18559,17'd19409,17'd22472,17'd22472,17'd20608,17'd26494,17'd27004,17'd30831,17'd39211,17'd32592,17'd51272,17'd53324,17'd53321,17'd53471,17'd53471,17'd53472,17'd53393,17'd53322,17'd52869,17'd53473,17'd35239,17'd33875,17'd31765,17'd29330,17'd28106,17'd30076,17'd24539,17'd23169,17'd19533,17'd11275,17'd11274,17'd14931,17'd14810,17'd12720,17'd10605,17'd10854,17'd10853,17'd12262,17'd12858,17'd12419,17'd14131,17'd19645,17'd26497,17'd15940,17'd9480,17'd53474,17'd10174,17'd14674,17'd9620,17'd16549,17'd12116,17'd21503,17'd10330,17'd13886,17'd14673,17'd11667,17'd15054,17'd15184,17'd14130,17'd12580,17'd12580,17'd12580,17'd13761,17'd14131,17'd14808,17'd18679,17'd13762,17'd10478,17'd16071,17'd53475,17'd16801,17'd53476,17'd10179,17'd10340,17'd25147,17'd24547,17'd53477,17'd26261,17'd53478,17'd24215,17'd53479,17'd9350,17'd14136,17'd14937,17'd15442,17'd20320,17'd53480,17'd53481,17'd22487,17'd7980,17'd888,17'd542,17'd128,17'd132,17'd5593,17'd53482,17'd53483,17'd53484,17'd53485,17'd44824,17'd51160,17'd33802,17'd53486,17'd53487,17'd50993,17'd49678,17'd53488,17'd53489,17'd51157,17'd51163,17'd43012,17'd43146,17'd43146,17'd51163,17'd53490,17'd41724,17'd40509,17'd44932,17'd42298,17'd35152,17'd32354,17'd53491,17'd33321,17'd32017,17'd32356,17'd31354,17'd31503,17'd28134,17'd29106,17'd49579,17'd33489,17'd31506,17'd30736,17'd30280,17'd49790,17'd29690,17'd29979,17'd30280,17'd30280,17'd30280,17'd30131,17'd30131,17'd30736,17'd30736,17'd30131,17'd30884,17'd53491,17'd33164,17'd29247,17'd28728,17'd31196,17'd28856,17'd28133,17'd28255,17'd47633,17'd27884,17'd32507,17'd32507,17'd40051,17'd40366,17'd45370,17'd43688,17'd47054,17'd49586,17'd49478,17'd50160,17'd51741,17'd52169,17'd52001,17'd50736,17'd48995,17'd49483,17'd49572,17'd49977,17'd48037,17'd43425,17'd43694,17'd43836,17'd33483,17'd34467,17'd23386,17'd23216,17'd36288,17'd31656,17'd29973,17'd23566,17'd29100,17'd23561,17'd24895,17'd28368,17'd30431,17'd23566,17'd29828,17'd23389,17'd22678,17'd22506,17'd35292,17'd50987,17'd35293,17'd51922,17'd53492,17'd53493,17'd53494,17'd51817,17'd21530,17'd35014,17'd53416,17'd53495,17'd53496,17'd51551,17'd53497,17'd53498,17'd53499,17'd53500,17'd53277,17'd53501,17'd22233,17'd53502,17'd23789,17'd53503,17'd53504,17'd7165,17'd5913,17'd5611,17'd5478,17'd4992,17'd53280,17'd53505,17'd53506,17'd6381,17'd4995,17'd4687,17'd5335,17'd27935,17'd9091,17'd9091,17'd29740,17'd29740,17'd9091,17'd32073,17'd6554,17'd6390,17'd6219,17'd6219,17'd6390,17'd6554,17'd36586,17'd32073,17'd32073,17'd9091,17'd7499,17'd7499,17'd7499,17'd7499,17'd9091,17'd9091,17'd29740,17'd27696,17'd8780,17'd6390,17'd5614,17'd30180,17'd31716,17'd5004,17'd5165,17'd50282,17'd5616,17'd5014,17'd51327,17'd53507,17'd53508,17'd53509,17'd46988,17'd53510,17'd45780,17'd53511,17'd24160,17'd53512,17'd53513,17'd53514,17'd53515,17'd2225,17'd41312,17'd53516,17'd20262,17'd52019,17'd3703,17'd42043,17'd5626,17'd41159,17'd5354,17'd18142,17'd5496,17'd38857,17'd53150,17'd53150,17'd53068,17'd5497,17'd2558,17'd4398,17'd38071,17'd38071,17'd5628,17'd3711,17'd3071,17'd3071,17'd235,17'd796,17'd4059,17'd53068,17'd6239,17'd2557,17'd53152,17'd52773,17'd53517,17'd53437,17'd53518,17'd53438,17'd53439,17'd53226,17'd53366,17'd53519
},
'{
17'd53228,17'd3592,17'd11609,17'd3429,17'd2936,17'd1416,17'd652,17'd27,17'd26,17'd285,17'd285,17'd467,17'd467,17'd2937,17'd467,17'd467,17'd7385,17'd7385,17'd7060,17'd7060,17'd4430,17'd4430,17'd4431,17'd4431,17'd6278,17'd6278,17'd11210,17'd3434,17'd5379,17'd5657,17'd5806,17'd32729,17'd5381,17'd4897,17'd32730,17'd33542,17'd24969,17'd49010,17'd48075,17'd14876,17'd46481,17'd14084,17'd53443,17'd23830,17'd53520,17'd16157,17'd18166,17'd53521,17'd53446,17'd12530,17'd12955,17'd15516,17'd12357,17'd14469,17'd14469,17'd12357,17'd22802,17'd22802,17'd22802,17'd11762,17'd11084,17'd11084,17'd13460,17'd14620,17'd14620,17'd12214,17'd10937,17'd13209,17'd14890,17'd12955,17'd12679,17'd12527,17'd13093,17'd13211,17'd13969,17'd22630,17'd20886,17'd28205,17'd17941,17'd17941,17'd18655,17'd17689,17'd16986,17'd20585,17'd13721,17'd14624,17'd48299,17'd34178,17'd50094,17'd53301,17'd53522,17'd53523,17'd53524,17'd3958,17'd3133,17'd2653,17'd53525,17'd53526,17'd43201,17'd6320,17'd42061,17'd43751,17'd53527,17'd53528,17'd53529,17'd6328,17'd51022,17'd50765,17'd50934,17'd43892,17'd53453,17'd48192,17'd47388,17'd48933,17'd53530,17'd53531,17'd53239,17'd49615,17'd51424,17'd53532,17'd25266,17'd23673,17'd53312,17'd53533,17'd10444,17'd17001,17'd53534,17'd53535,17'd19403,17'd15669,17'd10714,17'd53536,17'd53384,17'd53537,17'd53538,17'd53539,17'd17713,17'd26142,17'd11651,17'd12099,17'd12245,17'd12098,17'd21202,17'd24850,17'd53540,17'd53387,17'd53541,17'd53389,17'd53542,17'd17234,17'd16560,17'd16914,17'd15571,17'd14930,17'd13643,17'd13760,17'd12995,17'd13252,17'd17602,17'd19409,17'd21361,17'd22472,17'd21362,17'd23170,17'd24859,17'd29778,17'd29645,17'd31761,17'd50111,17'd51881,17'd53321,17'd53471,17'd53543,17'd53544,17'd53393,17'd53393,17'd53321,17'd53545,17'd52400,17'd35239,17'd31287,17'd30972,17'd30829,17'd29476,17'd28231,17'd21361,17'd19643,17'd14671,17'd11808,17'd11274,17'd14931,17'd12720,17'd14810,17'd10990,17'd10853,17'd18560,17'd18447,17'd12420,17'd12414,17'd14131,17'd53546,17'd26497,17'd19642,17'd15295,17'd9191,17'd25525,17'd9344,17'd16549,17'd11277,17'd18916,17'd17719,17'd14518,17'd10990,17'd11395,17'd15299,17'd13882,17'd13761,17'd11959,17'd16321,17'd12106,17'd11958,17'd12419,17'd14808,17'd13364,17'd18917,17'd12862,17'd53547,17'd8732,17'd53548,17'd7617,17'd48656,17'd16917,17'd26380,17'd11405,17'd26155,17'd23173,17'd37734,17'd24215,17'd7946,17'd34825,17'd25410,17'd15192,17'd19536,17'd53549,17'd53550,17'd53551,17'd53552,17'd52140,17'd888,17'd1481,17'd130,17'd132,17'd5593,17'd53553,17'd53554,17'd53555,17'd52086,17'd32999,17'd53556,17'd53557,17'd53558,17'd53559,17'd53126,17'd52256,17'd48995,17'd50365,17'd50371,17'd50739,17'd50660,17'd51236,17'd52974,17'd50072,17'd42589,17'd40356,17'd43971,17'd46205,17'd37658,17'd27885,17'd32192,17'd33655,17'd33654,17'd28373,17'd32832,17'd31503,17'd47633,17'd28256,17'd29536,17'd49790,17'd31506,17'd31506,17'd31506,17'd30280,17'd30131,17'd30131,17'd30280,17'd30736,17'd30736,17'd33489,17'd33323,17'd33489,17'd31036,17'd30736,17'd29690,17'd52889,17'd33164,17'd33319,17'd32017,17'd32507,17'd29105,17'd29105,17'd28370,17'd27761,17'd31503,17'd32832,17'd32507,17'd32505,17'd35990,17'd40519,17'd43283,17'd53560,17'd47936,17'd48263,17'd49788,17'd51157,17'd52001,17'd52169,17'd51163,17'd49891,17'd48361,17'd53561,17'd53562,17'd53127,17'd53563,17'd43835,17'd43694,17'd43553,17'd34276,17'd23732,17'd29975,17'd30425,17'd22859,17'd41419,17'd29828,17'd23918,17'd34884,17'd28718,17'd32007,17'd28977,17'd31033,17'd23387,17'd23215,17'd32827,17'd22855,17'd53564,17'd22507,17'd53565,17'd51303,17'd21537,17'd53566,17'd53567,17'd52438,17'd21533,17'd34880,17'd35293,17'd51901,17'd53568,17'd53569,17'd47947,17'd53570,17'd31535,17'd53571,17'd53572,17'd53573,17'd53574,17'd53575,17'd22218,17'd53576,17'd53577,17'd26327,17'd7009,17'd5913,17'd5609,17'd4840,17'd5144,17'd4186,17'd33041,17'd4523,17'd4681,17'd4840,17'd5002,17'd28185,17'd6554,17'd9091,17'd32074,17'd29740,17'd29740,17'd9091,17'd32073,17'd6390,17'd6219,17'd9091,17'd32073,17'd32073,17'd32073,17'd32073,17'd32073,17'd9091,17'd9091,17'd29740,17'd27696,17'd7668,17'd7499,17'd9091,17'd9091,17'd7499,17'd7499,17'd6391,17'd6390,17'd28185,17'd53578,17'd28536,17'd5160,17'd5164,17'd5338,17'd53353,17'd53579,17'd53580,17'd53581,17'd48805,17'd53582,17'd37565,17'd53583,17'd53584,17'd53585,17'd23985,17'd35057,17'd53513,17'd53586,17'd53587,17'd53588,17'd53589,17'd53590,17'd52614,17'd41478,17'd3703,17'd4054,17'd53591,17'd41159,17'd5495,17'd5496,17'd5496,17'd38857,17'd53150,17'd53150,17'd4399,17'd52918,17'd2558,17'd38071,17'd628,17'd1120,17'd53592,17'd18144,17'd52461,17'd18144,17'd796,17'd447,17'd38071,17'd38071,17'd5628,17'd18144,17'd53593,17'd18758,17'd53594,17'd53437,17'd53595,17'd53596,17'd53597,17'd53598,17'd53599,17'd53600
},
'{
17'd53228,17'd3592,17'd11609,17'd3429,17'd2936,17'd1416,17'd653,17'd27,17'd27,17'd285,17'd285,17'd467,17'd2937,17'd2937,17'd2937,17'd467,17'd7385,17'd7385,17'd7060,17'd7060,17'd4430,17'd4430,17'd4431,17'd4431,17'd6278,17'd6278,17'd11210,17'd3434,17'd5379,17'd5657,17'd5806,17'd5806,17'd4742,17'd51415,17'd4435,17'd33542,17'd24969,17'd48813,17'd23661,17'd27102,17'd53601,17'd5822,17'd53602,17'd53603,17'd19002,17'd15636,17'd20289,17'd20883,17'd53604,17'd13969,17'd14621,17'd12813,17'd15516,17'd12357,17'd14469,17'd12357,17'd22802,17'd19127,17'd22802,17'd15763,17'd11084,17'd11084,17'd13460,17'd14620,17'd14620,17'd12214,17'd10937,17'd13599,17'd14621,17'd14621,17'd13093,17'd12679,17'd13093,17'd13211,17'd13969,17'd22630,17'd20886,17'd28205,17'd17941,17'd17941,17'd18655,17'd16766,17'd16410,17'd17319,17'd16659,17'd15261,17'd16030,17'd33857,17'd53605,17'd53606,17'd53607,17'd53608,17'd53609,17'd3303,17'd3293,17'd4468,17'd53610,17'd53611,17'd53612,17'd42797,17'd42663,17'd53613,17'd53527,17'd53528,17'd53529,17'd53614,17'd51022,17'd50765,17'd50934,17'd43892,17'd48390,17'd53615,17'd41786,17'd48193,17'd48475,17'd53531,17'd52118,17'd49615,17'd27606,17'd27109,17'd26859,17'd53455,17'd53616,17'd53617,17'd53177,17'd10444,17'd53618,17'd15797,17'd53619,17'd52214,17'd53620,17'd10831,17'd11253,17'd53537,17'd53621,17'd53622,17'd17835,17'd16678,17'd11651,17'd11651,17'd24356,17'd24356,17'd12098,17'd23844,17'd53623,17'd53182,17'd53624,17'd53625,17'd53626,17'd53391,17'd17013,17'd53102,17'd15571,17'd14672,17'd14523,17'd18684,17'd12995,17'd13252,17'd17474,17'd17602,17'd17722,17'd21361,17'd21363,17'd21505,17'd23515,17'd25672,17'd29480,17'd31764,17'd33088,17'd51512,17'd53320,17'd53471,17'd53627,17'd53544,17'd53393,17'd53628,17'd53393,17'd53629,17'd53545,17'd53630,17'd34545,17'd31941,17'd32122,17'd30673,17'd33726,17'd24209,17'd52220,17'd19643,17'd24029,17'd11808,17'd14931,17'd14810,17'd12862,17'd14931,17'd10853,17'd18560,17'd19412,17'd11958,17'd12109,17'd15184,17'd15183,17'd14133,17'd53631,17'd9741,17'd9338,17'd15187,17'd9480,17'd19279,17'd22131,17'd11136,17'd9885,17'd20756,17'd10476,17'd14931,17'd23338,17'd19645,17'd13363,17'd13883,17'd11958,17'd12719,17'd12581,17'd11958,17'd13364,17'd13364,17'd12719,17'd13762,17'd48579,17'd50864,17'd19418,17'd23177,17'd11534,17'd7954,17'd53632,17'd36204,17'd53633,17'd11405,17'd12119,17'd16072,17'd22648,17'd46612,17'd9485,17'd15192,17'd53634,17'd53635,17'd17731,17'd53636,17'd53637,17'd22307,17'd53638,17'd130,17'd130,17'd132,17'd11683,17'd53639,17'd53640,17'd52741,17'd53641,17'd51552,17'd53642,17'd53643,17'd53644,17'd53645,17'd52255,17'd53646,17'd49582,17'd50736,17'd50272,17'd43011,17'd50660,17'd52000,17'd53647,17'd49788,17'd40507,17'd48899,17'd45609,17'd46094,17'd36127,17'd53648,17'd53412,17'd33654,17'd33654,17'd28134,17'd27885,17'd30279,17'd27761,17'd28371,17'd29979,17'd30131,17'd33489,17'd33489,17'd33489,17'd33489,17'd30280,17'd30280,17'd30736,17'd30736,17'd31505,17'd31506,17'd33489,17'd30736,17'd33322,17'd30738,17'd30884,17'd53338,17'd32354,17'd27885,17'd28134,17'd28134,17'd53339,17'd28855,17'd28854,17'd26276,17'd30279,17'd28134,17'd32355,17'd39910,17'd41109,17'd47729,17'd39272,17'd53649,17'd48909,17'd49682,17'd50568,17'd51741,17'd51920,17'd52675,17'd50736,17'd49485,17'd48359,17'd49472,17'd52818,17'd46102,17'd43285,17'd43550,17'd43694,17'd38406,17'd29688,17'd34137,17'd23217,17'd39131,17'd36288,17'd32830,17'd29686,17'd23732,17'd28367,17'd34283,17'd32007,17'd29688,17'd23733,17'd23387,17'd32351,17'd22679,17'd36870,17'd23574,17'd30727,17'd33161,17'd46860,17'd52680,17'd53650,17'd52886,17'd53651,17'd53652,17'd34880,17'd42305,17'd53653,17'd53654,17'd53568,17'd53655,17'd53656,17'd53657,17'd53658,17'd53421,17'd23081,17'd53659,17'd43725,17'd22920,17'd53660,17'd53661,17'd29590,17'd7166,17'd5913,17'd5609,17'd4992,17'd4188,17'd40079,17'd5477,17'd4838,17'd6067,17'd4686,17'd5330,17'd27935,17'd32073,17'd32074,17'd32074,17'd32074,17'd29740,17'd7499,17'd32073,17'd6390,17'd6219,17'd9091,17'd32073,17'd32073,17'd32073,17'd32073,17'd9091,17'd9091,17'd9091,17'd27696,17'd27696,17'd7668,17'd7499,17'd9091,17'd9091,17'd9091,17'd7499,17'd6220,17'd5614,17'd5160,17'd31401,17'd28418,17'd5335,17'd5164,17'd5338,17'd5013,17'd53662,17'd49498,17'd53663,17'd53664,17'd53665,17'd47083,17'd53666,17'd42472,17'd53667,17'd53668,17'd53669,17'd53513,17'd53670,17'd2077,17'd53671,17'd53672,17'd3058,17'd45655,17'd51581,17'd4552,17'd5626,17'd53673,17'd41159,17'd5495,17'd38857,17'd5496,17'd38857,17'd53068,17'd53068,17'd4399,17'd52918,17'd4398,17'd38071,17'd628,17'd1944,17'd53592,17'd3071,17'd53674,17'd1943,17'd628,17'd1264,17'd53068,17'd4399,17'd4228,17'd53675,17'd36322,17'd52773,17'd53676,17'd53437,17'd53677,17'd53596,17'd53597,17'd53678,17'd53679,17'd53600
},
'{
17'd52704,17'd15496,17'd11609,17'd3429,17'd2596,17'd1416,17'd28,17'd980,17'd27,17'd27,17'd285,17'd467,17'd467,17'd467,17'd467,17'd2937,17'd1833,17'd286,17'd286,17'd27,17'd4248,17'd4248,17'd18037,17'd4431,17'd6278,17'd3910,17'd3434,17'd3434,17'd5658,17'd5658,17'd5210,17'd5054,17'd4742,17'd5057,17'd4433,17'd3917,17'd3601,17'd12932,17'd28077,17'd27102,17'd53680,17'd39793,17'd53681,17'd13445,17'd53682,17'd13082,17'd17931,17'd22459,17'd53683,17'd28554,17'd12530,17'd35352,17'd15516,17'd22802,17'd22802,17'd15763,17'd12679,17'd12527,17'd12679,17'd22802,17'd11084,17'd50503,17'd14216,17'd14620,17'd52468,17'd12214,17'd10937,17'd13092,17'd12955,17'd14621,17'd12065,17'd34938,17'd13093,17'd14621,17'd12361,17'd16658,17'd18884,17'd19006,17'd11362,17'd18412,17'd11915,17'd18174,17'd16410,17'd16289,17'd24348,17'd15009,17'd16031,17'd48387,17'd53684,17'd50094,17'd53685,17'd53686,17'd53687,17'd2975,17'd3958,17'd4930,17'd2658,17'd53688,17'd53689,17'd53690,17'd42663,17'd53691,17'd53692,17'd53693,17'd53694,17'd53695,17'd51022,17'd50765,17'd51105,17'd50848,17'd53173,17'd53696,17'd42669,17'd48193,17'd38895,17'd7435,17'd53697,17'd53380,17'd30513,17'd27331,17'd9594,17'd24982,17'd20302,17'd53312,17'd53313,17'd53698,17'd15796,17'd15927,17'd53699,17'd19403,17'd15419,17'd53700,17'd10832,17'd53384,17'd53701,17'd53702,17'd53703,17'd53704,17'd11651,17'd14514,17'd14514,17'd24356,17'd12403,17'd22294,17'd53705,17'd53540,17'd53387,17'd53541,17'd53706,17'd53707,17'd17476,17'd53708,17'd17013,17'd16686,17'd16799,17'd13512,17'd18684,17'd13518,17'd15433,17'd17602,17'd17722,17'd21361,17'd22992,17'd24362,17'd23168,17'd23856,17'd29778,17'd28686,17'd32437,17'd50863,17'd52133,17'd52870,17'd53471,17'd53471,17'd53322,17'd53628,17'd53709,17'd53544,17'd52868,17'd52400,17'd50111,17'd34203,17'd31765,17'd29779,17'd29476,17'd25925,17'd21362,17'd19921,17'd13516,17'd10989,17'd14931,17'd14931,17'd14673,17'd14673,17'd10737,17'd18682,17'd18330,17'd12260,17'd12580,17'd12253,17'd18450,17'd13366,17'd15182,17'd22296,17'd9472,17'd9341,17'd16549,17'd16549,17'd24998,17'd9619,17'd9741,17'd21503,17'd10991,17'd51273,17'd12720,17'd13885,17'd20313,17'd11806,17'd11806,17'd13135,17'd12996,17'd11961,17'd13363,17'd13135,17'd12996,17'd11666,17'd15181,17'd47298,17'd8732,17'd35512,17'd7955,17'd15439,17'd12590,17'd53710,17'd23687,17'd23864,17'd23864,17'd8251,17'd19418,17'd17351,17'd7789,17'd7790,17'd24714,17'd8891,17'd53711,17'd21371,17'd53712,17'd53713,17'd7980,17'd134,17'd1481,17'd133,17'd52157,17'd53714,17'd52963,17'd53715,17'd53716,17'd50733,17'd50362,17'd53486,17'd50462,17'd50821,17'd49388,17'd48909,17'd50468,17'd50272,17'd50273,17'd43011,17'd43146,17'd52000,17'd50574,17'd49484,17'd40673,17'd44223,17'd48035,17'd32005,17'd27885,17'd32192,17'd33164,17'd33654,17'd33654,17'd32192,17'd26522,17'd28854,17'd28133,17'd29537,17'd29978,17'd30280,17'd33489,17'd33323,17'd33489,17'd33489,17'd30280,17'd30736,17'd31505,17'd31505,17'd31506,17'd31506,17'd30280,17'd31036,17'd32019,17'd28857,17'd53717,17'd33164,17'd27885,17'd31354,17'd31503,17'd29379,17'd37513,17'd33952,17'd33001,17'd33001,17'd32354,17'd28373,17'd28373,17'd35854,17'd43547,17'd53718,17'd46104,17'd48153,17'd49288,17'd49683,17'd51157,17'd51741,17'd52169,17'd52000,17'd49985,17'd49182,17'd48142,17'd53719,17'd48614,17'd48258,17'd46426,17'd43549,17'd43157,17'd53720,17'd24087,17'd23387,17'd29973,17'd41419,17'd36288,17'd23217,17'd29376,17'd28852,17'd29240,17'd24898,17'd25031,17'd32659,17'd23918,17'd23388,17'd23218,17'd22678,17'd23741,17'd53721,17'd22009,17'd33797,17'd51468,17'd53722,17'd53723,17'd53724,17'd51067,17'd21530,17'd35154,17'd42747,17'd51394,17'd51563,17'd46860,17'd22340,17'd53725,17'd53726,17'd53727,17'd53728,17'd19961,17'd53729,17'd53730,17'd53731,17'd29883,17'd25877,17'd11013,17'd7327,17'd6212,17'd5326,17'd6381,17'd33365,17'd43584,17'd5754,17'd4837,17'd4683,17'd5002,17'd25627,17'd31717,17'd7499,17'd32074,17'd29740,17'd27696,17'd32074,17'd32073,17'd9091,17'd9091,17'd7499,17'd9091,17'd9091,17'd32074,17'd29740,17'd29740,17'd29740,17'd29740,17'd29740,17'd29740,17'd27696,17'd8780,17'd7499,17'd36586,17'd36586,17'd9091,17'd7668,17'd6219,17'd5614,17'd25627,17'd31552,17'd30180,17'd5335,17'd5165,17'd53732,17'd53733,17'd53427,17'd38706,17'd53734,17'd53735,17'd53736,17'd37298,17'd53737,17'd53738,17'd53739,17'd53740,17'd53741,17'd53742,17'd53670,17'd2077,17'd53743,17'd41769,17'd53744,17'd52916,17'd3380,17'd3703,17'd4054,17'd3870,17'd39179,17'd5495,17'd38857,17'd4399,17'd53068,17'd53068,17'd53068,17'd4399,17'd4399,17'd4398,17'd4059,17'd1120,17'd5775,17'd1943,17'd53674,17'd6867,17'd235,17'd959,17'd447,17'd4398,17'd4398,17'd5628,17'd18144,17'd53745,17'd53746,17'd53594,17'd53747,17'd53595,17'd53748,17'd53749,17'd53750,17'd53751,17'd53752
},
'{
17'd52704,17'd3592,17'd11609,17'd3429,17'd2597,17'd1414,17'd288,17'd652,17'd27,17'd27,17'd285,17'd467,17'd467,17'd467,17'd467,17'd467,17'd1833,17'd286,17'd286,17'd286,17'd4248,17'd4248,17'd18037,17'd4431,17'd6278,17'd3910,17'd3434,17'd3434,17'd5658,17'd5658,17'd5210,17'd4739,17'd13819,17'd50757,17'd2608,17'd3917,17'd3603,17'd12659,17'd27829,17'd15749,17'd53753,17'd4752,17'd5987,17'd53754,17'd13080,17'd21805,17'd18290,17'd53755,17'd45069,17'd28438,17'd13969,17'd34015,17'd15516,17'd22802,17'd22802,17'd15763,17'd12679,17'd12527,17'd12679,17'd12527,17'd12062,17'd50503,17'd14216,17'd14620,17'd52468,17'd12214,17'd10937,17'd12954,17'd13211,17'd14621,17'd12065,17'd34938,17'd13093,17'd14621,17'd12361,17'd16658,17'd18884,17'd18884,17'd11362,17'd18412,17'd11915,17'd18174,17'd16410,17'd16289,17'd24348,17'd15770,17'd14624,17'd48387,17'd53605,17'd53301,17'd53756,17'd53757,17'd53758,17'd3131,17'd3303,17'd2979,17'd2471,17'd5265,17'd53759,17'd53760,17'd53691,17'd6155,17'd6012,17'd53693,17'd53694,17'd53695,17'd50193,17'd50847,17'd50765,17'd41501,17'd53761,17'd53762,17'd42669,17'd53763,17'd47674,17'd48935,17'd53697,17'd8393,17'd51423,17'd27606,17'd53532,17'd24982,17'd20302,17'd53616,17'd53617,17'd53764,17'd53765,17'd10827,17'd53766,17'd53767,17'd53768,17'd53769,17'd53770,17'd53771,17'd53702,17'd53772,17'd53773,17'd25402,17'd11941,17'd14514,17'd14514,17'd24356,17'd12407,17'd21497,17'd24697,17'd53386,17'd53182,17'd53774,17'd53775,17'd53776,17'd17476,17'd53708,17'd17724,17'd16560,17'd13134,17'd18807,17'd18684,17'd13760,17'd15570,17'd17602,17'd17722,17'd21361,17'd22992,17'd24362,17'd22819,17'd23512,17'd29778,17'd29066,17'd47403,17'd31589,17'd52867,17'd52800,17'd53321,17'd53321,17'd53322,17'd53709,17'd53777,17'd53709,17'd53321,17'd53473,17'd35239,17'd33875,17'd30834,17'd31587,17'd30673,17'd26872,17'd24209,17'd14258,17'd18444,17'd13516,17'd11274,17'd11274,17'd14673,17'd14673,17'd10736,17'd10737,17'd18560,17'd12260,17'd16321,17'd12253,17'd16324,17'd14130,17'd13764,17'd10604,17'd15300,17'd17012,17'd9619,17'd19279,17'd33083,17'd15187,17'd10742,17'd10992,17'd11134,17'd10477,17'd10605,17'd15182,17'd11666,17'd11963,17'd11963,17'd12996,17'd12422,17'd12996,17'd11806,17'd12996,17'd11806,17'd11520,17'd52726,17'd28577,17'd23861,17'd8581,17'd8735,17'd16567,17'd24869,17'd14390,17'd12726,17'd17850,17'd24215,17'd8250,17'd18203,17'd7786,17'd14681,17'd22135,17'd9891,17'd8427,17'd17131,17'd16211,17'd53778,17'd53779,17'd12275,17'd131,17'd542,17'd16090,17'd53780,17'd20929,17'd21389,17'd47835,17'd53781,17'd53405,17'd52888,17'd52967,17'd51736,17'd47436,17'd48792,17'd50467,17'd50268,17'd50661,17'd50273,17'd50273,17'd50661,17'd50476,17'd49891,17'd43147,17'd43831,17'd44593,17'd39740,17'd39437,17'd33319,17'd33164,17'd33319,17'd28134,17'd28134,17'd32192,17'd28981,17'd28856,17'd29380,17'd29536,17'd29978,17'd30280,17'd33323,17'd33323,17'd33323,17'd33489,17'd30280,17'd30736,17'd31506,17'd31506,17'd31506,17'd30736,17'd31036,17'd30738,17'd29831,17'd29380,17'd33654,17'd32354,17'd27642,17'd31353,17'd31352,17'd28727,17'd28979,17'd28980,17'd33952,17'd33001,17'd32192,17'd28373,17'd40367,17'd40961,17'd41416,17'd44472,17'd48901,17'd48535,17'd50822,17'd50365,17'd51830,17'd52671,17'd52675,17'd50272,17'd49693,17'd45742,17'd47825,17'd53782,17'd50152,17'd42884,17'd43835,17'd43694,17'd42302,17'd34276,17'd23918,17'd32191,17'd36426,17'd36288,17'd32830,17'd30128,17'd23733,17'd29100,17'd27763,17'd24898,17'd32007,17'd23916,17'd23565,17'd23388,17'd23218,17'd22678,17'd53564,17'd35292,17'd31832,17'd35154,17'd53783,17'd53784,17'd53723,17'd53785,17'd46775,17'd21531,17'd42747,17'd51479,17'd53786,17'd47069,17'd53787,17'd53788,17'd53789,17'd53790,17'd53791,17'd35743,17'd23434,17'd53792,17'd53793,17'd53731,17'd30028,17'd25221,17'd10627,17'd7327,17'd23799,17'd7008,17'd24148,17'd33365,17'd5477,17'd4523,17'd4682,17'd32552,17'd5002,17'd30638,17'd6554,17'd7499,17'd34658,17'd29740,17'd27696,17'd32074,17'd32073,17'd9091,17'd7499,17'd7499,17'd9091,17'd9091,17'd29740,17'd29740,17'd29740,17'd29740,17'd29740,17'd29740,17'd29740,17'd9933,17'd8780,17'd9091,17'd36586,17'd36586,17'd9091,17'd6391,17'd5615,17'd5762,17'd5005,17'd31716,17'd30637,17'd5166,17'd53794,17'd5617,17'd53579,17'd4372,17'd39617,17'd53795,17'd53796,17'd3363,17'd46695,17'd45063,17'd53797,17'd53798,17'd53799,17'd53800,17'd53801,17'd53802,17'd53803,17'd53671,17'd38713,17'd53744,17'd52916,17'd41479,17'd41480,17'd5626,17'd51857,17'd39179,17'd18142,17'd38857,17'd53068,17'd53068,17'd53068,17'd53068,17'd4399,17'd4399,17'd4398,17'd4059,17'd1944,17'd1944,17'd18144,17'd53674,17'd6867,17'd1943,17'd796,17'd795,17'd4399,17'd4399,17'd4228,17'd2557,17'd36322,17'd53746,17'd53594,17'd53747,17'd53595,17'd53748,17'd53749,17'd53678,17'd53804,17'd53752
},
'{
17'd52704,17'd3592,17'd10925,17'd3429,17'd2597,17'd22965,17'd652,17'd652,17'd27,17'd27,17'd286,17'd1833,17'd285,17'd467,17'd467,17'd467,17'd467,17'd285,17'd286,17'd286,17'd4248,17'd4248,17'd4431,17'd4431,17'd10269,17'd3910,17'd3434,17'd4249,17'd5210,17'd5210,17'd25790,17'd25790,17'd13819,17'd13820,17'd37171,17'd1707,17'd33851,17'd3110,17'd53805,17'd28920,17'd53806,17'd32888,17'd14877,17'd53807,17'd19619,17'd12942,17'd16276,17'd53808,17'd29621,17'd19892,17'd22630,17'd23154,17'd15516,17'd12527,17'd22802,17'd22802,17'd12527,17'd12527,17'd13093,17'd12527,17'd12062,17'd50503,17'd14216,17'd14620,17'd14620,17'd12214,17'd12062,17'd13092,17'd12955,17'd14621,17'd12065,17'd11626,17'd34938,17'd13094,17'd13969,17'd22630,17'd18884,17'd18884,17'd12681,17'd18412,17'd11915,17'd18174,17'd17318,17'd16289,17'd24348,17'd17322,17'd15009,17'd15641,17'd53809,17'd50094,17'd53810,17'd53811,17'd53812,17'd53813,17'd3478,17'd3791,17'd53814,17'd4617,17'd53815,17'd53816,17'd53817,17'd53374,17'd53818,17'd53819,17'd53820,17'd53821,17'd50193,17'd50394,17'd50847,17'd50765,17'd53822,17'd53823,17'd53824,17'd41786,17'd40278,17'd48475,17'd53825,17'd52118,17'd51502,17'd28929,17'd52210,17'd26990,17'd23673,17'd53616,17'd18071,17'd53617,17'd10578,17'd10710,17'd53826,17'd53382,17'd18674,17'd16545,17'd53827,17'd53828,17'd53829,17'd53830,17'd53831,17'd24698,17'd11792,17'd11942,17'd14514,17'd24356,17'd12402,17'd18800,17'd21976,17'd25271,17'd53832,17'd53387,17'd53468,17'd53626,17'd53391,17'd53708,17'd17724,17'd17013,17'd17015,17'd44647,17'd14523,17'd14809,17'd21506,17'd50779,17'd12106,17'd17722,17'd18198,17'd14130,17'd21671,17'd23512,17'd27004,17'd30830,17'd40133,17'd32283,17'd51118,17'd52867,17'd52799,17'd53321,17'd53321,17'd53393,17'd53833,17'd53833,17'd53393,17'd52868,17'd50952,17'd31590,17'd33568,17'd30221,17'd29330,17'd28345,17'd24856,17'd29781,17'd20609,17'd16326,17'd11964,17'd13516,17'd11964,17'd14262,17'd10736,17'd10736,17'd10989,17'd13362,17'd13883,17'd15184,17'd12253,17'd15184,17'd13363,17'd11520,17'd11133,17'd21503,17'd9741,17'd22131,17'd33083,17'd15569,17'd17011,17'd9885,17'd16796,17'd10991,17'd13001,17'd12720,17'd29331,17'd11520,17'd11667,17'd11667,17'd13362,17'd13362,17'd12996,17'd11806,17'd13253,17'd11520,17'd20908,17'd14666,17'd17716,17'd25147,17'd53834,17'd53835,17'd15438,17'd17852,17'd25004,17'd15440,17'd16446,17'd53836,17'd15435,17'd17484,17'd15302,17'd14938,17'd24868,17'd25293,17'd12868,17'd9893,17'd18093,17'd53837,17'd52959,17'd17363,17'd889,17'd20464,17'd53838,17'd53839,17'd53840,17'd22007,17'd40960,17'd33802,17'd52967,17'd53841,17'd51154,17'd47044,17'd47641,17'd51916,17'd50272,17'd50660,17'd50739,17'd50272,17'd50739,17'd50370,17'd50822,17'd48155,17'd44936,17'd42298,17'd36542,17'd27642,17'd33319,17'd33319,17'd30279,17'd32832,17'd28854,17'd28981,17'd28856,17'd31196,17'd28857,17'd29831,17'd29978,17'd30131,17'd33323,17'd33323,17'd30131,17'd30131,17'd30280,17'd30280,17'd30280,17'd30736,17'd30280,17'd30280,17'd32019,17'd36132,17'd32017,17'd32354,17'd32832,17'd31503,17'd29245,17'd28486,17'd27027,17'd27027,17'd27027,17'd28979,17'd37513,17'd33001,17'd32192,17'd32832,17'd35291,17'd41582,17'd53842,17'd48990,17'd46956,17'd48264,17'd49692,17'd50272,17'd51741,17'd52671,17'd53843,17'd49986,17'd52170,17'd53844,17'd47443,17'd53845,17'd53846,17'd43017,17'd43694,17'd44105,17'd51392,17'd35159,17'd23566,17'd23217,17'd23740,17'd33316,17'd29973,17'd29530,17'd24086,17'd34884,17'd34283,17'd25030,17'd25032,17'd24249,17'd29099,17'd30128,17'd36986,17'd22332,17'd22160,17'd49096,17'd35295,17'd51479,17'd53847,17'd53848,17'd53849,17'd53850,17'd51726,17'd21530,17'd52985,17'd51562,17'd47163,17'd53851,17'd53852,17'd53853,17'd53854,17'd53855,17'd53856,17'd53857,17'd53858,17'd22402,17'd53859,17'd22752,17'd23969,17'd26326,17'd10198,17'd7327,17'd23799,17'd6702,17'd7005,17'd53278,17'd4523,17'd4837,17'd4840,17'd4845,17'd25627,17'd28185,17'd6219,17'd9091,17'd34658,17'd29740,17'd7499,17'd9091,17'd9091,17'd9091,17'd7499,17'd7499,17'd29740,17'd29740,17'd29740,17'd29740,17'd29740,17'd29740,17'd27696,17'd27696,17'd29740,17'd9933,17'd7668,17'd9091,17'd6554,17'd6390,17'd6219,17'd6220,17'd5614,17'd5336,17'd4842,17'd28536,17'd5009,17'd5166,17'd51930,17'd53353,17'd53662,17'd53860,17'd52185,17'd38063,17'd37703,17'd53861,17'd53862,17'd53863,17'd53864,17'd53865,17'd53866,17'd53867,17'd53868,17'd53869,17'd53803,17'd40858,17'd51182,17'd53870,17'd52916,17'd3217,17'd4053,17'd4394,17'd40099,17'd4710,17'd18035,17'd4398,17'd38071,17'd38071,17'd53068,17'd4399,17'd4398,17'd38071,17'd38071,17'd38071,17'd5775,17'd1120,17'd236,17'd237,17'd52462,17'd451,17'd234,17'd2587,17'd4398,17'd4398,17'd5628,17'd2557,17'd53152,17'd35206,17'd53594,17'd53747,17'd53871,17'd53872,17'd53873,17'd53750,17'd53751,17'd53752
},
'{
17'd5511,17'd3592,17'd10925,17'd3429,17'd2597,17'd2257,17'd29,17'd652,17'd27,17'd27,17'd286,17'd286,17'd285,17'd285,17'd467,17'd467,17'd467,17'd285,17'd286,17'd286,17'd4430,17'd4430,17'd4431,17'd4431,17'd10269,17'd3910,17'd3434,17'd3104,17'd4250,17'd4739,17'd25790,17'd3106,17'd53874,17'd2432,17'd39630,17'd1706,17'd3917,17'd3440,17'd2797,17'd39632,17'd53875,17'd53876,17'd53877,17'd53878,17'd21034,17'd12941,17'd53879,17'd21647,17'd46482,17'd19892,17'd28554,17'd13094,17'd12813,17'd12527,17'd22802,17'd22802,17'd12527,17'd13093,17'd12955,17'd13093,17'd12677,17'd12062,17'd13461,17'd13460,17'd14620,17'd12355,17'd12062,17'd12954,17'd14621,17'd14764,17'd12065,17'd11626,17'd34938,17'd13094,17'd13969,17'd28554,17'd19006,17'd18884,17'd12532,17'd18412,17'd11915,17'd18174,17'd17318,17'd16519,17'd15524,17'd16769,17'd15009,17'd16030,17'd53809,17'd53301,17'd53880,17'd53811,17'd53812,17'd53881,17'd3478,17'd3958,17'd4773,17'd2658,17'd5699,17'd53882,17'd53883,17'd53884,17'd53885,17'd53886,17'd53887,17'd53888,17'd53889,17'd51022,17'd50847,17'd41177,17'd41648,17'd53173,17'd53615,17'd42669,17'd50195,17'd53890,17'd35080,17'd52118,17'd51502,17'd30513,17'd51263,17'd52120,17'd23673,17'd53891,17'd53616,17'd18071,17'd53764,17'd17112,17'd10827,17'd53459,17'd53892,17'd53893,17'd53894,17'd53895,17'd15036,17'd15036,17'd25920,17'd24698,17'd11791,17'd11941,17'd11942,17'd12245,17'd12989,17'd12989,17'd12244,17'd53896,17'd24021,17'd53897,17'd53898,17'd53899,17'd53900,17'd17476,17'd17013,17'd17013,17'd17014,17'd16686,17'd14672,17'd13643,17'd13518,17'd15685,17'd12106,17'd18198,17'd18198,17'd21671,17'd22819,17'd23512,17'd25672,17'd30524,17'd53901,17'd39211,17'd31442,17'd51272,17'd53187,17'd52799,17'd53321,17'd53393,17'd53709,17'd53833,17'd53628,17'd52799,17'd51881,17'd50951,17'd31590,17'd33568,17'd31439,17'd29779,17'd28227,17'd23512,17'd20608,17'd18443,17'd19158,17'd13762,17'd11964,17'd11964,17'd14262,17'd14262,17'd10989,17'd11964,17'd13520,17'd13761,17'd12109,17'd12414,17'd13882,17'd12861,17'd14931,17'd10328,17'd9473,17'd22131,17'd15298,17'd16549,17'd15048,17'd9741,17'd18916,17'd11134,17'd14666,17'd10605,17'd12720,17'd11519,17'd11666,17'd13764,17'd11667,17'd12262,17'd16204,17'd13253,17'd11395,17'd11666,17'd11395,17'd17121,17'd14928,17'd8726,17'd12589,17'd10610,17'd13378,17'd14816,17'd9891,17'd8257,17'd16919,17'd16803,17'd53902,17'd25286,17'd15302,17'd7621,17'd11969,17'd11814,17'd7958,17'd15195,17'd18336,17'd53903,17'd53904,17'd11152,17'd888,17'd23537,17'd53905,17'd21228,17'd34880,17'd22500,17'd30431,17'd38406,17'd53906,17'd50461,17'd52163,17'd53907,17'd48793,17'd49980,17'd50739,17'd43143,17'd50273,17'd50736,17'd50370,17'd49984,17'd48264,17'd45870,17'd44698,17'd42890,17'd31352,17'd30279,17'd32354,17'd32354,17'd27885,17'd27885,17'd28854,17'd29104,17'd31196,17'd30884,17'd29690,17'd29979,17'd29978,17'd29978,17'd30131,17'd33323,17'd30131,17'd30131,17'd30131,17'd30131,17'd30280,17'd30280,17'd30280,17'd30130,17'd36132,17'd28372,17'd32354,17'd27885,17'd31503,17'd28727,17'd28486,17'd26902,17'd27259,17'd28725,17'd26902,17'd26901,17'd37513,17'd33319,17'd32354,17'd32356,17'd34274,17'd43844,17'd53908,17'd45987,17'd53909,17'd43419,17'd50271,17'd51163,17'd51741,17'd53843,17'd51995,17'd49582,17'd45742,17'd53910,17'd51739,17'd53911,17'd48037,17'd43285,17'd43976,17'd53332,17'd33802,17'd24087,17'd30128,17'd29973,17'd32514,17'd32514,17'd29828,17'd29099,17'd23731,17'd28008,17'd24897,17'd25030,17'd25032,17'd34467,17'd34137,17'd30128,17'd32827,17'd22333,17'd35292,17'd21848,17'd33946,17'd51377,17'd53912,17'd53913,17'd21540,17'd53914,17'd21839,17'd21529,17'd51562,17'd53786,17'd53915,17'd53916,17'd53917,17'd53918,17'd53919,17'd53920,17'd53921,17'd53922,17'd43178,17'd53923,17'd53924,17'd23267,17'd24303,17'd53925,17'd7824,17'd23799,17'd25082,17'd7006,17'd53926,17'd6839,17'd5322,17'd6067,17'd4686,17'd5329,17'd31553,17'd31717,17'd7499,17'd9091,17'd34658,17'd32074,17'd9091,17'd9091,17'd9091,17'd7499,17'd7668,17'd7499,17'd29740,17'd29740,17'd29740,17'd29740,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd9933,17'd7668,17'd32073,17'd31717,17'd6390,17'd6219,17'd5615,17'd5336,17'd5335,17'd28536,17'd28418,17'd5163,17'd5163,17'd5338,17'd53353,17'd53927,17'd4201,17'd53928,17'd53929,17'd53930,17'd53931,17'd53932,17'd42327,17'd53933,17'd53934,17'd53935,17'd53936,17'd53937,17'd53938,17'd53939,17'd53940,17'd2726,17'd53870,17'd52916,17'd3217,17'd4053,17'd4394,17'd3871,17'd4710,17'd5936,17'd38071,17'd4059,17'd4059,17'd53068,17'd4399,17'd38071,17'd38071,17'd4059,17'd4398,17'd5775,17'd796,17'd237,17'd237,17'd52462,17'd235,17'd628,17'd795,17'd4399,17'd4399,17'd4228,17'd2557,17'd53152,17'd35206,17'd53594,17'd53941,17'd53942,17'd53872,17'd53873,17'd53678,17'd53804,17'd53752
},
'{
17'd15877,17'd3901,17'd10925,17'd3429,17'd2597,17'd22965,17'd652,17'd652,17'd27,17'd27,17'd286,17'd286,17'd285,17'd285,17'd285,17'd467,17'd467,17'd285,17'd286,17'd286,17'd4430,17'd4430,17'd4431,17'd4091,17'd6278,17'd3910,17'd3434,17'd3104,17'd4251,17'd2604,17'd4739,17'd2945,17'd50679,17'd2432,17'd39630,17'd1706,17'd3917,17'd3440,17'd2797,17'd53943,17'd53944,17'd53945,17'd5396,17'd53946,17'd13824,17'd19002,17'd18403,17'd21647,17'd53947,17'd53948,17'd53949,17'd12362,17'd12813,17'd12527,17'd15763,17'd22802,17'd12527,17'd13093,17'd12955,17'd13093,17'd12678,17'd12062,17'd14344,17'd13460,17'd13460,17'd12355,17'd12677,17'd12954,17'd14621,17'd12530,17'd12814,17'd12065,17'd34938,17'd13094,17'd13969,17'd28554,17'd20292,17'd29048,17'd12532,17'd12681,17'd17941,17'd18174,17'd21185,17'd19011,17'd18776,17'd16769,17'd15009,17'd16167,17'd53809,17'd50094,17'd53950,17'd53951,17'd53952,17'd53953,17'd53954,17'd3790,17'd2650,17'd2470,17'd53610,17'd53955,17'd53956,17'd53884,17'd53957,17'd53958,17'd53959,17'd53960,17'd53961,17'd50193,17'd50847,17'd41177,17'd51023,17'd53822,17'd53453,17'd53962,17'd45199,17'd48826,17'd53454,17'd53963,17'd53380,17'd49615,17'd51342,17'd52210,17'd53964,17'd20302,17'd53616,17'd53312,17'd53617,17'd10578,17'd10710,17'd53965,17'd53966,17'd53967,17'd13871,17'd14915,17'd53968,17'd15036,17'd53969,17'd53970,17'd24851,17'd11940,17'd53971,17'd53971,17'd17226,17'd12711,17'd19775,17'd53972,17'd53973,17'd53974,17'd13509,17'd53975,17'd53976,17'd45933,17'd17476,17'd17476,17'd17013,17'd17014,17'd16686,17'd32138,17'd14809,17'd13252,17'd12106,17'd12106,17'd20314,17'd21671,17'd23168,17'd23512,17'd27347,17'd27346,17'd30218,17'd28686,17'd31941,17'd36213,17'd53977,17'd53187,17'd52799,17'd53393,17'd53472,17'd53709,17'd53628,17'd53322,17'd52868,17'd53473,17'd35239,17'd34037,17'd31761,17'd31285,17'd30673,17'd24856,17'd23170,17'd20608,17'd16442,17'd15185,17'd16326,17'd13516,17'd11397,17'd14673,17'd11274,17'd10989,17'd13762,17'd12861,17'd12419,17'd12577,17'd12577,17'd13363,17'd11520,17'd10474,17'd10856,17'd18196,17'd22131,17'd9619,17'd15048,17'd12116,17'd18441,17'd16796,17'd14518,17'd11132,17'd10990,17'd14931,17'd16068,17'd16064,17'd11667,17'd11964,17'd13516,17'd11807,17'd14262,17'd11395,17'd14262,17'd12720,17'd10479,17'd9041,17'd25411,17'd13891,17'd22299,17'd13894,17'd53978,17'd18086,17'd14680,17'd23345,17'd21988,17'd16334,17'd53979,17'd14679,17'd18205,17'd53980,17'd53981,17'd10031,17'd22140,17'd14686,17'd53982,17'd53983,17'd889,17'd53984,17'd53985,17'd21538,17'd48274,17'd31195,17'd28368,17'd38282,17'd48895,17'd53986,17'd49374,17'd47538,17'd49684,17'd50072,17'd43143,17'd43143,17'd50476,17'd50365,17'd49984,17'd48995,17'd53987,17'd41415,17'd45484,17'd36127,17'd27642,17'd31354,17'd27885,17'd28134,17'd28134,17'd33319,17'd28854,17'd29247,17'd28857,17'd29979,17'd49790,17'd49790,17'd29978,17'd29978,17'd30131,17'd30131,17'd30131,17'd30131,17'd30131,17'd30131,17'd30131,17'd30131,17'd30738,17'd30130,17'd32018,17'd33654,17'd28258,17'd31354,17'd31035,17'd26782,17'd26902,17'd27259,17'd27640,17'd27259,17'd26902,17'd28486,17'd29246,17'd27885,17'd30279,17'd36264,17'd43560,17'd45481,17'd45750,17'd43420,17'd49082,17'd49093,17'd50574,17'd51741,17'd51741,17'd53197,17'd50468,17'd49183,17'd53988,17'd53989,17'd51555,17'd53990,17'd53563,17'd46659,17'd53486,17'd51392,17'd29688,17'd23918,17'd23215,17'd30425,17'd32514,17'd32504,17'd23386,17'd23733,17'd30879,17'd34884,17'd25032,17'd25180,17'd25032,17'd24415,17'd34137,17'd32351,17'd22331,17'd22160,17'd35153,17'd51749,17'd52172,17'd47749,17'd53991,17'd53992,17'd51641,17'd51468,17'd22153,17'd53993,17'd51726,17'd53915,17'd53994,17'd53995,17'd53996,17'd53997,17'd53998,17'd53999,17'd54000,17'd20360,17'd54001,17'd22402,17'd28416,17'd54002,17'd24642,17'd11294,17'd23975,17'd5608,17'd24647,17'd53506,17'd7004,17'd4677,17'd5756,17'd4995,17'd4687,17'd5329,17'd31553,17'd6554,17'd7499,17'd32073,17'd9091,17'd9091,17'd6219,17'd6390,17'd9091,17'd7668,17'd27696,17'd29740,17'd29740,17'd29740,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd9933,17'd7499,17'd36586,17'd31717,17'd6554,17'd5615,17'd5614,17'd5335,17'd25627,17'd31716,17'd28418,17'd5166,17'd5163,17'd5169,17'd53733,17'd54003,17'd54004,17'd51491,17'd38708,17'd54005,17'd54006,17'd54007,17'd54008,17'd54009,17'd54010,17'd54011,17'd54012,17'd54013,17'd53802,17'd2077,17'd40713,17'd41769,17'd53870,17'd52916,17'd51252,17'd40562,17'd5494,17'd54014,17'd54015,17'd5936,17'd38071,17'd4059,17'd38071,17'd38071,17'd38071,17'd38071,17'd4059,17'd4059,17'd2558,17'd1944,17'd1121,17'd797,17'd237,17'd630,17'd448,17'd628,17'd1120,17'd4398,17'd4399,17'd6239,17'd2557,17'd53152,17'd35206,17'd53594,17'd53747,17'd53871,17'd53872,17'd53873,17'd53598,17'd53751,17'd53752
},
'{
17'd15877,17'd3901,17'd10925,17'd3429,17'd2597,17'd2425,17'd29,17'd652,17'd980,17'd27,17'd286,17'd286,17'd285,17'd285,17'd285,17'd467,17'd467,17'd285,17'd286,17'd286,17'd4430,17'd4430,17'd4431,17'd4091,17'd6278,17'd3756,17'd3435,17'd2944,17'd2604,17'd2946,17'd2946,17'd1975,17'd2432,17'd2433,17'd44851,17'd1705,17'd1978,17'd3600,17'd13072,17'd29759,17'd15881,17'd2802,17'd20876,17'd20417,17'd54016,17'd13825,17'd54017,17'd54018,17'd54019,17'd53948,17'd32102,17'd13969,17'd12065,17'd12527,17'd15763,17'd12527,17'd12813,17'd13093,17'd14621,17'd13211,17'd12812,17'd12357,17'd14344,17'd13460,17'd13460,17'd12355,17'd12677,17'd12813,17'd12218,17'd12530,17'd12814,17'd12065,17'd11626,17'd13094,17'd12361,17'd22630,17'd20292,17'd28667,17'd12532,17'd11362,17'd11915,17'd17205,17'd19255,17'd27833,17'd18776,17'd15524,17'd16032,17'd47673,17'd53809,17'd53301,17'd54020,17'd54021,17'd53686,17'd53953,17'd53954,17'd3478,17'd54022,17'd54023,17'd54024,17'd54025,17'd54026,17'd53816,17'd53885,17'd54027,17'd54028,17'd54029,17'd46493,17'd50193,17'd53306,17'd54030,17'd54031,17'd54032,17'd54033,17'd53824,17'd41786,17'd48933,17'd50398,17'd52555,17'd49418,17'd49615,17'd28929,17'd51263,17'd54034,17'd23673,17'd25917,17'd53616,17'd18071,17'd53764,17'd15796,17'd54035,17'd54036,17'd54037,17'd13872,17'd54038,17'd54039,17'd53830,17'd53969,17'd11502,17'd24532,17'd24851,17'd12712,17'd12712,17'd17226,17'd12711,17'd12094,17'd23676,17'd20897,17'd24357,17'd54040,17'd54041,17'd54042,17'd54043,17'd17234,17'd17476,17'd17013,17'd17013,17'd17013,17'd16914,17'd13643,17'd13760,17'd13252,17'd12106,17'd20314,17'd22818,17'd23512,17'd24859,17'd24537,17'd27004,17'd28816,17'd29066,17'd31587,17'd31127,17'd54044,17'd52867,17'd52868,17'd53321,17'd53472,17'd53709,17'd53628,17'd53322,17'd52868,17'd53473,17'd50951,17'd34545,17'd32283,17'd30972,17'd30971,17'd26873,17'd24538,17'd25926,17'd21361,17'd16325,17'd15185,17'd16326,17'd11397,17'd11396,17'd14673,17'd11274,17'd11395,17'd11666,17'd11961,17'd12110,17'd12414,17'd12109,17'd11806,17'd10854,17'd10023,17'd18196,17'd15431,17'd14928,17'd14928,17'd11276,17'd18916,17'd10167,17'd10991,17'd11132,17'd10854,17'd10990,17'd14673,17'd13137,17'd13764,17'd11807,17'd11964,17'd11807,17'd16069,17'd11808,17'd11520,17'd10736,17'd10479,17'd24361,17'd22993,17'd15946,17'd8737,17'd54045,17'd15950,17'd14683,17'd16567,17'd15060,17'd21988,17'd54046,17'd54047,17'd25681,17'd54048,17'd54049,17'd54050,17'd54051,17'd54052,17'd24052,17'd22484,17'd54053,17'd53258,17'd53838,17'd54054,17'd54055,17'd54056,17'd54057,17'd32353,17'd43157,17'd49171,17'd54058,17'd53844,17'd48536,17'd50164,17'd50907,17'd43279,17'd43012,17'd50736,17'd49683,17'd49390,17'd47641,17'd46946,17'd53336,17'd32826,17'd27642,17'd31503,17'd31503,17'd27885,17'd28134,17'd33654,17'd32192,17'd29247,17'd28372,17'd29536,17'd30131,17'd34117,17'd49790,17'd29979,17'd36132,17'd29978,17'd30131,17'd30131,17'd30131,17'd30131,17'd30131,17'd30131,17'd30131,17'd30738,17'd36132,17'd32193,17'd32354,17'd32506,17'd31353,17'd26782,17'd27883,17'd27640,17'd27514,17'd27514,17'd27259,17'd26902,17'd31035,17'd29379,17'd31503,17'd31503,17'd33476,17'd44103,17'd45152,17'd45479,17'd47054,17'd48904,17'd49478,17'd50272,17'd52675,17'd51830,17'd51995,17'd50267,17'd48361,17'd48152,17'd54059,17'd51387,17'd54060,17'd50153,17'd46659,17'd53486,17'd54061,17'd23917,17'd23566,17'd29973,17'd36426,17'd39132,17'd36987,17'd23565,17'd24086,17'd30879,17'd24743,17'd32007,17'd25180,17'd24895,17'd24415,17'd34137,17'd32351,17'd22680,17'd22159,17'd23222,17'd22864,17'd48164,17'd54062,17'd53723,17'd53992,17'd21387,17'd21535,17'd53653,17'd54063,17'd51911,17'd54064,17'd54065,17'd54066,17'd54067,17'd54068,17'd54069,17'd54070,17'd54071,17'd26820,17'd54072,17'd53923,17'd54073,17'd54074,17'd25877,17'd11294,17'd5608,17'd4839,17'd5322,17'd7822,17'd24475,17'd24149,17'd5323,17'd4841,17'd5002,17'd5004,17'd30333,17'd6554,17'd9091,17'd32073,17'd9091,17'd9091,17'd6219,17'd6390,17'd9091,17'd7668,17'd27696,17'd29740,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd7499,17'd37152,17'd31891,17'd6554,17'd5614,17'd27935,17'd5335,17'd30180,17'd31552,17'd4842,17'd5166,17'd5166,17'd5012,17'd53733,17'd52011,17'd54075,17'd48726,17'd54076,17'd54077,17'd54006,17'd54078,17'd54079,17'd54080,17'd54081,17'd54082,17'd54083,17'd54084,17'd53938,17'd54085,17'd40997,17'd54086,17'd53870,17'd52916,17'd51252,17'd40562,17'd3567,17'd54014,17'd54015,17'd6239,17'd4059,17'd38071,17'd38071,17'd38071,17'd4059,17'd4059,17'd4059,17'd38071,17'd2558,17'd1120,17'd960,17'd797,17'd237,17'd630,17'd448,17'd628,17'd38071,17'd4399,17'd4399,17'd6239,17'd6084,17'd53152,17'd35206,17'd53594,17'd53941,17'd53942,17'd53872,17'd53873,17'd54087,17'd53804,17'd53752
},
'{
17'd15877,17'd3427,17'd10802,17'd3429,17'd2258,17'd27442,17'd652,17'd652,17'd980,17'd27,17'd286,17'd286,17'd285,17'd285,17'd285,17'd467,17'd285,17'd285,17'd286,17'd286,17'd4430,17'd4430,17'd4431,17'd4091,17'd6278,17'd3910,17'd3434,17'd2944,17'd17300,17'd2265,17'd2265,17'd1974,17'd1840,17'd2433,17'd1424,17'd1706,17'd1707,17'd3600,17'd36605,17'd54088,17'd14753,17'd2802,17'd5531,17'd54089,17'd54016,17'd13825,17'd13588,17'd54090,17'd54091,17'd42485,17'd54092,17'd22630,17'd12814,17'd24345,17'd15763,17'd22802,17'd11476,17'd11626,17'd14621,17'd12955,17'd12678,17'd12357,17'd14344,17'd13461,17'd13460,17'd12355,17'd12677,17'd12954,17'd14621,17'd12530,17'd12360,17'd12065,17'd12065,17'd23154,17'd12362,17'd22630,17'd28438,17'd28667,17'd12532,17'd12681,17'd17204,17'd17205,17'd19255,17'd27833,17'd18776,17'd18776,17'd16165,17'd47673,17'd34179,17'd50005,17'd48932,17'd54093,17'd53757,17'd54094,17'd54095,17'd54096,17'd2979,17'd54023,17'd54097,17'd5263,17'd54098,17'd54099,17'd53885,17'd53958,17'd54100,17'd54101,17'd46253,17'd53889,17'd53306,17'd54030,17'd54102,17'd54103,17'd54104,17'd53762,17'd48192,17'd6792,17'd38895,17'd37597,17'd54105,17'd50098,17'd30662,17'd54106,17'd52037,17'd22805,17'd26356,17'd25917,17'd53312,17'd53764,17'd53765,17'd54107,17'd11106,17'd54108,17'd54109,17'd13991,17'd54039,17'd11502,17'd11502,17'd11502,17'd54110,17'd24852,17'd11939,17'd12711,17'd17226,17'd12710,17'd20903,17'd54111,17'd54112,17'd21200,17'd53623,17'd54113,17'd53899,17'd54114,17'd18331,17'd17476,17'd53708,17'd53708,17'd17724,17'd16560,17'd30378,17'd13643,17'd13252,17'd12106,17'd17474,17'd12107,17'd23512,17'd24859,17'd24856,17'd27004,17'd26370,17'd29923,17'd29645,17'd30676,17'd34380,17'd50952,17'd52301,17'd54115,17'd53032,17'd54116,17'd53393,17'd53321,17'd52869,17'd52401,17'd50951,17'd49525,17'd33875,17'd30677,17'd31285,17'd28691,17'd27123,17'd22819,17'd22992,17'd14261,17'd11806,17'd16326,17'd21985,17'd11396,17'd11523,17'd14810,17'd11519,17'd16198,17'd12112,17'd12110,17'd12418,17'd12109,17'd11961,17'd14673,17'd17720,17'd17839,17'd25530,17'd19642,17'd10479,17'd11528,17'd9883,17'd10167,17'd11133,17'd19282,17'd11399,17'd11524,17'd11274,17'd16069,17'd14669,17'd17125,17'd11807,17'd11807,17'd17125,17'd11275,17'd14262,17'd14931,17'd17720,17'd53547,17'd8732,17'd16076,17'd54117,17'd54118,17'd13771,17'd15061,17'd12728,17'd19036,17'd25152,17'd54046,17'd16447,17'd15303,17'd54048,17'd54119,17'd53981,17'd54120,17'd21510,17'd54121,17'd54122,17'd11004,17'd19655,17'd54123,17'd54124,17'd54125,17'd54126,17'd54127,17'd54128,17'd48695,17'd54129,17'd53989,17'd48360,17'd49691,17'd50907,17'd54130,17'd43417,17'd43012,17'd50164,17'd51648,17'd39575,17'd53560,17'd39903,17'd41271,17'd31352,17'd29977,17'd27642,17'd27642,17'd27885,17'd32192,17'd33655,17'd33321,17'd29380,17'd28728,17'd29831,17'd29978,17'd49790,17'd49579,17'd29831,17'd36132,17'd29978,17'd29978,17'd29978,17'd29978,17'd29978,17'd29978,17'd29978,17'd29978,17'd36132,17'd28372,17'd33654,17'd32832,17'd39437,17'd26781,17'd33815,17'd27514,17'd26530,17'd26530,17'd27514,17'd27640,17'd26902,17'd31035,17'd31352,17'd31352,17'd38025,17'd43696,17'd43974,17'd44587,17'd45369,17'd47343,17'd49382,17'd49683,17'd50371,17'd53341,17'd51830,17'd50468,17'd49389,17'd54131,17'd48252,17'd54132,17'd54133,17'd54134,17'd53116,17'd54135,17'd52742,17'd48987,17'd30275,17'd29830,17'd32667,17'd32830,17'd32504,17'd23923,17'd23733,17'd23732,17'd30879,17'd24742,17'd32007,17'd25032,17'd24745,17'd24090,17'd34137,17'd29828,17'd22856,17'd22683,17'd48912,17'd32010,17'd48276,17'd54136,17'd54137,17'd53913,17'd53131,17'd21999,17'd53495,17'd54138,17'd54139,17'd51903,17'd54140,17'd54141,17'd54142,17'd54143,17'd54144,17'd54145,17'd54146,17'd54147,17'd54148,17'd54149,17'd54073,17'd48172,17'd22413,17'd8608,17'd5757,17'd4525,17'd5754,17'd54150,17'd23974,17'd4679,17'd4682,17'd4687,17'd5002,17'd5004,17'd30638,17'd6390,17'd9091,17'd9091,17'd6219,17'd6219,17'd6390,17'd6390,17'd9091,17'd7668,17'd27696,17'd35052,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd7499,17'd7668,17'd6219,17'd31891,17'd30333,17'd27935,17'd27935,17'd28185,17'd5335,17'd28536,17'd31552,17'd4842,17'd5166,17'd5167,17'd5011,17'd53733,17'd49705,17'd49103,17'd3684,17'd54151,17'd54077,17'd54152,17'd54153,17'd54154,17'd54155,17'd54156,17'd54157,17'd54158,17'd54159,17'd54160,17'd54161,17'd54162,17'd41476,17'd53870,17'd52916,17'd51252,17'd40562,17'd3567,17'd54014,17'd54163,17'd3711,17'd3874,17'd38071,17'd38071,17'd4059,17'd52698,17'd4059,17'd4059,17'd4398,17'd2558,17'd628,17'd1265,17'd237,17'd237,17'd236,17'd629,17'd1120,17'd4398,17'd4399,17'd4399,17'd6239,17'd6084,17'd53152,17'd35206,17'd53594,17'd53747,17'd53871,17'd53872,17'd54164,17'd53598,17'd54165,17'd54166
},
'{
17'd15877,17'd3427,17'd10802,17'd3429,17'd2258,17'd2425,17'd29,17'd652,17'd652,17'd980,17'd27,17'd286,17'd285,17'd285,17'd467,17'd467,17'd285,17'd285,17'd1833,17'd286,17'd4430,17'd4430,17'd4431,17'd4091,17'd3910,17'd3910,17'd3434,17'd2601,17'd2265,17'd19874,17'd19874,17'd1702,17'd1840,17'd2433,17'd1424,17'd35772,17'd1707,17'd3600,17'd3110,17'd30050,17'd14993,17'd13956,17'd4591,17'd20877,17'd54167,17'd13959,17'd13587,17'd54168,17'd54169,17'd42485,17'd54170,17'd19382,17'd12956,17'd24345,17'd15763,17'd15763,17'd11476,17'd11626,17'd12218,17'd14890,17'd15516,17'd12357,17'd13597,17'd13461,17'd12214,17'd12355,17'd12677,17'd12813,17'd12218,17'd11627,17'd12530,17'd12218,17'd12814,17'd23154,17'd12815,17'd16658,17'd28438,17'd18884,17'd18884,17'd17204,17'd11087,17'd16766,17'd25512,17'd27833,17'd18776,17'd15902,17'd14765,17'd47673,17'd34357,17'd48819,17'd54171,17'd54172,17'd53757,17'd53522,17'd53448,17'd54173,17'd2978,17'd54174,17'd54175,17'd2476,17'd54176,17'd54026,17'd53884,17'd53958,17'd5862,17'd54177,17'd54178,17'd54179,17'd54180,17'd54181,17'd54181,17'd54182,17'd6650,17'd54183,17'd53615,17'd54184,17'd40278,17'd50398,17'd54185,17'd52938,17'd51423,17'd27840,17'd51782,17'd27223,17'd22289,17'd26249,17'd53312,17'd54186,17'd15926,17'd54187,17'd54188,17'd54189,17'd19636,17'd14247,17'd54039,17'd25669,17'd54190,17'd11502,17'd54191,17'd12090,17'd11788,17'd12710,17'd12570,17'd12711,17'd20902,17'd13131,17'd54192,17'd20897,17'd24697,17'd53466,17'd53468,17'd53976,17'd39072,17'd17969,17'd53708,17'd53708,17'd17724,17'd53102,17'd13642,17'd30378,17'd15570,17'd17348,17'd17474,17'd12107,17'd23512,17'd24537,17'd24856,17'd27004,17'd26370,17'd28816,17'd28460,17'd29330,17'd31289,17'd31590,17'd50951,17'd53545,17'd52800,17'd53320,17'd52799,17'd52799,17'd52869,17'd52302,17'd52300,17'd50111,17'd31590,17'd33568,17'd30972,17'd31290,17'd26873,17'd23512,17'd25926,17'd24995,17'd11960,17'd12582,17'd19643,17'd11396,17'd16068,17'd12720,17'd11519,17'd11666,17'd13363,17'd12110,17'd12253,17'd12579,17'd11960,17'd11807,17'd10739,17'd10741,17'd11528,17'd10479,17'd9883,17'd11528,17'd10329,17'd20754,17'd10329,17'd19532,17'd11132,17'd21206,17'd21206,17'd11274,17'd13137,17'd17125,17'd13762,17'd13762,17'd17125,17'd11274,17'd11130,17'd14931,17'd10991,17'd15187,17'd24214,17'd16333,17'd10996,17'd54193,17'd14818,17'd17133,17'd13894,17'd19646,17'd16447,17'd12589,17'd16447,17'd13377,17'd18205,17'd54194,17'd54195,17'd16694,17'd14142,17'd54196,17'd18337,17'd54197,17'd54198,17'd51986,17'd54199,17'd54200,17'd40224,17'd54201,17'd54202,17'd53906,17'd54203,17'd48451,17'd49289,17'd49986,17'd42874,17'd43143,17'd54130,17'd43012,17'd49987,17'd48536,17'd40814,17'd49078,17'd45483,17'd35011,17'd31503,17'd32354,17'd27642,17'd27642,17'd32832,17'd32354,17'd53491,17'd32193,17'd28372,17'd29536,17'd29978,17'd29978,17'd49790,17'd49579,17'd29831,17'd36132,17'd29978,17'd29978,17'd29978,17'd29978,17'd29978,17'd29978,17'd30130,17'd31038,17'd28857,17'd28855,17'd33319,17'd32356,17'd28486,17'd28009,17'd27639,17'd25949,17'd27767,17'd26062,17'd27514,17'd43290,17'd26781,17'd31035,17'd30735,17'd31035,17'd32005,17'd45484,17'd39583,17'd44100,17'd48609,17'd48535,17'd50467,17'd50468,17'd52000,17'd52675,17'd50268,17'd49794,17'd49090,17'd54204,17'd49472,17'd51310,17'd54205,17'd54206,17'd53486,17'd54135,17'd53193,17'd34883,17'd28976,17'd32352,17'd36426,17'd36426,17'd32352,17'd29242,17'd31033,17'd28722,17'd28852,17'd24742,17'd32007,17'd25032,17'd24744,17'd29100,17'd29242,17'd29828,17'd22332,17'd32009,17'd48912,17'd22512,17'd54207,17'd53115,17'd54208,17'd54209,17'd52594,17'd54210,17'd54211,17'd54212,17'd54213,17'd54214,17'd54215,17'd54216,17'd54217,17'd54218,17'd54219,17'd54220,17'd54221,17'd54222,17'd54148,17'd54223,17'd54224,17'd54225,17'd11692,17'd8608,17'd24648,17'd4837,17'd4521,17'd54226,17'd4677,17'd24796,17'd4683,17'd5002,17'd5004,17'd30637,17'd28185,17'd6390,17'd32073,17'd9091,17'd6220,17'd6219,17'd6390,17'd32073,17'd7499,17'd27696,17'd27696,17'd35052,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd7499,17'd7668,17'd6390,17'd33369,17'd31553,17'd28185,17'd27935,17'd5160,17'd5334,17'd5152,17'd31716,17'd4842,17'd5166,17'd5169,17'd37944,17'd4693,17'd54227,17'd54228,17'd54229,17'd38197,17'd54230,17'd54231,17'd54232,17'd54233,17'd54234,17'd54235,17'd54236,17'd54237,17'd2072,17'd54238,17'd54161,17'd41621,17'd54086,17'd53870,17'd54239,17'd51252,17'd40562,17'd3567,17'd39326,17'd5627,17'd3711,17'd3874,17'd38071,17'd38071,17'd4059,17'd52698,17'd52698,17'd4059,17'd2558,17'd5775,17'd796,17'd237,17'd237,17'd237,17'd236,17'd628,17'd38071,17'd4398,17'd4399,17'd4399,17'd6239,17'd54240,17'd53152,17'd35206,17'd53594,17'd53747,17'd53871,17'd53872,17'd54164,17'd54241,17'd54165,17'd54166
},
'{
17'd54242,17'd10925,17'd10670,17'd3429,17'd2258,17'd2425,17'd17,17'd3905,17'd652,17'd652,17'd27,17'd286,17'd285,17'd285,17'd7385,17'd7385,17'd285,17'd285,17'd285,17'd285,17'd7060,17'd7060,17'd4430,17'd4430,17'd4091,17'd3755,17'd3434,17'd2601,17'd2785,17'd2600,17'd2121,17'd2121,17'd1702,17'd1283,17'd1284,17'd18150,17'd1560,17'd1708,17'd3440,17'd30504,17'd54243,17'd28663,17'd3767,17'd54244,17'd49410,17'd24515,17'd13314,17'd54245,17'd21648,17'd48077,17'd54246,17'd25512,17'd11629,17'd54247,17'd22802,17'd22802,17'd11476,17'd11626,17'd11477,17'd11477,17'd19127,17'd12357,17'd13597,17'd14344,17'd54248,17'd13716,17'd12062,17'd10941,17'd15640,17'd11362,17'd12532,17'd16765,17'd13211,17'd12955,17'd13094,17'd13969,17'd20422,17'd20148,17'd20886,17'd17204,17'd10944,17'd19754,17'd30511,17'd54249,17'd17690,17'd14347,17'd14346,17'd15900,17'd54250,17'd54251,17'd54252,17'd54253,17'd54254,17'd54255,17'd53163,17'd53953,17'd54256,17'd54257,17'd54258,17'd54259,17'd5094,17'd54260,17'd54261,17'd54262,17'd5861,17'd54263,17'd54264,17'd54265,17'd54266,17'd54267,17'd54268,17'd54181,17'd54182,17'd53822,17'd53615,17'd54269,17'd54270,17'd54271,17'd54272,17'd50198,17'd30207,17'd27606,17'd28085,17'd28444,17'd50301,17'd26357,17'd19910,17'd54186,17'd18670,17'd15796,17'd15927,17'd10828,17'd54273,17'd11109,17'd26362,17'd26489,17'd53702,17'd53829,17'd54274,17'd54275,17'd23677,17'd17833,17'd17226,17'd12570,17'd13638,17'd20903,17'd13359,17'd21980,17'd23508,17'd24696,17'd54276,17'd54277,17'd54278,17'd38503,17'd38367,17'd18685,17'd40136,17'd40136,17'd17349,17'd38239,17'd14526,17'd13252,17'd12106,17'd12106,17'd14807,17'd12254,17'd24856,17'd26370,17'd26370,17'd28816,17'd27857,17'd28818,17'd29067,17'd34381,17'd34545,17'd49033,17'd51603,17'd51513,17'd52303,17'd54279,17'd52402,17'd52401,17'd52400,17'd53394,17'd34705,17'd33095,17'd34835,17'd30974,17'd28462,17'd26629,17'd24859,17'd29781,17'd21671,17'd17722,17'd18681,17'd11964,17'd10989,17'd10989,17'd14262,17'd11667,17'd11960,17'd12580,17'd12579,17'd12414,17'd13882,17'd12861,17'd10737,17'd27859,17'd10326,17'd10478,17'd10329,17'd10329,17'd20756,17'd11134,17'd11134,17'd10330,17'd10330,17'd10991,17'd10991,17'd19532,17'd12720,17'd13000,17'd11666,17'd10989,17'd11520,17'd16069,17'd11524,17'd11132,17'd10476,17'd11277,17'd9046,17'd26262,17'd15692,17'd54280,17'd20051,17'd24049,17'd7463,17'd20049,17'd21058,17'd21210,17'd52405,17'd19536,17'd14683,17'd7958,17'd15307,17'd54281,17'd9353,17'd54282,17'd20758,17'd54283,17'd54284,17'd52072,17'd53417,17'd54285,17'd24421,17'd37390,17'd54202,17'd54286,17'd53989,17'd48153,17'd49692,17'd50072,17'd52506,17'd50370,17'd42875,17'd50475,17'd54287,17'd40507,17'd54288,17'd44226,17'd30726,17'd31354,17'd33001,17'd38813,17'd38813,17'd39284,17'd27885,17'd28134,17'd28134,17'd32017,17'd32018,17'd34285,17'd32508,17'd32508,17'd29690,17'd29690,17'd29831,17'd29831,17'd29979,17'd49579,17'd30130,17'd30130,17'd29831,17'd36132,17'd31038,17'd29537,17'd33654,17'd33001,17'd32356,17'd35426,17'd28482,17'd30734,17'd28720,17'd28594,17'd28602,17'd26062,17'd26530,17'd28725,17'd33163,17'd28486,17'd26901,17'd32343,17'd40826,17'd46546,17'd45609,17'd43422,17'd49174,17'd43281,17'd50267,17'd50268,17'd52675,17'd51741,17'd50568,17'd49484,17'd46656,17'd54289,17'd51311,17'd54290,17'd54291,17'd52743,17'd53486,17'd52669,17'd34282,17'd24086,17'd29830,17'd38976,17'd32830,17'd39278,17'd23385,17'd28975,17'd29100,17'd28975,17'd24743,17'd28851,17'd32007,17'd32007,17'd24417,17'd28975,17'd38669,17'd39590,17'd34454,17'd31497,17'd41726,17'd34280,17'd54292,17'd54293,17'd54294,17'd54295,17'd54296,17'd21533,17'd51067,17'd54297,17'd54298,17'd51980,17'd54299,17'd54300,17'd54301,17'd54302,17'd54303,17'd54304,17'd54305,17'd22906,17'd54306,17'd54307,17'd54308,17'd47848,17'd12741,17'd54309,17'd9502,17'd23457,17'd54310,17'd54311,17'd4679,17'd6067,17'd4687,17'd4842,17'd30637,17'd5160,17'd28185,17'd27935,17'd6390,17'd6220,17'd9091,17'd32073,17'd32073,17'd32074,17'd29740,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd29593,17'd31888,17'd31888,17'd31888,17'd31888,17'd27696,17'd7499,17'd7499,17'd6554,17'd31400,17'd5167,17'd5166,17'd5163,17'd5161,17'd34921,17'd5155,17'd34791,17'd5008,17'd5165,17'd5170,17'd37697,17'd52522,17'd38571,17'd47264,17'd54312,17'd3191,17'd54313,17'd54314,17'd54315,17'd54316,17'd54317,17'd54318,17'd54319,17'd54320,17'd2072,17'd54321,17'd54322,17'd40997,17'd53672,17'd54323,17'd54324,17'd51252,17'd40410,17'd54325,17'd2390,17'd38856,17'd3874,17'd1120,17'd38071,17'd4059,17'd54326,17'd54326,17'd1264,17'd795,17'd1944,17'd629,17'd18144,17'd52461,17'd237,17'd630,17'd628,17'd1120,17'd1402,17'd1402,17'd4398,17'd4398,17'd53293,17'd54240,17'd54327,17'd35206,17'd54328,17'd54329,17'd53518,17'd54330,17'd54331,17'd54241,17'd54332,17'd54333
},
'{
17'd16010,17'd10925,17'd10802,17'd3593,17'd3429,17'd2258,17'd1414,17'd1416,17'd653,17'd652,17'd27,17'd27,17'd26,17'd26,17'd7385,17'd7385,17'd285,17'd285,17'd285,17'd285,17'd7060,17'd7060,17'd4430,17'd4430,17'd4091,17'd3755,17'd3434,17'd2601,17'd2785,17'd2121,17'd1971,17'd1971,17'd1702,17'd1283,17'd1284,17'd18150,17'd18150,17'd1560,17'd34168,17'd48292,17'd54334,17'd54335,17'd27717,17'd54336,17'd54337,17'd49411,17'd16508,17'd54338,17'd21182,17'd48473,17'd54339,17'd27833,17'd19754,17'd10690,17'd12527,17'd22802,17'd11476,17'd54340,17'd54341,17'd11477,17'd54342,17'd22802,17'd12357,17'd13597,17'd13838,17'd13716,17'd11762,17'd10281,17'd12066,17'd11362,17'd18884,17'd29048,17'd13211,17'd12955,17'd12218,17'd11628,17'd18774,17'd19893,17'd20886,17'd19893,17'd11231,17'd21964,17'd30511,17'd54249,17'd16169,17'd14346,17'd15641,17'd54343,17'd54344,17'd54345,17'd54346,17'd54347,17'd54348,17'd54349,17'd54350,17'd54094,17'd3636,17'd3638,17'd54351,17'd3490,17'd3963,17'd54352,17'd54353,17'd54354,17'd54355,17'd54356,17'd54357,17'd54358,17'd54359,17'd54360,17'd54268,17'd54361,17'd54181,17'd41648,17'd53615,17'd54269,17'd54362,17'd54363,17'd54364,17'd54365,17'd50851,17'd29766,17'd28557,17'd54366,17'd50100,17'd25807,17'd54367,17'd18431,17'd10578,17'd10579,17'd15665,17'd10711,17'd15284,17'd11377,17'd26362,17'd54368,17'd53701,17'd54369,17'd54274,17'd54275,17'd54370,17'd23848,17'd11650,17'd12570,17'd13638,17'd20903,17'd13131,17'd54111,17'd54371,17'd24022,17'd54372,17'd54373,17'd54374,17'd39072,17'd38503,17'd18685,17'd40136,17'd40136,17'd54375,17'd40744,17'd14809,17'd13517,17'd12106,17'd12106,17'd14807,17'd12254,17'd24856,17'd26370,17'd29778,17'd28816,17'd28104,17'd27857,17'd28461,17'd31440,17'd48660,17'd38498,17'd54376,17'd35100,17'd52134,17'd54377,17'd52303,17'd52302,17'd53473,17'd53473,17'd53394,17'd36936,17'd33568,17'd30677,17'd31768,17'd28460,17'd27004,17'd28817,17'd22819,17'd20314,17'd18443,17'd16326,17'd13516,17'd10989,17'd11964,17'd15185,17'd15053,17'd14130,17'd12579,17'd12414,17'd13882,17'd20313,17'd15810,17'd41193,17'd10474,17'd14518,17'd10330,17'd10330,17'd11528,17'd10479,17'd11135,17'd19642,17'd9883,17'd11528,17'd11133,17'd24996,17'd14810,17'd12862,17'd11666,17'd14262,17'd11520,17'd16068,17'd11524,17'd11132,17'd10739,17'd9883,17'd17607,17'd37734,17'd54378,17'd54379,17'd21212,17'd15697,17'd54380,17'd12729,17'd54381,17'd54382,17'd15946,17'd19536,17'd14816,17'd14817,17'd15951,17'd54281,17'd9353,17'd11815,17'd21372,17'd54383,17'd54384,17'd54385,17'd21698,17'd23924,17'd29528,17'd33793,17'd54386,17'd54387,17'd54388,17'd43541,17'd49984,17'd50574,17'd50271,17'd49985,17'd50907,17'd54389,17'd54390,17'd47239,17'd44697,17'd44700,17'd54391,17'd26652,17'd33001,17'd38672,17'd38813,17'd54392,17'd27885,17'd27885,17'd28134,17'd32355,17'd29248,17'd29249,17'd32833,17'd32508,17'd29690,17'd29690,17'd29536,17'd29536,17'd29690,17'd30280,17'd30130,17'd29690,17'd29831,17'd36132,17'd28728,17'd28981,17'd33001,17'd31354,17'd37908,17'd28853,17'd28481,17'd27638,17'd28130,17'd28600,17'd28602,17'd26062,17'd27514,17'd28853,17'd30586,17'd26902,17'd26902,17'd32006,17'd41270,17'd53336,17'd39433,17'd43152,17'd49279,17'd49093,17'd50164,17'd51157,17'd51741,17'd50272,17'd49890,17'd49288,17'd52750,17'd51155,17'd53782,17'd54393,17'd50361,17'd50154,17'd52967,17'd54394,17'd33317,17'd34137,17'd29531,17'd32504,17'd36426,17'd23217,17'd29972,17'd23562,17'd28601,17'd34884,17'd24743,17'd25032,17'd25180,17'd25030,17'd24744,17'd29100,17'd42449,17'd39590,17'd31834,17'd21845,17'd54395,17'd35294,17'd54396,17'd54397,17'd54398,17'd54399,17'd21999,17'd21702,17'd51067,17'd51468,17'd54400,17'd52594,17'd54401,17'd29139,17'd54402,17'd54403,17'd54404,17'd54405,17'd54406,17'd54407,17'd54408,17'd22751,17'd54409,17'd54410,17'd53925,17'd26583,17'd54411,17'd23277,17'd24147,17'd7822,17'd4837,17'd42910,17'd4686,17'd4842,17'd30637,17'd25627,17'd28185,17'd27935,17'd6390,17'd6219,17'd32073,17'd32073,17'd34658,17'd32074,17'd29740,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd29593,17'd29593,17'd31888,17'd31888,17'd31888,17'd27696,17'd7668,17'd6220,17'd30638,17'd31400,17'd5167,17'd5009,17'd5163,17'd5161,17'd4530,17'd49804,17'd34791,17'd5008,17'd5164,17'd5170,17'd37697,17'd51177,17'd52689,17'd53216,17'd54412,17'd54413,17'd54414,17'd54415,17'd54416,17'd54417,17'd54418,17'd54318,17'd54319,17'd54320,17'd54419,17'd54321,17'd54420,17'd54421,17'd41902,17'd54323,17'd54324,17'd51252,17'd40410,17'd54422,17'd53675,17'd1943,17'd628,17'd628,17'd38071,17'd4059,17'd54326,17'd54326,17'd1264,17'd1402,17'd1944,17'd629,17'd6867,17'd36902,17'd237,17'd630,17'd628,17'd1120,17'd1402,17'd1402,17'd4398,17'd4398,17'd53293,17'd54240,17'd54327,17'd35058,17'd54328,17'd54329,17'd54423,17'd54330,17'd54424,17'd54425,17'd54332,17'd54426
},
'{
17'd16010,17'd10924,17'd10802,17'd3429,17'd2258,17'd2426,17'd1414,17'd1416,17'd653,17'd652,17'd27,17'd27,17'd26,17'd26,17'd285,17'd285,17'd285,17'd285,17'd285,17'd285,17'd7060,17'd7060,17'd4430,17'd4430,17'd4091,17'd3755,17'd3434,17'd2601,17'd2785,17'd2600,17'd2121,17'd1971,17'd1702,17'd1283,17'd1284,17'd18150,17'd18150,17'd1560,17'd1561,17'd32254,17'd30050,17'd13308,17'd28663,17'd54427,17'd54428,17'd49714,17'd19374,17'd17194,17'd21806,17'd48473,17'd54429,17'd17445,17'd10944,17'd11914,17'd12679,17'd14469,17'd12527,17'd11626,17'd11360,17'd11477,17'd54342,17'd14469,17'd13597,17'd13718,17'd15135,17'd13716,17'd10687,17'd10281,17'd12066,17'd18412,17'd19006,17'd16027,17'd15383,17'd19890,17'd14621,17'd14471,17'd20422,17'd17689,17'd20886,17'd17317,17'd16766,17'd21649,17'd30511,17'd54249,17'd16411,17'd15641,17'd15641,17'd24195,17'd54344,17'd54430,17'd54431,17'd54432,17'd54433,17'd54434,17'd53756,17'd53952,17'd54435,17'd54436,17'd54437,17'd2998,17'd2660,17'd2160,17'd54438,17'd5698,17'd54439,17'd54440,17'd54441,17'd54442,17'd54443,17'd54444,17'd54268,17'd54445,17'd54446,17'd54103,17'd54033,17'd54447,17'd54448,17'd50008,17'd53454,17'd54449,17'd54450,17'd54451,17'd27965,17'd29461,17'd9455,17'd9716,17'd10135,17'd53764,17'd54452,17'd10579,17'd54453,17'd54454,17'd54455,17'd14369,17'd15286,17'd53701,17'd53621,17'd54456,17'd53969,17'd54275,17'd54275,17'd20601,17'd54457,17'd54458,17'd19914,17'd12093,17'd13506,17'd13131,17'd23676,17'd23675,17'd54459,17'd54460,17'd54461,17'd53707,17'd45933,17'd17969,17'd53708,17'd53708,17'd17476,17'd16686,17'd14525,17'd13517,17'd15685,17'd15685,17'd17348,17'd12254,17'd24856,17'd26370,17'd28816,17'd28816,17'd28104,17'd28104,17'd35372,17'd29067,17'd31761,17'd36490,17'd35933,17'd34833,17'd51432,17'd52134,17'd51693,17'd51693,17'd52401,17'd51602,17'd51603,17'd53250,17'd34203,17'd31767,17'd31285,17'd28345,17'd28103,17'd36935,17'd23512,17'd19408,17'd16325,17'd16326,17'd11397,17'd11274,17'd11964,17'd16326,17'd18917,17'd11960,17'd12109,17'd12109,17'd13882,17'd15564,17'd15186,17'd20910,17'd16555,17'd10476,17'd11670,17'd10330,17'd11528,17'd10479,17'd19642,17'd51697,17'd9883,17'd11134,17'd10326,17'd10166,17'd10604,17'd12720,17'd11666,17'd11395,17'd11395,17'd16068,17'd11524,17'd11399,17'd10739,17'd17839,17'd16067,17'd23343,17'd16207,17'd53635,17'd54462,17'd54463,17'd54464,17'd8112,17'd14388,17'd54465,17'd21508,17'd25681,17'd14266,17'd14684,17'd7795,17'd54466,17'd7959,17'd54467,17'd54468,17'd54469,17'd54470,17'd54471,17'd54472,17'd54473,17'd30424,17'd34459,17'd54474,17'd54132,17'd49581,17'd49693,17'd50659,17'd50370,17'd49987,17'd49985,17'd42874,17'd54475,17'd54476,17'd48358,17'd48897,17'd33942,17'd31494,17'd26523,17'd33001,17'd32354,17'd30279,17'd29977,17'd30279,17'd30279,17'd28134,17'd32355,17'd32507,17'd33486,17'd29690,17'd29690,17'd29690,17'd30884,17'd28857,17'd29536,17'd29979,17'd30738,17'd29979,17'd30884,17'd36132,17'd29536,17'd29105,17'd27636,17'd33952,17'd35570,17'd33163,17'd41999,17'd27513,17'd28594,17'd27765,17'd28600,17'd26064,17'd25949,17'd27515,17'd28853,17'd27027,17'd27371,17'd28725,17'd33478,17'd44228,17'd48044,17'd39737,17'd42596,17'd47937,17'd51648,17'd50365,17'd51830,17'd50371,17'd50072,17'd51077,17'd52676,17'd54477,17'd49472,17'd54478,17'd54479,17'd54480,17'd50154,17'd52967,17'd33802,17'd31033,17'd29826,17'd42744,17'd33651,17'd29973,17'd23388,17'd23384,17'd28852,17'd34467,17'd24743,17'd24743,17'd25031,17'd25180,17'd24895,17'd28851,17'd29100,17'd41874,17'd46966,17'd36566,17'd31658,17'd23042,17'd42440,17'd54481,17'd54482,17'd54483,17'd54484,17'd54485,17'd54486,17'd51563,17'd51631,17'd54487,17'd54488,17'd54489,17'd54490,17'd54491,17'd54492,17'd54493,17'd54494,17'd20361,17'd35463,17'd22402,17'd54495,17'd54496,17'd12443,17'd53925,17'd26111,17'd23108,17'd23456,17'd9764,17'd54497,17'd4837,17'd4995,17'd4686,17'd4842,17'd30637,17'd25627,17'd28185,17'd27935,17'd6390,17'd6219,17'd32073,17'd32073,17'd32074,17'd29740,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd29593,17'd29593,17'd31888,17'd31888,17'd27696,17'd27696,17'd8780,17'd6219,17'd32553,17'd30180,17'd42031,17'd37153,17'd5162,17'd27697,17'd4690,17'd49804,17'd40397,17'd37029,17'd5164,17'd5011,17'd54498,17'd54499,17'd54500,17'd51179,17'd54501,17'd54502,17'd54503,17'd54504,17'd54505,17'd54506,17'd54507,17'd54508,17'd54509,17'd54510,17'd54511,17'd54321,17'd54512,17'd54513,17'd53672,17'd51182,17'd52614,17'd3217,17'd40410,17'd54514,17'd2557,17'd18144,17'd629,17'd628,17'd38071,17'd4059,17'd54326,17'd54326,17'd795,17'd8015,17'd54515,17'd448,17'd36748,17'd36902,17'd237,17'd235,17'd628,17'd628,17'd1402,17'd1825,17'd4398,17'd4398,17'd6239,17'd54516,17'd54327,17'd35058,17'd54517,17'd54329,17'd54518,17'd54519,17'd54424,17'd1938,17'd54520,17'd54426
},
'{
17'd16010,17'd10925,17'd10670,17'd10669,17'd52621,17'd2426,17'd1414,17'd2257,17'd289,17'd653,17'd980,17'd27,17'd26,17'd26,17'd285,17'd285,17'd285,17'd285,17'd285,17'd285,17'd7060,17'd7060,17'd4430,17'd4430,17'd4091,17'd3755,17'd3434,17'd2601,17'd2785,17'd2600,17'd2121,17'd1971,17'd1702,17'd1557,17'd14449,17'd17553,17'd17553,17'd18150,17'd2611,17'd3437,17'd54521,17'd13441,17'd13955,17'd54522,17'd54523,17'd49012,17'd24008,17'd17310,17'd54524,17'd30509,17'd54525,17'd17810,17'd17318,17'd10691,17'd11626,17'd12527,17'd12813,17'd11626,17'd11360,17'd11360,17'd24345,17'd12527,17'd12678,17'd15762,17'd14098,17'd13838,17'd10687,17'd10281,17'd12066,17'd18412,17'd19006,17'd16765,17'd14621,17'd14621,17'd12218,17'd11628,17'd25258,17'd17689,17'd18884,17'd17317,17'd16766,17'd21649,17'd27461,17'd54526,17'd14768,17'd15384,17'd15767,17'd54527,17'd54344,17'd54430,17'd54528,17'd54529,17'd54530,17'd54531,17'd54532,17'd54533,17'd54435,17'd2297,17'd54534,17'd54535,17'd54535,17'd3490,17'd54536,17'd54537,17'd54538,17'd54539,17'd54540,17'd54541,17'd54542,17'd54543,17'd54544,17'd54545,17'd54546,17'd54102,17'd54547,17'd54548,17'd54447,17'd54549,17'd48475,17'd54550,17'd54551,17'd54552,17'd28672,17'd28085,17'd54553,17'd27967,17'd23506,17'd22123,17'd17112,17'd10579,17'd54554,17'd53965,17'd54555,17'd19636,17'd54556,17'd53829,17'd53621,17'd53464,17'd11379,17'd54191,17'd11378,17'd54274,17'd11649,17'd11788,17'd19914,17'd12243,17'd12849,17'd14374,17'd13507,17'd54557,17'd54558,17'd54559,17'd54560,17'd54374,17'd54561,17'd17969,17'd17844,17'd17844,17'd17476,17'd16686,17'd14672,17'd12416,17'd15570,17'd15685,17'd17348,17'd12254,17'd24856,17'd26370,17'd28343,17'd29923,17'd30222,17'd30222,17'd28460,17'd29645,17'd31587,17'd31761,17'd48660,17'd34833,17'd33243,17'd51432,17'd51513,17'd51602,17'd52401,17'd51694,17'd51694,17'd53250,17'd34203,17'd34835,17'd30972,17'd29779,17'd28460,17'd35519,17'd23856,17'd23168,17'd22992,17'd19158,17'd11397,17'd14673,17'd11964,17'd11964,17'd12422,17'd13883,17'd12109,17'd12110,17'd14131,17'd14808,17'd12861,17'd10989,17'd11131,17'd11132,17'd11670,17'd10330,17'd10479,17'd11134,17'd19642,17'd28576,17'd11134,17'd17719,17'd10330,17'd10328,17'd10739,17'd14810,17'd11520,17'd11395,17'd11520,17'd16068,17'd17236,17'd11524,17'd10990,17'd10479,17'd15684,17'd19923,17'd53325,17'd54562,17'd54563,17'd9749,17'd54564,17'd8112,17'd17852,17'd21058,17'd15302,17'd14140,17'd53549,17'd15061,17'd54281,17'd11535,17'd7959,17'd7465,17'd54565,17'd54566,17'd54567,17'd21688,17'd23395,17'd34894,17'd33652,17'd34113,17'd54568,17'd53561,17'd52170,17'd49985,17'd50659,17'd52506,17'd50271,17'd49985,17'd54569,17'd54570,17'd39122,17'd54571,17'd42886,17'd37908,17'd26524,17'd26278,17'd29977,17'd32354,17'd27885,17'd30279,17'd30279,17'd30279,17'd32354,17'd32355,17'd32507,17'd33486,17'd30884,17'd30884,17'd30884,17'd30884,17'd28857,17'd29536,17'd30130,17'd29979,17'd30884,17'd29979,17'd36132,17'd29380,17'd53339,17'd26277,17'd31353,17'd36690,17'd27515,17'd52508,17'd30734,17'd28594,17'd27765,17'd28594,17'd30606,17'd25949,17'd28724,17'd28978,17'd28725,17'd27640,17'd28724,17'd43838,17'd48256,17'd46760,17'd43545,17'd41860,17'd43147,17'd50267,17'd50736,17'd51830,17'd50268,17'd49890,17'd54572,17'd54573,17'd48252,17'd54574,17'd54575,17'd54576,17'd50154,17'd52743,17'd52888,17'd28977,17'd23384,17'd48257,17'd42744,17'd32504,17'd29828,17'd23566,17'd24902,17'd29100,17'd24415,17'd24743,17'd24744,17'd29976,17'd25180,17'd25180,17'd24416,17'd24090,17'd35166,17'd23739,17'd34638,17'd31830,17'd54577,17'd51164,17'd54578,17'd54579,17'd54580,17'd22152,17'd54581,17'd54582,17'd54583,17'd51631,17'd51922,17'd54584,17'd54585,17'd54586,17'd54587,17'd54588,17'd54589,17'd54590,17'd54591,17'd43038,17'd22404,17'd54592,17'd54593,17'd11830,17'd26826,17'd25767,17'd23455,17'd23627,17'd54311,17'd6210,17'd6067,17'd4841,17'd28418,17'd4842,17'd30637,17'd25627,17'd28185,17'd27935,17'd6390,17'd6219,17'd32073,17'd32073,17'd32074,17'd29740,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd29593,17'd29593,17'd31888,17'd31888,17'd27696,17'd7668,17'd6391,17'd5614,17'd31245,17'd30637,17'd5162,17'd37432,17'd4848,17'd34921,17'd49804,17'd49804,17'd40397,17'd29024,17'd5009,17'd5011,17'd50918,17'd54227,17'd52185,17'd53735,17'd54594,17'd44736,17'd54595,17'd54596,17'd54417,17'd54597,17'd54598,17'd54599,17'd54600,17'd54601,17'd54511,17'd54321,17'd54512,17'd54513,17'd54162,17'd54602,17'd52916,17'd54603,17'd40410,17'd6236,17'd6084,17'd18144,17'd448,17'd628,17'd4059,17'd52698,17'd54326,17'd52615,17'd1402,17'd2410,17'd54604,17'd630,17'd37043,17'd37043,17'd236,17'd448,17'd628,17'd4059,17'd1824,17'd1824,17'd4398,17'd4398,17'd3390,17'd54516,17'd54327,17'd35058,17'd54517,17'd54329,17'd54518,17'd54605,17'd54606,17'd2086,17'd54165,17'd54607
},
'{
17'd16010,17'd10925,17'd10670,17'd10669,17'd52621,17'd2426,17'd1414,17'd1416,17'd653,17'd653,17'd980,17'd980,17'd27,17'd27,17'd285,17'd285,17'd285,17'd285,17'd285,17'd285,17'd286,17'd27,17'd4430,17'd4430,17'd4091,17'd3755,17'd3255,17'd2940,17'd2602,17'd2600,17'd22615,17'd1838,17'd2121,17'd1557,17'd1137,17'd19244,17'd19244,17'd17553,17'd2787,17'd1979,17'd54608,17'd23660,17'd38337,17'd54609,17'd54610,17'd14607,17'd24340,17'd16154,17'd54611,17'd47672,17'd54525,17'd17810,17'd54612,17'd10427,17'd23154,17'd12813,17'd12813,17'd11626,17'd11360,17'd11360,17'd12065,17'd12679,17'd13092,17'd13597,17'd13716,17'd12355,17'd10687,17'd10281,17'd11229,17'd18412,17'd19382,17'd16658,17'd12361,17'd12361,17'd12362,17'd11764,17'd25258,17'd19753,17'd19006,17'd17317,17'd16766,17'd21649,17'd19007,17'd17320,17'd14768,17'd47972,17'd15767,17'd54527,17'd54613,17'd54614,17'd54615,17'd54616,17'd54617,17'd54618,17'd54347,17'd54619,17'd54620,17'd2297,17'd2158,17'd54621,17'd54622,17'd3000,17'd54623,17'd54624,17'd54625,17'd54626,17'd54627,17'd54628,17'd54629,17'd54630,17'd54182,17'd54545,17'd54631,17'd54632,17'd54633,17'd54634,17'd54635,17'd53763,17'd54636,17'd54637,17'd54638,17'd54639,17'd29766,17'd27723,17'd54640,17'd25918,17'd24690,17'd52211,17'd52291,17'd16539,17'd10710,17'd10445,17'd10711,17'd54641,17'd13872,17'd13239,17'd53464,17'd53180,17'd53384,17'd11502,17'd24985,17'd54642,17'd11648,17'd16901,17'd12243,17'd12243,17'd12400,17'd12849,17'd13359,17'd21358,17'd21201,17'd54643,17'd54644,17'd54645,17'd54278,17'd18331,17'd17969,17'd19031,17'd19031,17'd17013,17'd15571,17'd14930,17'd13517,17'd13252,17'd16321,17'd12579,17'd23855,17'd28107,17'd28227,17'd28943,17'd28943,17'd28943,17'd28943,17'd29066,17'd28686,17'd31587,17'd31289,17'd33568,17'd34833,17'd36936,17'd51603,17'd52134,17'd51602,17'd51694,17'd51694,17'd34705,17'd34037,17'd31289,17'd30974,17'd30074,17'd28461,17'd28230,17'd23856,17'd24030,17'd24362,17'd16442,17'd11396,17'd14673,17'd14673,17'd11964,17'd17604,17'd13135,17'd13761,17'd13882,17'd12577,17'd30682,17'd13363,17'd13762,17'd10854,17'd11132,17'd11670,17'd10330,17'd11276,17'd11276,17'd16070,17'd48579,17'd16070,17'd16796,17'd10330,17'd10328,17'd10475,17'd14931,17'd11395,17'd11395,17'd11520,17'd11395,17'd14673,17'd17236,17'd14931,17'd20756,17'd10174,17'd9887,17'd16690,17'd54646,17'd54647,17'd18924,17'd54648,17'd8263,17'd24552,17'd54381,17'd21058,17'd14140,17'd15437,17'd20320,17'd54649,17'd54650,17'd14142,17'd54651,17'd54652,17'd54653,17'd54654,17'd22318,17'd22505,17'd50733,17'd33482,17'd54655,17'd54656,17'd49483,17'd51077,17'd50273,17'd42142,17'd54657,17'd50370,17'd50271,17'd54658,17'd43419,17'd54659,17'd48697,17'd32826,17'd30279,17'd28980,17'd27642,17'd30279,17'd27885,17'd27885,17'd30279,17'd27885,17'd27885,17'd32354,17'd32017,17'd28372,17'd29106,17'd30884,17'd29691,17'd29691,17'd30884,17'd29536,17'd29831,17'd31038,17'd28857,17'd29536,17'd29831,17'd28372,17'd28856,17'd28854,17'd47633,17'd38025,17'd27258,17'd27767,17'd33507,17'd28598,17'd28594,17'd28594,17'd27638,17'd28602,17'd25833,17'd28724,17'd28724,17'd27515,17'd26530,17'd35012,17'd42885,17'd48698,17'd46954,17'd54660,17'd47343,17'd49093,17'd50164,17'd50736,17'd50371,17'd50736,17'd49692,17'd54661,17'd48353,17'd48033,17'd51555,17'd53203,17'd53333,17'd53262,17'd54135,17'd53720,17'd34467,17'd28976,17'd29975,17'd37117,17'd38976,17'd23923,17'd29242,17'd23731,17'd24415,17'd29100,17'd24252,17'd25030,17'd27637,17'd25178,17'd25179,17'd24743,17'd23917,17'd35166,17'd45614,17'd40523,17'd54662,17'd48269,17'd46862,17'd54209,17'd51298,17'd52514,17'd29725,17'd54663,17'd54664,17'd51067,17'd51067,17'd51748,17'd54299,17'd54665,17'd54666,17'd54667,17'd54668,17'd35184,17'd54669,17'd22554,17'd54670,17'd53730,17'd54671,17'd25877,17'd54672,17'd11158,17'd24644,17'd24307,17'd23627,17'd54497,17'd24795,17'd4995,17'd4841,17'd28418,17'd4842,17'd5004,17'd25627,17'd28185,17'd27935,17'd6390,17'd6390,17'd32073,17'd9091,17'd29740,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd31888,17'd31888,17'd29593,17'd29593,17'd31888,17'd31888,17'd27696,17'd7668,17'd6220,17'd27935,17'd30796,17'd4842,17'd4847,17'd28778,17'd5157,17'd4846,17'd54673,17'd49804,17'd4527,17'd51176,17'd38059,17'd4850,17'd51931,17'd38446,17'd54674,17'd47478,17'd54675,17'd54676,17'd54677,17'd54678,17'd54679,17'd54680,17'd54681,17'd54682,17'd54683,17'd54684,17'd54685,17'd54686,17'd54512,17'd54513,17'd54162,17'd50923,17'd52193,17'd3867,17'd6082,17'd54687,17'd7341,17'd18144,17'd448,17'd629,17'd628,17'd52698,17'd2113,17'd795,17'd8015,17'd8015,17'd629,17'd236,17'd54688,17'd36902,17'd630,17'd448,17'd447,17'd2587,17'd3072,17'd1824,17'd2558,17'd38071,17'd3390,17'd54689,17'd54690,17'd35206,17'd54328,17'd53155,17'd54518,17'd54691,17'd54692,17'd53597,17'd54520,17'd54607
},
'{
17'd16010,17'd10925,17'd10670,17'd10669,17'd52621,17'd52621,17'd2596,17'd1414,17'd468,17'd653,17'd652,17'd980,17'd980,17'd27,17'd26,17'd285,17'd285,17'd285,17'd285,17'd285,17'd286,17'd27,17'd6744,17'd4430,17'd4091,17'd3755,17'd3255,17'd2941,17'd2602,17'd2600,17'd22615,17'd1838,17'd2121,17'd1282,17'd1137,17'd824,17'd824,17'd824,17'd827,17'd2437,17'd54693,17'd32732,17'd38868,17'd41163,17'd54694,17'd54695,17'd54696,17'd13702,17'd54697,17'd54698,17'd32415,17'd18175,17'd46889,17'd10564,17'd12957,17'd12813,17'd12813,17'd17096,17'd24347,17'd12815,17'd13211,17'd13093,17'd13092,17'd12678,17'd13597,17'd12355,17'd10687,17'd10281,17'd9572,17'd11230,17'd32261,17'd19006,17'd12532,17'd12361,17'd12680,17'd11764,17'd54699,17'd25258,17'd19006,17'd17317,17'd19893,17'd16766,17'd21649,17'd17320,17'd15384,17'd47972,17'd15767,17'd32100,17'd54613,17'd54700,17'd54701,17'd54702,17'd54703,17'd54704,17'd54705,17'd54706,17'd54707,17'd3482,17'd3309,17'd54621,17'd54708,17'd2664,17'd3314,17'd54709,17'd54710,17'd54711,17'd54712,17'd54713,17'd54714,17'd54715,17'd53090,17'd54632,17'd54716,17'd54546,17'd54717,17'd54718,17'd54719,17'd53763,17'd54720,17'd54721,17'd54722,17'd54551,17'd54451,17'd27606,17'd51782,17'd50600,17'd24690,17'd54723,17'd54724,17'd54725,17'd18551,17'd54726,17'd54188,17'd54555,17'd23160,17'd12982,17'd54456,17'd53241,17'd11380,17'd53771,17'd13239,17'd14506,17'd54727,17'd54728,17'd20304,17'd12093,17'd12568,17'd12849,17'd14374,17'd21980,17'd22126,17'd54729,17'd54372,17'd54730,17'd54731,17'd18199,17'd18331,17'd19031,17'd19031,17'd17013,17'd17235,17'd15687,17'd12418,17'd12995,17'd16321,17'd14807,17'd12255,17'd28107,17'd28227,17'd28943,17'd29066,17'd29066,17'd28943,17'd28943,17'd28818,17'd31768,17'd30974,17'd34381,17'd54732,17'd34833,17'd53250,17'd51603,17'd51602,17'd51602,17'd51694,17'd51603,17'd35644,17'd34203,17'd34381,17'd30974,17'd29330,17'd29480,17'd40597,17'd24537,17'd24992,17'd16325,17'd11522,17'd14673,17'd14673,17'd14673,17'd11964,17'd12996,17'd13883,17'd13761,17'd12577,17'd12413,17'd13761,17'd13253,17'd14931,17'd19282,17'd11670,17'd10330,17'd11671,17'd11671,17'd14928,17'd25530,17'd25530,17'd9885,17'd11134,17'd10167,17'd19282,17'd16320,17'd14931,17'd14262,17'd11520,17'd16068,17'd11523,17'd11523,17'd14810,17'd26037,17'd17716,17'd11404,17'd24044,17'd48212,17'd19783,17'd54733,17'd54734,17'd54735,17'd10748,17'd54736,17'd19288,17'd19288,17'd10862,17'd54737,17'd7960,17'd54738,17'd8587,17'd54739,17'd54740,17'd54741,17'd54742,17'd36544,17'd22502,17'd30578,17'd54743,17'd54744,17'd54745,17'd48262,17'd54746,17'd42875,17'd42142,17'd50475,17'd54657,17'd54747,17'd49389,17'd49278,17'd47052,17'd42599,17'd39437,17'd40681,17'd29379,17'd27642,17'd27642,17'd30279,17'd29977,17'd29977,17'd27885,17'd28134,17'd32192,17'd32017,17'd28372,17'd29106,17'd29691,17'd29691,17'd53122,17'd29691,17'd29536,17'd36132,17'd29831,17'd29536,17'd29831,17'd28372,17'd29105,17'd29104,17'd28255,17'd26525,17'd35011,17'd25949,17'd31055,17'd28599,17'd28598,17'd27638,17'd28594,17'd30606,17'd25833,17'd28252,17'd28724,17'd27515,17'd26530,17'd28602,17'd43978,17'd52343,17'd49978,17'd54748,17'd48609,17'd47641,17'd49478,17'd50365,17'd50272,17'd50272,17'd49890,17'd45150,17'd54749,17'd54750,17'd54059,17'd54290,17'd54751,17'd53333,17'd53563,17'd48695,17'd34276,17'd24902,17'd29687,17'd36987,17'd29973,17'd37117,17'd29242,17'd28849,17'd34467,17'd23916,17'd29100,17'd24252,17'd29976,17'd27637,17'd25178,17'd25179,17'd24743,17'd23917,17'd42449,17'd32363,17'd34882,17'd32665,17'd52986,17'd54752,17'd54753,17'd54754,17'd51903,17'd54755,17'd54663,17'd54664,17'd51563,17'd51563,17'd47163,17'd54756,17'd54757,17'd54758,17'd54759,17'd54760,17'd54761,17'd20817,17'd54762,17'd54763,17'd22750,17'd30329,17'd25360,17'd54672,17'd23628,17'd54764,17'd24307,17'd6839,17'd6210,17'd5322,17'd4840,17'd4686,17'd28418,17'd4842,17'd5004,17'd25627,17'd28185,17'd27935,17'd6390,17'd6390,17'd32073,17'd9091,17'd29740,17'd27696,17'd27696,17'd27696,17'd27696,17'd27696,17'd31888,17'd31888,17'd29593,17'd29593,17'd31888,17'd31888,17'd27696,17'd7668,17'd6390,17'd5160,17'd31716,17'd28536,17'd28778,17'd34791,17'd4846,17'd5156,17'd54765,17'd49804,17'd4527,17'd51176,17'd5007,17'd54498,17'd49997,17'd38706,17'd54766,17'd37566,17'd54767,17'd43873,17'd54768,17'd54769,17'd54680,17'd54770,17'd54508,17'd54771,17'd54772,17'd54773,17'd54774,17'd54686,17'd54775,17'd54513,17'd54162,17'd53744,17'd52019,17'd3867,17'd6082,17'd54776,17'd54777,17'd18144,17'd448,17'd448,17'd796,17'd54778,17'd1264,17'd1402,17'd8015,17'd3248,17'd235,17'd797,17'd54688,17'd36902,17'd235,17'd629,17'd2587,17'd1402,17'd1824,17'd1824,17'd2558,17'd4228,17'd54779,17'd54780,17'd54781,17'd1663,17'd54782,17'd54783,17'd54518,17'd54784,17'd54785,17'd2086,17'd54786,17'd53599
},
'{
17'd16010,17'd10924,17'd10670,17'd10669,17'd52621,17'd2426,17'd2257,17'd2257,17'd1416,17'd4089,17'd653,17'd652,17'd980,17'd27,17'd27,17'd286,17'd285,17'd285,17'd285,17'd285,17'd286,17'd27,17'd6744,17'd4430,17'd4091,17'd4091,17'd3595,17'd2941,17'd2602,17'd2600,17'd22615,17'd22615,17'd16966,17'd1282,17'd991,17'd992,17'd824,17'd825,17'd826,17'd828,17'd54787,17'd54788,17'd54789,17'd29307,17'd54790,17'd54791,17'd54792,17'd54793,17'd54794,17'd54795,17'd54796,17'd18175,17'd48297,17'd30356,17'd12680,17'd23154,17'd12813,17'd13093,17'd23154,17'd12815,17'd13211,17'd13093,17'd12527,17'd12678,17'd13462,17'd12062,17'd11762,17'd11086,17'd10814,17'd12066,17'd27218,17'd19382,17'd18884,17'd12531,17'd12680,17'd11913,17'd27218,17'd25258,17'd17941,17'd19893,17'd17204,17'd17689,17'd21649,17'd15899,17'd15384,17'd47972,17'd15641,17'd32101,17'd54797,17'd54798,17'd54799,17'd54800,17'd54801,17'd54802,17'd54803,17'd54804,17'd54253,17'd54805,17'd1873,17'd54621,17'd54806,17'd2483,17'd54807,17'd54808,17'd5855,17'd54809,17'd54810,17'd54811,17'd54812,17'd54813,17'd42508,17'd54814,17'd54716,17'd54815,17'd54816,17'd54817,17'd54818,17'd47388,17'd54819,17'd54271,17'd54637,17'd54638,17'd30060,17'd27466,17'd27222,17'd54640,17'd54820,17'd50403,17'd51593,17'd17829,17'd10444,17'd18551,17'd15665,17'd10711,17'd21975,17'd14919,17'd11502,17'd11380,17'd53241,17'd53385,17'd53969,17'd14506,17'd12395,17'd12395,17'd12237,17'd12089,17'd20304,17'd12849,17'd12400,17'd13247,17'd54371,17'd23675,17'd54821,17'd54822,17'd54823,17'd54824,17'd45933,17'd54825,17'd18685,17'd17726,17'd17724,17'd16560,17'd16799,17'd14809,17'd13252,17'd15570,17'd12108,17'd24991,17'd28343,17'd28943,17'd29066,17'd30071,17'd28943,17'd29923,17'd28227,17'd28345,17'd29198,17'd30677,17'd31289,17'd34203,17'd54376,17'd54826,17'd53630,17'd51693,17'd51602,17'd51513,17'd51432,17'd33243,17'd33568,17'd34835,17'd30677,17'd28686,17'd30524,17'd24856,17'd24208,17'd24995,17'd14264,17'd14673,17'd14673,17'd16068,17'd11395,17'd13762,17'd13135,17'd13761,17'd12414,17'd12414,17'd14130,17'd15299,17'd16068,17'd11132,17'd12863,17'd10330,17'd11671,17'd11671,17'd12116,17'd26759,17'd26759,17'd10992,17'd9883,17'd10167,17'd19532,17'd10739,17'd10990,17'd14810,17'd11519,17'd14262,17'd14673,17'd11523,17'd13138,17'd21205,17'd16065,17'd12264,17'd13375,17'd9051,17'd24373,17'd54827,17'd19538,17'd8264,17'd21825,17'd54828,17'd13654,17'd19646,17'd54829,17'd12430,17'd54830,17'd54831,17'd18207,17'd54832,17'd54833,17'd54834,17'd54835,17'd22507,17'd24421,17'd29375,17'd54836,17'd54837,17'd54838,17'd48995,17'd50474,17'd50475,17'd42142,17'd50475,17'd54389,17'd54839,17'd40206,17'd46946,17'd43975,17'd36690,17'd27642,17'd33952,17'd30279,17'd29977,17'd27642,17'd29379,17'd28980,17'd28980,17'd26276,17'd27884,17'd28370,17'd28257,17'd29380,17'd28372,17'd29106,17'd31196,17'd31196,17'd29106,17'd29537,17'd49286,17'd29537,17'd36848,17'd28728,17'd29105,17'd53339,17'd26522,17'd27642,17'd30586,17'd26903,17'd27513,17'd33000,17'd25567,17'd25567,17'd27638,17'd30606,17'd26062,17'd25707,17'd28724,17'd27515,17'd28482,17'd28481,17'd28723,17'd43425,17'd54840,17'd50902,17'd48522,17'd47828,17'd43281,17'd50267,17'd50568,17'd50476,17'd50574,17'd49693,17'd54841,17'd54842,17'd54843,17'd54844,17'd54205,17'd54845,17'd50068,17'd50154,17'd53557,17'd23916,17'd29689,17'd29830,17'd38976,17'd29973,17'd32191,17'd23564,17'd29100,17'd32659,17'd23916,17'd24090,17'd24742,17'd25178,17'd25568,17'd25177,17'd25030,17'd24742,17'd24087,17'd54846,17'd45614,17'd34759,17'd32997,17'd51479,17'd53344,17'd54847,17'd54848,17'd54849,17'd53655,17'd47749,17'd54583,17'd51394,17'd54664,17'd54850,17'd54851,17'd54852,17'd54853,17'd54854,17'd54855,17'd54856,17'd54857,17'd54858,17'd54859,17'd22750,17'd54860,17'd25483,17'd26583,17'd24793,17'd54764,17'd23627,17'd23974,17'd24148,17'd5323,17'd32552,17'd4686,17'd28418,17'd5005,17'd5004,17'd25627,17'd28185,17'd27935,17'd6390,17'd6554,17'd9091,17'd7499,17'd27696,17'd27696,17'd27696,17'd27696,17'd31888,17'd31888,17'd31888,17'd31888,17'd29593,17'd31888,17'd27696,17'd29740,17'd7499,17'd6391,17'd30638,17'd5004,17'd28536,17'd5327,17'd54861,17'd4526,17'd4689,17'd5155,17'd54765,17'd54862,17'd49995,17'd50586,17'd50835,17'd54003,17'd51489,17'd54500,17'd46987,17'd54863,17'd39784,17'd54864,17'd54865,17'd54866,17'd54867,17'd54868,17'd54869,17'd54870,17'd54010,17'd54773,17'd54871,17'd54872,17'd54873,17'd54874,17'd41312,17'd38456,17'd54875,17'd54876,17'd6082,17'd54776,17'd54777,17'd38856,17'd448,17'd448,17'd1121,17'd1121,17'd1264,17'd3072,17'd5775,17'd628,17'd630,17'd239,17'd449,17'd243,17'd448,17'd629,17'd2587,17'd1402,17'd3898,17'd1824,17'd2558,17'd38071,17'd53151,17'd54877,17'd54878,17'd1663,17'd54879,17'd53296,17'd53677,17'd54784,17'd24494,17'd2086,17'd54786,17'd53751
},
'{
17'd11609,17'd10924,17'd10670,17'd10669,17'd52621,17'd10547,17'd2597,17'd2257,17'd1416,17'd1416,17'd653,17'd652,17'd980,17'd980,17'd27,17'd286,17'd285,17'd285,17'd285,17'd285,17'd286,17'd27,17'd6744,17'd4430,17'd4091,17'd3755,17'd3255,17'd2941,17'd2602,17'd2600,17'd22615,17'd23658,17'd16966,17'd19499,17'd992,17'd992,17'd825,17'd825,17'd826,17'd828,17'd54787,17'd54880,17'd2795,17'd22970,17'd54881,17'd54882,17'd49410,17'd49715,17'd54883,17'd54884,17'd54796,17'd18175,17'd16169,17'd10693,17'd10815,17'd13094,17'd34938,17'd12813,17'd23154,17'd12815,17'd13211,17'd17096,17'd12813,17'd15516,17'd14469,17'd12062,17'd11762,17'd11086,17'd10108,17'd12066,17'd27218,17'd19753,17'd17204,17'd18884,17'd43599,17'd12680,17'd27218,17'd54885,17'd18774,17'd19893,17'd19382,17'd17689,17'd21649,17'd15899,17'd15384,17'd33548,17'd14893,17'd24194,17'd54886,17'd54887,17'd54888,17'd54889,17'd54890,17'd54891,17'd54892,17'd54893,17'd54894,17'd54895,17'd54896,17'd54897,17'd54898,17'd54899,17'd2666,17'd54900,17'd54901,17'd54902,17'd54903,17'd54904,17'd54905,17'd54906,17'd54907,17'd54908,17'd54546,17'd54815,17'd54909,17'd54910,17'd54911,17'd42217,17'd54912,17'd54913,17'd54914,17'd54915,17'd54916,17'd51189,17'd50684,17'd51782,17'd28086,17'd54917,17'd50854,17'd54918,17'd17829,17'd10444,17'd16784,17'd10959,17'd10960,17'd54919,17'd54642,17'd53384,17'd53241,17'd53180,17'd54369,17'd54642,17'd11647,17'd54920,17'd13238,17'd11649,17'd20304,17'd18799,17'd13996,17'd12567,17'd54111,17'd54921,17'd23675,17'd54922,17'd54923,17'd54924,17'd54561,17'd18331,17'd18685,17'd28232,17'd17724,17'd17013,17'd14524,17'd13643,17'd15570,17'd15433,17'd12108,17'd24991,17'd28343,17'd28943,17'd30071,17'd29329,17'd30831,17'd30218,17'd28343,17'd27984,17'd28686,17'd30974,17'd54925,17'd31288,17'd54926,17'd54927,17'd34556,17'd51602,17'd51602,17'd51602,17'd51513,17'd53250,17'd33720,17'd34203,17'd34835,17'd30220,17'd51601,17'd27346,17'd24857,17'd24362,17'd14259,17'd11397,17'd11274,17'd12720,17'd11395,17'd11964,17'd12996,17'd13761,17'd12414,17'd12109,17'd14130,17'd15054,17'd16069,17'd21206,17'd11400,17'd10330,17'd11671,17'd11671,17'd12116,17'd16070,17'd26759,17'd13255,17'd9884,17'd21503,17'd10330,17'd10476,17'd11399,17'd14931,17'd14931,17'd10990,17'd11397,17'd12583,17'd13138,17'd26630,17'd33083,17'd8725,17'd50418,17'd11140,17'd54928,17'd54929,17'd17854,17'd19538,17'd19784,17'd22481,17'd54930,17'd19419,17'd10343,17'd13771,17'd54931,17'd17854,17'd20323,17'd54932,17'd54933,17'd54934,17'd54935,17'd22680,17'd29527,17'd30431,17'd54936,17'd54937,17'd44929,17'd49478,17'd50474,17'd54569,17'd42142,17'd42142,17'd50573,17'd54572,17'd52340,17'd46556,17'd45878,17'd31353,17'd29246,17'd29977,17'd40681,17'd33952,17'd31353,17'd29245,17'd28726,17'd44703,17'd26277,17'd27884,17'd28133,17'd28371,17'd30587,17'd29380,17'd28372,17'd29106,17'd31196,17'd28372,17'd29537,17'd49285,17'd52429,17'd52429,17'd29104,17'd53339,17'd26522,17'd26523,17'd26781,17'd28725,17'd40965,17'd28599,17'd33000,17'd28369,17'd27765,17'd28598,17'd30606,17'd25949,17'd26903,17'd26903,17'd28482,17'd40965,17'd30606,17'd28721,17'd50153,17'd54938,17'd54939,17'd39736,17'd47446,17'd48363,17'd49794,17'd50568,17'd50907,17'd54747,17'd49389,17'd46656,17'd54940,17'd54941,17'd51387,17'd54942,17'd54480,17'd52343,17'd48695,17'd40964,17'd28722,17'd23385,17'd29975,17'd38976,17'd23216,17'd23387,17'd28849,17'd24252,17'd28851,17'd34467,17'd24415,17'd24744,17'd27512,17'd25709,17'd25177,17'd28974,17'd28851,17'd24087,17'd54943,17'd34277,17'd30581,17'd22864,17'd51067,17'd51384,17'd54944,17'd54945,17'd54946,17'd30164,17'd54947,17'd47652,17'd46775,17'd46862,17'd54948,17'd54949,17'd54950,17'd54951,17'd54952,17'd35326,17'd26210,17'd54953,17'd54954,17'd22058,17'd54955,17'd30484,17'd12135,17'd54956,17'd54957,17'd54958,17'd23457,17'd23974,17'd24148,17'd5323,17'd4688,17'd4841,17'd28418,17'd5005,17'd5004,17'd25627,17'd28185,17'd27935,17'd6390,17'd6554,17'd9091,17'd7499,17'd27696,17'd27696,17'd27696,17'd27696,17'd31888,17'd31888,17'd31888,17'd31888,17'd31888,17'd31888,17'd27696,17'd29740,17'd7499,17'd6220,17'd30333,17'd5005,17'd5328,17'd47174,17'd54959,17'd5156,17'd4689,17'd49804,17'd54960,17'd54961,17'd39015,17'd4528,17'd50835,17'd52011,17'd49599,17'd51094,17'd54962,17'd54963,17'd44736,17'd54964,17'd54965,17'd54966,17'd54967,17'd54968,17'd54969,17'd54970,17'd54971,17'd54972,17'd54871,17'd54872,17'd54973,17'd54874,17'd41312,17'd54974,17'd51252,17'd54876,17'd54975,17'd54877,17'd54689,17'd38856,17'd448,17'd448,17'd1121,17'd1121,17'd795,17'd3745,17'd5775,17'd796,17'd236,17'd239,17'd239,17'd243,17'd629,17'd628,17'd795,17'd3072,17'd3898,17'd3898,17'd2558,17'd4228,17'd6406,17'd54877,17'd54878,17'd19361,17'd54879,17'd53365,17'd53677,17'd54976,17'd24494,17'd54977,17'd54786,17'd53751
},
'{
17'd54978,17'd54978,17'd10802,17'd10669,17'd10547,17'd52621,17'd2597,17'd1414,17'd1416,17'd16,17'd18,17'd3905,17'd28,17'd652,17'd1278,17'd27,17'd467,17'd285,17'd285,17'd285,17'd286,17'd27,17'd6744,17'd4430,17'd4431,17'd4431,17'd3595,17'd2941,17'd2601,17'd2263,17'd2600,17'd54979,17'd1282,17'd19499,17'd992,17'd827,17'd57,17'd57,17'd827,17'd18275,17'd41628,17'd39038,17'd2620,17'd34932,17'd27101,17'd54980,17'd54981,17'd54696,17'd54982,17'd54983,17'd54984,17'd54985,17'd16411,17'd29905,17'd11629,17'd13094,17'd34938,17'd11626,17'd23154,17'd13094,17'd12815,17'd13094,17'd11626,17'd12527,17'd15516,17'd15516,17'd11762,17'd11086,17'd10108,17'd12956,17'd18412,17'd54885,17'd17689,17'd19893,17'd10815,17'd14472,17'd12681,17'd48930,17'd18655,17'd19893,17'd19006,17'd20422,17'd21649,17'd16028,17'd14768,17'd15519,17'd15520,17'd32101,17'd54986,17'd54344,17'd54987,17'd54988,17'd54989,17'd54990,17'd54991,17'd54992,17'd54993,17'd54618,17'd1872,17'd54994,17'd54995,17'd54996,17'd54997,17'd54998,17'd54999,17'd55000,17'd55001,17'd55002,17'd55003,17'd55004,17'd55005,17'd55006,17'd55007,17'd54815,17'd55008,17'd55009,17'd55010,17'd54718,17'd55011,17'd55012,17'd55013,17'd55014,17'd55015,17'd50939,17'd50940,17'd27110,17'd27724,17'd55016,17'd51109,17'd52211,17'd17112,17'd16897,17'd55017,17'd54453,17'd10711,17'd21975,17'd16195,17'd53970,17'd55018,17'd53180,17'd55019,17'd55020,17'd54920,17'd55021,17'd54727,17'd12091,17'd15172,17'd20304,17'd14373,17'd14373,17'd13247,17'd55022,17'd54921,17'd55023,17'd55024,17'd55025,17'd55026,17'd45814,17'd18685,17'd37738,17'd18685,17'd19031,17'd17014,17'd44647,17'd14526,17'd15433,17'd19407,17'd18200,17'd27121,17'd30222,17'd30370,17'd31940,17'd30071,17'd29923,17'd28816,17'd28816,17'd28461,17'd31440,17'd31767,17'd33409,17'd33721,17'd34545,17'd54826,17'd53630,17'd52302,17'd51602,17'd51694,17'd51513,17'd53250,17'd34833,17'd54732,17'd30677,17'd28686,17'd28103,17'd24859,17'd24992,17'd28112,17'd11396,17'd11274,17'd14810,17'd11520,17'd11964,17'd16204,17'd13883,17'd12109,17'd12414,17'd12579,17'd13882,17'd16064,17'd14931,17'd19282,17'd10330,17'd11671,17'd9884,17'd15566,17'd16549,17'd32916,17'd17011,17'd9885,17'd16796,17'd10330,17'd14518,17'd11132,17'd16320,17'd16320,17'd14931,17'd11397,17'd19533,17'd17838,17'd21205,17'd50112,17'd20176,17'd16072,17'd55027,17'd20049,17'd55028,17'd55029,17'd54463,17'd10612,17'd24371,17'd20049,17'd13528,17'd13259,17'd21510,17'd7467,17'd55030,17'd55031,17'd55032,17'd55033,17'd55034,17'd55035,17'd32008,17'd45763,17'd55036,17'd55037,17'd55038,17'd43281,17'd54839,17'd54747,17'd54389,17'd42142,17'd42873,17'd55039,17'd40951,17'd46844,17'd43834,17'd36542,17'd29379,17'd31353,17'd31352,17'd40681,17'd33952,17'd27368,17'd25945,17'd26898,17'd25557,17'd26652,17'd27761,17'd28854,17'd28370,17'd28257,17'd28257,17'd29247,17'd29247,17'd29104,17'd29247,17'd28371,17'd52429,17'd33320,17'd32354,17'd40681,17'd29977,17'd27642,17'd28979,17'd35578,17'd55040,17'd38671,17'd28597,17'd27882,17'd28369,17'd25567,17'd27638,17'd28602,17'd26174,17'd27515,17'd26530,17'd27767,17'd27767,17'd28598,17'd44229,17'd55041,17'd54290,17'd47732,17'd47735,17'd47937,17'd49184,17'd49980,17'd50271,17'd54747,17'd49988,17'd55042,17'd55043,17'd55044,17'd55045,17'd50901,17'd50361,17'd53333,17'd52817,17'd50155,17'd34467,17'd29972,17'd29827,17'd29975,17'd37117,17'd23388,17'd23566,17'd23916,17'd24745,17'd24416,17'd24743,17'd24252,17'd25032,17'd25177,17'd25709,17'd25438,17'd24898,17'd35159,17'd23732,17'd55046,17'd44110,17'd33945,17'd33946,17'd55047,17'd55048,17'd55049,17'd55050,17'd21999,17'd51562,17'd51817,17'd51067,17'd21703,17'd53852,17'd55051,17'd55052,17'd55053,17'd54759,17'd55054,17'd55055,17'd55056,17'd22555,17'd55057,17'd55058,17'd22565,17'd55059,17'd12135,17'd55060,17'd23453,17'd23455,17'd23457,17'd6840,17'd4680,17'd5607,17'd32552,17'd5328,17'd5002,17'd4842,17'd30637,17'd5335,17'd5614,17'd27935,17'd31717,17'd6554,17'd7499,17'd7668,17'd27696,17'd27696,17'd31888,17'd31888,17'd31888,17'd29593,17'd29593,17'd31888,17'd29593,17'd31888,17'd29740,17'd29740,17'd7668,17'd5615,17'd25627,17'd4842,17'd4684,17'd54861,17'd41891,17'd44614,17'd55061,17'd54765,17'd4369,17'd4369,17'd49896,17'd50918,17'd54003,17'd51403,17'd54004,17'd55062,17'd55063,17'd55064,17'd55065,17'd55066,17'd55067,17'd55068,17'd55069,17'd54770,17'd55070,17'd54772,17'd55071,17'd55072,17'd55073,17'd55074,17'd54973,17'd55075,17'd39027,17'd55076,17'd51251,17'd55077,17'd55078,17'd55079,17'd3071,17'd1121,17'd448,17'd235,17'd447,17'd2587,17'd1402,17'd3072,17'd1944,17'd235,17'd449,17'd450,17'd238,17'd242,17'd234,17'd2587,17'd626,17'd625,17'd11590,17'd3898,17'd4398,17'd628,17'd3071,17'd55080,17'd55081,17'd19238,17'd55082,17'd53365,17'd55083,17'd55084,17'd24494,17'd2086,17'd54786,17'd53366
},
'{
17'd54978,17'd54978,17'd10802,17'd10669,17'd10547,17'd52621,17'd2597,17'd2596,17'd2257,17'd17,17'd17,17'd3905,17'd652,17'd652,17'd1278,17'd27,17'd467,17'd285,17'd285,17'd285,17'd286,17'd286,17'd6744,17'd4430,17'd4431,17'd4431,17'd3595,17'd2941,17'd2601,17'd2263,17'd2600,17'd55085,17'd1134,17'd19609,17'd827,17'd481,17'd59,17'd56,17'd667,17'd18275,17'd41628,17'd2950,17'd55086,17'd2796,17'd27325,17'd48472,17'd55087,17'd54792,17'd16757,17'd55088,17'd33061,17'd54985,17'd24192,17'd16767,17'd11087,17'd12956,17'd10814,17'd11626,17'd23154,17'd13094,17'd12815,17'd13094,17'd11626,17'd11476,17'd10941,17'd15516,17'd11762,17'd11625,17'd10941,17'd11360,17'd18412,17'd19891,17'd16986,17'd21964,17'd19621,17'd10815,17'd12681,17'd32102,17'd19511,17'd27834,17'd19006,17'd20422,17'd21649,17'd16028,17'd14346,17'd15519,17'd24194,17'd32101,17'd34177,17'd54613,17'd54993,17'd55089,17'd55090,17'd55091,17'd55092,17'd55093,17'd54893,17'd54895,17'd55094,17'd55095,17'd55096,17'd55097,17'd55098,17'd55099,17'd55100,17'd5552,17'd54999,17'd55101,17'd55102,17'd55103,17'd55104,17'd53091,17'd55105,17'd55106,17'd55107,17'd55108,17'd55109,17'd55110,17'd55111,17'd55011,17'd55112,17'd55113,17'd55114,17'd55115,17'd55116,17'd27109,17'd27332,17'd55117,17'd51873,17'd21811,17'd19770,17'd17112,17'd55118,17'd10710,17'd10959,17'd10960,17'd54109,17'd14506,17'd53621,17'd53180,17'd55119,17'd53970,17'd21496,17'd54920,17'd14506,17'd11648,17'd15172,17'd20304,17'd14373,17'd14373,17'd13129,17'd22293,17'd23676,17'd55120,17'd55121,17'd55122,17'd55123,17'd45933,17'd19031,17'd17725,17'd18685,17'd19031,17'd19031,17'd16686,17'd21057,17'd51039,17'd13515,17'd23855,17'd27121,17'd30222,17'd30071,17'd31940,17'd30370,17'd29066,17'd28816,17'd40597,17'd29480,17'd29330,17'd33884,17'd33727,17'd33721,17'd35644,17'd34556,17'd53394,17'd52401,17'd52401,17'd51694,17'd51694,17'd34705,17'd54376,17'd54926,17'd34385,17'd30220,17'd29480,17'd27346,17'd24030,17'd24995,17'd17478,17'd11274,17'd14673,17'd11395,17'd14262,17'd13362,17'd11806,17'd12110,17'd12414,17'd12579,17'd15184,17'd13764,17'd14810,17'd11669,17'd24996,17'd10329,17'd9884,17'd15566,17'd16549,17'd24998,17'd9479,17'd9741,17'd9741,17'd11276,17'd11527,17'd15176,17'd13886,17'd13886,17'd14931,17'd11397,17'd19533,17'd13138,17'd26037,17'd51790,17'd26874,17'd8580,17'd55124,17'd19647,17'd18922,17'd54827,17'd55125,17'd14014,17'd54051,17'd55126,17'd16079,17'd24047,17'd17732,17'd17855,17'd55127,17'd55128,17'd55129,17'd55130,17'd55131,17'd55132,17'd31190,17'd39916,17'd55133,17'd55134,17'd55135,17'd48363,17'd45033,17'd50474,17'd50659,17'd42873,17'd50474,17'd41409,17'd49379,17'd50366,17'd40218,17'd31352,17'd33952,17'd35426,17'd31352,17'd29977,17'd30279,17'd25553,17'd25430,17'd27145,17'd25944,17'd26523,17'd27761,17'd28854,17'd28133,17'd28370,17'd29104,17'd29247,17'd28371,17'd28487,17'd28487,17'd29247,17'd28854,17'd44826,17'd37513,17'd29379,17'd29379,17'd28727,17'd26902,17'd27514,17'd26064,17'd28599,17'd28597,17'd27882,17'd25567,17'd28598,17'd30606,17'd26062,17'd26174,17'd25833,17'd25949,17'd40965,17'd27513,17'd27765,17'd44105,17'd55136,17'd53782,17'd55137,17'd46321,17'd43281,17'd49381,17'd49787,17'd49891,17'd49984,17'd49390,17'd55138,17'd55139,17'd55140,17'd53194,17'd52426,17'd55141,17'd52817,17'd53558,17'd34459,17'd23732,17'd29827,17'd29975,17'd42744,17'd29828,17'd29686,17'd23565,17'd28851,17'd24898,17'd24744,17'd24252,17'd24742,17'd25030,17'd25709,17'd33000,17'd25438,17'd24898,17'd32659,17'd23384,17'd44107,17'd55142,17'd31658,17'd52172,17'd55143,17'd55144,17'd55145,17'd55146,17'd21534,17'd51655,17'd46775,17'd53786,17'd47749,17'd55147,17'd55148,17'd55149,17'd55150,17'd55151,17'd55152,17'd55153,17'd20817,17'd28053,17'd55154,17'd43725,17'd55155,17'd55059,17'd55156,17'd22933,17'd23453,17'd23107,17'd23457,17'd8911,17'd24476,17'd5607,17'd4840,17'd5328,17'd5002,17'd5005,17'd5004,17'd5335,17'd27935,17'd28185,17'd31717,17'd6554,17'd7499,17'd7499,17'd27696,17'd27696,17'd31888,17'd31888,17'd31888,17'd29593,17'd29593,17'd35052,17'd31888,17'd31888,17'd32074,17'd7499,17'd6391,17'd5614,17'd5005,17'd4841,17'd41459,17'd54861,17'd33841,17'd5001,17'd49597,17'd54765,17'd4369,17'd4370,17'd49896,17'd50488,17'd51931,17'd54499,17'd39474,17'd55157,17'd55158,17'd55159,17'd55160,17'd55066,17'd55067,17'd55161,17'd55162,17'd55070,17'd54870,17'd54772,17'd55163,17'd55164,17'd55073,17'd55074,17'd54973,17'd40713,17'd55165,17'd50385,17'd51411,17'd55166,17'd55078,17'd55167,17'd3222,17'd1121,17'd448,17'd1121,17'd447,17'd2587,17'd1402,17'd3072,17'd1944,17'd960,17'd632,17'd450,17'd238,17'd630,17'd959,17'd795,17'd446,17'd625,17'd11590,17'd1824,17'd38071,17'd3711,17'd7341,17'd55080,17'd55168,17'd55169,17'd55170,17'd53365,17'd55171,17'd55084,17'd24494,17'd2086,17'd54786,17'd53366
},
'{
17'd54978,17'd54978,17'd10802,17'd10669,17'd10547,17'd52621,17'd2597,17'd2596,17'd2257,17'd1416,17'd17,17'd17,17'd18,17'd3905,17'd3905,17'd1128,17'd285,17'd1832,17'd285,17'd285,17'd286,17'd286,17'd7060,17'd27444,17'd4430,17'd4431,17'd3755,17'd3254,17'd2944,17'd2263,17'd2600,17'd55085,17'd21949,17'd22967,17'd481,17'd482,17'd60,17'd303,17'd480,17'd16637,17'd2438,17'd1709,17'd39038,17'd2620,17'd27956,17'd3766,17'd55172,17'd49410,17'd55173,17'd55174,17'd32891,17'd55175,17'd24012,17'd55176,17'd10692,17'd11361,17'd10814,17'd10813,17'd11626,17'd13094,17'd12362,17'd12815,17'd55177,17'd55178,17'd11476,17'd11476,17'd11625,17'd11625,17'd10941,17'd11360,17'd18412,17'd19891,17'd19008,17'd23156,17'd19512,17'd10815,17'd12532,17'd32261,17'd25512,17'd27601,17'd55179,17'd19128,17'd16986,17'd16880,17'd14219,17'd15008,17'd37827,17'd54527,17'd34521,17'd54613,17'd55180,17'd55181,17'd55090,17'd55182,17'd55183,17'd55184,17'd55185,17'd55185,17'd55186,17'd55187,17'd55188,17'd55189,17'd55190,17'd3968,17'd55191,17'd55192,17'd55193,17'd55194,17'd5564,17'd55195,17'd55196,17'd54265,17'd54267,17'd55197,17'd55198,17'd55199,17'd54909,17'd55200,17'd54718,17'd55201,17'd55202,17'd55203,17'd55204,17'd55205,17'd50939,17'd50852,17'd51425,17'd27332,17'd51029,17'd52715,17'd19147,17'd19770,17'd54452,17'd15796,17'd55206,17'd55207,17'd54037,17'd16059,17'd53829,17'd53240,17'd55119,17'd24698,17'd14506,17'd21496,17'd13495,17'd54642,17'd16901,17'd12088,17'd13996,17'd14373,17'd12706,17'd13358,17'd55208,17'd55209,17'd55210,17'd55211,17'd55212,17'd54561,17'd18331,17'd19031,17'd17969,17'd17969,17'd19031,17'd16686,17'd14525,17'd52797,17'd13515,17'd25279,17'd25528,17'd28104,17'd35372,17'd28686,17'd29330,17'd31768,17'd30222,17'd55213,17'd55214,17'd29645,17'd30972,17'd31588,17'd33721,17'd52305,17'd51603,17'd55215,17'd52401,17'd53473,17'd51694,17'd51694,17'd51603,17'd53250,17'd36936,17'd31591,17'd30221,17'd36347,17'd28103,17'd24537,17'd24992,17'd16325,17'd11522,17'd14673,17'd14262,17'd14262,17'd13362,17'd13135,17'd12420,17'd12414,17'd12253,17'd15184,17'd19645,17'd11520,17'd11131,17'd24996,17'd26152,17'd12116,17'd16549,17'd16549,17'd33083,17'd15187,17'd11809,17'd12116,17'd11276,17'd20756,17'd12863,17'd14518,17'd14518,17'd13886,17'd24029,17'd19533,17'd17236,17'd26037,17'd27482,17'd11402,17'd8419,17'd55124,17'd22301,17'd55216,17'd55217,17'd55218,17'd55219,17'd7301,17'd55220,17'd55221,17'd15308,17'd26042,17'd17734,17'd55222,17'd55223,17'd55224,17'd55225,17'd55226,17'd55227,17'd55228,17'd45763,17'd55229,17'd55230,17'd46955,17'd49289,17'd45033,17'd52972,17'd52972,17'd44928,17'd49682,17'd39122,17'd43545,17'd48710,17'd32826,17'd29245,17'd29379,17'd31352,17'd31352,17'd29977,17'd31503,17'd25311,17'd36000,17'd25430,17'd26279,17'd26780,17'd26276,17'd26522,17'd28370,17'd28134,17'd28258,17'd32831,17'd39910,17'd40051,17'd32831,17'd30279,17'd44826,17'd37513,17'd29246,17'd28727,17'd26901,17'd30586,17'd29535,17'd26174,17'd28598,17'd28597,17'd28597,17'd28597,17'd25567,17'd27638,17'd28720,17'd27766,17'd26174,17'd26174,17'd26064,17'd38671,17'd28598,17'd29970,17'd53486,17'd55231,17'd47924,17'd51915,17'd46199,17'd48536,17'd49989,17'd49691,17'd49583,17'd49582,17'd45261,17'd41105,17'd49678,17'd55232,17'd51075,17'd50462,17'd55141,17'd52817,17'd54394,17'd29534,17'd34137,17'd23387,17'd42744,17'd32352,17'd23923,17'd29827,17'd23731,17'd32007,17'd25030,17'd24744,17'd24417,17'd24745,17'd25178,17'd25709,17'd28597,17'd27511,17'd24898,17'd23916,17'd23385,17'd34124,17'd50991,17'd34457,17'd21839,17'd55233,17'd21394,17'd55234,17'd55235,17'd55236,17'd55237,17'd51394,17'd55238,17'd55239,17'd55240,17'd55241,17'd55242,17'd55243,17'd55244,17'd55245,17'd55246,17'd21741,17'd22726,17'd55247,17'd55248,17'd55249,17'd55059,17'd55250,17'd23972,17'd23972,17'd23453,17'd23457,17'd8289,17'd5912,17'd4992,17'd4840,17'd4847,17'd4842,17'd30637,17'd5160,17'd5336,17'd28185,17'd30638,17'd31717,17'd6390,17'd7499,17'd7499,17'd27696,17'd9933,17'd31888,17'd31888,17'd29593,17'd29593,17'd9933,17'd32074,17'd27696,17'd27696,17'd32073,17'd7499,17'd6221,17'd5335,17'd29024,17'd4684,17'd39612,17'd55251,17'd49295,17'd4835,17'd4369,17'd55252,17'd55253,17'd50176,17'd55254,17'd55255,17'd4371,17'd49897,17'd55256,17'd55257,17'd55258,17'd55259,17'd55260,17'd55261,17'd55262,17'd55263,17'd55068,17'd55264,17'd54970,17'd55265,17'd55266,17'd55267,17'd55268,17'd53061,17'd54973,17'd40713,17'd21322,17'd55269,17'd50677,17'd55270,17'd54776,17'd37167,17'd3071,17'd1121,17'd796,17'd1121,17'd959,17'd1402,17'd3072,17'd3072,17'd1120,17'd236,17'd449,17'd450,17'd243,17'd235,17'd447,17'd1402,17'd625,17'd1119,17'd5357,17'd1824,17'd4059,17'd53151,17'd54777,17'd36600,17'd39176,17'd55169,17'd55271,17'd55272,17'd55273,17'd55084,17'd24494,17'd2086,17'd54786,17'd53366
},
'{
17'd54978,17'd54978,17'd10802,17'd10669,17'd10547,17'd52621,17'd2597,17'd2597,17'd2257,17'd1414,17'd17,17'd17,17'd3905,17'd3905,17'd3905,17'd1128,17'd285,17'd1832,17'd285,17'd285,17'd286,17'd286,17'd7060,17'd27444,17'd4430,17'd4431,17'd3755,17'd3254,17'd2944,17'd2264,17'd2600,17'd55274,17'd55275,17'd821,17'd58,17'd22616,17'd20869,17'd60,17'd482,17'd16637,17'd994,17'd1710,17'd55276,17'd55086,17'd34932,17'd27101,17'd26241,17'd20730,17'd49411,17'd6456,17'd32566,17'd34355,17'd55277,17'd49014,17'd10945,17'd10563,17'd10942,17'd54340,17'd54247,17'd12362,17'd20885,17'd12362,17'd54340,17'd55177,17'd55177,17'd11476,17'd15516,17'd11625,17'd11086,17'd54247,17'd17204,17'd17572,17'd17690,17'd19384,17'd16518,17'd17317,17'd12531,17'd20423,17'd28668,17'd41320,17'd30510,17'd30510,17'd17206,17'd20585,17'd16769,17'd15008,17'd55278,17'd32100,17'd34522,17'd54613,17'd55279,17'd55280,17'd55090,17'd55281,17'd55282,17'd55283,17'd55284,17'd54992,17'd55285,17'd55286,17'd55287,17'd55288,17'd55289,17'd55290,17'd3002,17'd55291,17'd55292,17'd55293,17'd55294,17'd55295,17'd5866,17'd55296,17'd55297,17'd55298,17'd55299,17'd55199,17'd55199,17'd55300,17'd55010,17'd55301,17'd55302,17'd55303,17'd55304,17'd55305,17'd55306,17'd55307,17'd55308,17'd9454,17'd26991,17'd26249,17'd52122,17'd19147,17'd54452,17'd55309,17'd16784,17'd55310,17'd55311,17'd54109,17'd14656,17'd53771,17'd55119,17'd55019,17'd12090,17'd54275,17'd13495,17'd13495,17'd54728,17'd12237,17'd12236,17'd13996,17'd13996,17'd13130,17'd55312,17'd55313,17'd55314,17'd54372,17'd55315,17'd55316,17'd45814,17'd19031,17'd17969,17'd17969,17'd38238,17'd17013,17'd15811,17'd21057,17'd13515,17'd13515,17'd24991,17'd27737,17'd35372,17'd28686,17'd29330,17'd31285,17'd28571,17'd55317,17'd55318,17'd47011,17'd34551,17'd30676,17'd31942,17'd54044,17'd52798,17'd51694,17'd52401,17'd52401,17'd51602,17'd51694,17'd53630,17'd34705,17'd34556,17'd33243,17'd34385,17'd30220,17'd34390,17'd28107,17'd24030,17'd24995,17'd14264,17'd11397,17'd10989,17'd14262,17'd13362,17'd12996,17'd11958,17'd12577,17'd12414,17'd12109,17'd13364,17'd11667,17'd11808,17'd24996,17'd26152,17'd9741,17'd11809,17'd11809,17'd15569,17'd9345,17'd11809,17'd16549,17'd11277,17'd11135,17'd11670,17'd11527,17'd10991,17'd13886,17'd24029,17'd18326,17'd16687,17'd10478,17'd27482,17'd9193,17'd18919,17'd15947,17'd19646,17'd21061,17'd55319,17'd55320,17'd55321,17'd21514,17'd19649,17'd19649,17'd15576,17'd54196,17'd55322,17'd55323,17'd55324,17'd55325,17'd55326,17'd55327,17'd46452,17'd33801,17'd35577,17'd55328,17'd47435,17'd39423,17'd45150,17'd55329,17'd52972,17'd44928,17'd51077,17'd49382,17'd42295,17'd46665,17'd46425,17'd36542,17'd31352,17'd27642,17'd31352,17'd29245,17'd29246,17'd31352,17'd25704,17'd25832,17'd25172,17'd26279,17'd25558,17'd26278,17'd26276,17'd28854,17'd28258,17'd32831,17'd28258,17'd27885,17'd29977,17'd37513,17'd44704,17'd38537,17'd44703,17'd28727,17'd28486,17'd27259,17'd28482,17'd27513,17'd28599,17'd33000,17'd28597,17'd28597,17'd28598,17'd28598,17'd28594,17'd27766,17'd25708,17'd25708,17'd28602,17'd28598,17'd28599,17'd27882,17'd43553,17'd55330,17'd55331,17'd47639,17'd51740,17'd48535,17'd49184,17'd49479,17'd49484,17'd49682,17'd49484,17'd55332,17'd55333,17'd49572,17'd55334,17'd54938,17'd54845,17'd55335,17'd53558,17'd34459,17'd24086,17'd23566,17'd30128,17'd37117,17'd29975,17'd29242,17'd28722,17'd30126,17'd29976,17'd28254,17'd24896,17'd24896,17'd24898,17'd25177,17'd28597,17'd28597,17'd27511,17'd24895,17'd23731,17'd28976,17'd31350,17'd34454,17'd43697,17'd46860,17'd55336,17'd54579,17'd55337,17'd55338,17'd55339,17'd55340,17'd46775,17'd54581,17'd55341,17'd55342,17'd23224,17'd55343,17'd55344,17'd55345,17'd55346,17'd55347,17'd21891,17'd26104,17'd22744,17'd54307,17'd53576,17'd24474,17'd22932,17'd23973,17'd55348,17'd23453,17'd23798,17'd24645,17'd24647,17'd4683,17'd4684,17'd37153,17'd31245,17'd5004,17'd5335,17'd5336,17'd28185,17'd30638,17'd31717,17'd6219,17'd7499,17'd7668,17'd27696,17'd9933,17'd29593,17'd29593,17'd29593,17'd29593,17'd9933,17'd32074,17'd27696,17'd27696,17'd32073,17'd6220,17'd5919,17'd5329,17'd4847,17'd4526,17'd55349,17'd55350,17'd4835,17'd4368,17'd55351,17'd55351,17'd55253,17'd49997,17'd55254,17'd52011,17'd54499,17'd38446,17'd51094,17'd55352,17'd55353,17'd55354,17'd55355,17'd55261,17'd55356,17'd55357,17'd55068,17'd55264,17'd54970,17'd55071,17'd54972,17'd55358,17'd55268,17'd55359,17'd55360,17'd40713,17'd55361,17'd55362,17'd3387,17'd55363,17'd54776,17'd53674,17'd960,17'd1121,17'd796,17'd1121,17'd1264,17'd1402,17'd3072,17'd3072,17'd796,17'd55364,17'd631,17'd450,17'd243,17'd235,17'd447,17'd1825,17'd1119,17'd2586,17'd50843,17'd4399,17'd3390,17'd6406,17'd54780,17'd55365,17'd39176,17'd55366,17'd55367,17'd53942,17'd55273,17'd55368,17'd2230,17'd2086,17'd54786,17'd53227
},
'{
17'd10670,17'd54978,17'd10802,17'd10669,17'd10547,17'd52621,17'd2597,17'd2597,17'd2257,17'd1414,17'd17,17'd17,17'd3905,17'd3905,17'd18,17'd1128,17'd285,17'd1832,17'd285,17'd285,17'd286,17'd286,17'd7060,17'd27444,17'd4430,17'd4430,17'd4091,17'd3254,17'd2941,17'd2430,17'd1973,17'd23658,17'd1695,17'd820,17'd14749,17'd61,17'd21022,17'd60,17'd482,17'd16637,17'd994,17'd995,17'd17554,17'd2950,17'd2620,17'd23661,17'd22274,17'd55369,17'd20283,17'd46701,17'd55370,17'd55371,17'd39042,17'd14768,17'd16289,17'd11915,17'd25124,17'd54340,17'd54247,17'd12680,17'd16765,17'd12362,17'd11477,17'd55372,17'd55177,17'd11626,17'd15516,17'd11625,17'd11086,17'd54340,17'd10563,17'd17572,17'd22980,17'd18060,17'd21649,17'd17317,17'd12531,17'd19006,17'd41320,17'd41771,17'd36756,17'd27834,17'd17572,17'd16767,17'd15899,17'd15008,17'd48642,17'd55373,17'd34357,17'd55374,17'd55375,17'd55184,17'd55376,17'd55377,17'd55378,17'd55379,17'd55380,17'd54803,17'd55381,17'd55382,17'd55383,17'd55384,17'd55385,17'd55385,17'd4134,17'd55386,17'd55387,17'd55388,17'd55389,17'd55390,17'd55391,17'd55392,17'd55393,17'd55394,17'd55395,17'd55107,17'd55396,17'd55397,17'd55398,17'd55399,17'd55400,17'd55401,17'd55402,17'd55403,17'd55404,17'd55405,17'd55406,17'd55407,17'd55408,17'd52121,17'd53456,17'd53533,17'd55409,17'd55118,17'd54187,17'd55410,17'd15163,17'd15284,17'd13123,17'd53830,17'd55119,17'd17835,17'd11939,17'd12090,17'd55411,17'd21496,17'd54727,17'd12239,17'd11936,17'd14125,17'd14373,17'd13996,17'd13247,17'd55412,17'd22292,17'd55413,17'd55414,17'd55415,17'd55416,17'd17969,17'd18331,17'd55417,17'd55417,17'd17844,17'd53102,17'd52299,17'd21207,17'd52797,17'd12415,17'd17846,17'd28345,17'd28686,17'd31587,17'd30972,17'd31587,17'd29645,17'd30674,17'd30674,17'd47107,17'd31439,17'd31128,17'd36213,17'd52798,17'd55418,17'd52302,17'd52302,17'd52401,17'd51602,17'd51694,17'd51603,17'd34705,17'd53250,17'd33096,17'd30678,17'd36347,17'd28103,17'd24537,17'd30229,17'd14259,17'd11396,17'd10989,17'd14262,17'd13362,17'd13362,17'd12113,17'd12110,17'd12414,17'd12109,17'd13364,17'd13253,17'd11274,17'd10474,17'd10328,17'd10856,17'd17011,17'd15187,17'd24361,17'd15944,17'd14674,17'd11809,17'd12116,17'd14928,17'd11671,17'd11528,17'd10606,17'd10477,17'd11275,17'd18326,17'd14134,17'd15943,17'd15688,17'd17964,17'd12867,17'd55419,17'd20456,17'd55420,17'd12869,17'd55421,17'd23875,17'd55422,17'd55423,17'd15815,17'd55424,17'd55425,17'd55424,17'd55426,17'd55427,17'd55428,17'd55429,17'd55430,17'd33794,17'd31033,17'd55431,17'd55432,17'd55433,17'd43687,17'd55434,17'd54746,17'd52972,17'd55329,17'd41721,17'd40669,17'd46844,17'd48145,17'd42598,17'd36542,17'd31352,17'd27642,17'd29379,17'd29246,17'd29245,17'd30586,17'd25705,17'd25434,17'd27640,17'd30586,17'd32016,17'd31354,17'd27885,17'd32832,17'd32506,17'd31354,17'd27642,17'd28727,17'd34767,17'd46431,17'd34767,17'd28726,17'd34767,17'd26781,17'd26902,17'd26903,17'd26064,17'd31055,17'd31366,17'd28597,17'd28597,17'd28598,17'd30734,17'd27513,17'd26064,17'd25708,17'd25708,17'd28602,17'd27765,17'd33484,17'd27882,17'd27511,17'd55435,17'd55436,17'd55437,17'd55438,17'd45478,17'd43147,17'd49478,17'd49682,17'd49484,17'd49093,17'd43541,17'd55439,17'd49678,17'd48443,17'd50266,17'd48988,17'd55335,17'd55141,17'd50155,17'd35159,17'd23918,17'd29530,17'd37386,17'd29828,17'd23386,17'd29378,17'd24416,17'd25179,17'd25178,17'd25029,17'd34283,17'd24897,17'd27637,17'd25438,17'd25567,17'd25567,17'd29103,17'd30126,17'd28722,17'd23918,17'd31350,17'd30728,17'd43983,17'd52964,17'd55440,17'd21542,17'd55441,17'd21528,17'd55340,17'd53568,17'd51817,17'd55442,17'd55443,17'd55444,17'd55445,17'd55446,17'd55447,17'd55448,17'd55449,17'd55450,17'd27925,17'd26104,17'd55451,17'd22739,17'd30484,17'd55250,17'd23796,17'd23973,17'd55348,17'd23453,17'd8607,17'd8143,17'd5607,17'd4683,17'd4684,17'd29024,17'd53578,17'd5004,17'd5336,17'd5336,17'd30638,17'd30638,17'd6554,17'd6220,17'd7499,17'd27696,17'd9933,17'd9933,17'd29593,17'd29593,17'd29593,17'd29593,17'd27696,17'd32074,17'd29740,17'd29740,17'd9091,17'd6220,17'd5763,17'd4848,17'd4527,17'd49804,17'd55452,17'd55453,17'd55454,17'd55453,17'd55455,17'd55456,17'd38569,17'd49997,17'd52011,17'd55457,17'd53580,17'd55458,17'd52355,17'd55459,17'd55460,17'd55461,17'd55462,17'd55463,17'd55464,17'd55465,17'd55466,17'd55467,17'd55468,17'd55469,17'd55470,17'd55358,17'd55471,17'd55359,17'd55472,17'd40713,17'd55361,17'd19489,17'd55473,17'd8948,17'd37167,17'd36902,17'd630,17'd796,17'd796,17'd1121,17'd1264,17'd3072,17'd3072,17'd795,17'd1121,17'd631,17'd450,17'd238,17'd630,17'd448,17'd2587,17'd1824,17'd1119,17'd3423,17'd50843,17'd1825,17'd52698,17'd3071,17'd37167,17'd55365,17'd39176,17'd55366,17'd55474,17'd53942,17'd55475,17'd55084,17'd54785,17'd2086,17'd54786,17'd53227
},
'{
17'd10670,17'd54978,17'd10802,17'd10669,17'd10547,17'd52621,17'd2597,17'd2597,17'd1414,17'd2257,17'd17,17'd16,17'd3905,17'd3905,17'd18,17'd20404,17'd26,17'd55476,17'd26,17'd285,17'd286,17'd286,17'd7060,17'd27444,17'd4430,17'd4431,17'd3755,17'd3255,17'd2941,17'd2430,17'd1973,17'd23658,17'd1695,17'd1554,17'd21329,17'd14750,17'd55477,17'd21022,17'd61,17'd22616,17'd63,17'd995,17'd995,17'd1709,17'd55086,17'd34932,17'd54609,17'd55478,17'd55479,17'd44620,17'd55480,17'd55481,17'd34014,17'd14892,17'd15899,17'd10944,17'd10111,17'd9572,17'd10283,17'd20424,17'd20886,17'd20424,17'd25124,17'd55482,17'd54340,17'd11626,17'd12813,17'd15516,17'd11086,17'd54247,17'd10816,17'd16289,17'd16411,17'd17448,17'd17206,17'd17317,17'd12532,17'd17941,17'd21185,17'd27219,17'd27833,17'd21650,17'd17319,17'd16767,17'd15899,17'd14893,17'd50191,17'd55483,17'd50094,17'd55483,17'd55484,17'd55485,17'd55486,17'd55487,17'd55488,17'd55489,17'd55490,17'd55184,17'd54892,17'd55491,17'd55492,17'd55493,17'd55385,17'd55494,17'd54996,17'd55495,17'd55496,17'd55497,17'd55498,17'd55499,17'd55500,17'd55501,17'd55502,17'd6490,17'd55105,17'd55503,17'd55504,17'd55505,17'd55506,17'd55507,17'd55508,17'd55509,17'd55510,17'd55511,17'd55512,17'd55405,17'd55513,17'd55514,17'd25266,17'd26356,17'd26249,17'd53456,17'd19147,17'd55118,17'd55515,17'd15665,17'd55516,17'd55517,17'd14369,17'd55518,17'd54456,17'd16678,17'd11789,17'd11938,17'd54275,17'd21496,17'd21496,17'd54727,17'd12237,17'd18799,17'd13996,17'd12087,17'd13129,17'd18319,17'd20306,17'd23675,17'd55519,17'd55520,17'd55416,17'd17969,17'd17234,17'd18331,17'd55417,17'd17844,17'd17724,17'd16914,17'd21057,17'd15942,17'd14003,17'd17727,17'd28228,17'd29067,17'd30072,17'd31439,17'd30676,17'd30972,17'd47010,17'd46912,17'd47107,17'd47593,17'd30834,17'd31442,17'd52798,17'd55521,17'd52402,17'd52402,17'd52302,17'd52401,17'd51694,17'd51694,17'd51603,17'd35100,17'd32770,17'd32933,17'd29482,17'd30222,17'd27004,17'd25671,17'd24995,17'd17478,17'd13516,17'd14262,17'd12262,17'd13362,17'd12113,17'd12419,17'd12109,17'd12109,17'd13882,17'd20313,17'd14262,17'd16555,17'd10166,17'd12116,17'd11809,17'd9345,17'd15944,17'd8874,17'd15807,17'd15807,17'd11809,17'd12116,17'd9884,17'd11276,17'd15688,17'd14518,17'd28463,17'd18326,17'd11400,17'd20756,17'd40134,17'd55522,17'd8248,17'd55523,17'd20456,17'd55524,17'd55322,17'd55525,17'd55526,17'd55527,17'd55528,17'd8430,17'd55529,17'd55530,17'd55531,17'd55532,17'd55533,17'd55534,17'd55535,17'd23217,17'd32186,17'd28722,17'd55536,17'd54843,17'd40362,17'd55042,17'd55537,17'd50474,17'd44928,17'd45033,17'd50735,17'd48358,17'd46665,17'd43154,17'd32184,17'd35426,17'd32016,17'd31352,17'd33952,17'd29246,17'd29245,17'd27027,17'd24737,17'd25434,17'd26903,17'd33163,17'd35426,17'd35570,17'd31354,17'd32832,17'd27642,17'd28980,17'd34767,17'd46431,17'd46431,17'd34767,17'd28726,17'd34767,17'd28727,17'd26781,17'd27259,17'd25707,17'd32658,17'd28484,17'd27882,17'd25709,17'd28598,17'd27513,17'd40965,17'd27767,17'd26062,17'd26174,17'd27766,17'd27638,17'd25709,17'd27512,17'd27511,17'd33318,17'd55538,17'd48146,17'd55539,17'd51915,17'd48153,17'd49391,17'd49478,17'd49390,17'd48995,17'd48363,17'd52505,17'd55540,17'd49473,17'd55541,17'd53203,17'd54845,17'd48258,17'd50154,17'd32668,17'd23917,17'd29376,17'd29829,17'd38976,17'd29686,17'd34137,17'd29102,17'd25180,17'd25438,17'd27637,17'd28596,17'd34283,17'd25029,17'd25177,17'd27882,17'd25567,17'd25317,17'd25179,17'd28851,17'd28722,17'd31029,17'd44233,17'd32346,17'd21531,17'd52679,17'd55542,17'd21390,17'd55543,17'd51479,17'd55544,17'd53568,17'd51377,17'd55545,17'd30018,17'd55546,17'd55547,17'd55548,17'd33520,17'd55549,17'd55550,17'd33831,17'd55551,17'd55552,17'd28530,17'd23617,17'd24303,17'd53577,17'd55553,17'd55348,17'd55348,17'd23107,17'd7492,17'd7659,17'd5607,17'd5328,17'd37153,17'd29024,17'd31245,17'd25627,17'd5336,17'd5335,17'd30638,17'd28185,17'd6219,17'd7499,17'd29740,17'd27696,17'd9933,17'd9933,17'd29593,17'd29593,17'd29593,17'd29593,17'd29740,17'd29740,17'd29740,17'd9091,17'd6220,17'd5919,17'd5167,17'd4685,17'd39015,17'd55350,17'd55554,17'd55555,17'd49399,17'd39016,17'd55455,17'd55456,17'd38569,17'd55457,17'd52011,17'd49997,17'd54227,17'd52689,17'd54674,17'd55556,17'd55557,17'd55461,17'd55558,17'd55559,17'd54009,17'd55560,17'd55466,17'd55467,17'd55561,17'd53799,17'd55164,17'd27203,17'd55471,17'd55562,17'd55563,17'd54162,17'd2893,17'd54875,17'd9245,17'd55564,17'd37167,17'd52461,17'd960,17'd796,17'd796,17'd1121,17'd795,17'd3072,17'd1402,17'd1264,17'd960,17'd55364,17'd237,17'd243,17'd235,17'd796,17'd795,17'd1824,17'd2586,17'd3423,17'd4712,17'd53068,17'd38716,17'd6084,17'd54776,17'd55365,17'd39176,17'd55366,17'd55474,17'd53942,17'd55565,17'd55566,17'd55567,17'd54425,17'd54786,17'd53227
},
'{
17'd10670,17'd10670,17'd10802,17'd10669,17'd10547,17'd52621,17'd2597,17'd2597,17'd1414,17'd2257,17'd17,17'd17,17'd1416,17'd1416,17'd3905,17'd26127,17'd26,17'd55476,17'd26,17'd285,17'd286,17'd286,17'd7060,17'd27444,17'd4430,17'd4430,17'd4091,17'd3255,17'd2941,17'd2943,17'd2785,17'd22615,17'd40,17'd817,17'd15365,17'd55568,17'd55569,17'd55570,17'd20869,17'd483,17'd832,17'd1980,17'd2790,17'd17554,17'd998,17'd33544,17'd2958,17'd26241,17'd54981,17'd49411,17'd55571,17'd55572,17'd55573,17'd14893,17'd16034,17'd10944,17'd13841,17'd25124,17'd10283,17'd20424,17'd20886,17'd20424,17'd11229,17'd55574,17'd54340,17'd11626,17'd13093,17'd12812,17'd15516,17'd23154,17'd10816,17'd16164,17'd16411,17'd24192,17'd18656,17'd17317,17'd12532,17'd19382,17'd19259,17'd55575,17'd19010,17'd16519,17'd20585,17'd16767,17'd24348,17'd14892,17'd55483,17'd55576,17'd53301,17'd55577,17'd54700,17'd55578,17'd55579,17'd55580,17'd55581,17'd55582,17'd55583,17'd55380,17'd55184,17'd55584,17'd55585,17'd55586,17'd55290,17'd55494,17'd55587,17'd55588,17'd55496,17'd55589,17'd55590,17'd55591,17'd55592,17'd55593,17'd55594,17'd55595,17'd54103,17'd54546,17'd55596,17'd55505,17'd55597,17'd55598,17'd55599,17'd55509,17'd55600,17'd55601,17'd55305,17'd55602,17'd55603,17'd26613,17'd10134,17'd53964,17'd27333,17'd55604,17'd53533,17'd19770,17'd15796,17'd53618,17'd55310,17'd53382,17'd55605,17'd55606,17'd54190,17'd26254,17'd12099,17'd25272,17'd54728,17'd11647,17'd54920,17'd21496,17'd12237,17'd12088,17'd13996,17'd12087,17'd12706,17'd55607,17'd20307,17'd21976,17'd53244,17'd55608,17'd55609,17'd55610,17'd55611,17'd18199,17'd55417,17'd55612,17'd18685,17'd17013,17'd14930,17'd15942,17'd13517,17'd16913,17'd28350,17'd29201,17'd36491,17'd50021,17'd34704,17'd31588,17'd34202,17'd37606,17'd35931,17'd47593,17'd47403,17'd48747,17'd51272,17'd52867,17'd55613,17'd55613,17'd52402,17'd52401,17'd51694,17'd51694,17'd51513,17'd35100,17'd34387,17'd55614,17'd30372,17'd34390,17'd27121,17'd25670,17'd15055,17'd15185,17'd11964,17'd11964,17'd12262,17'd11963,17'd12113,17'd12420,17'd12109,17'd12577,17'd13364,17'd18679,17'd11520,17'd10854,17'd10326,17'd9739,17'd17011,17'd9345,17'd15944,17'd9189,17'd10174,17'd10173,17'd9480,17'd11809,17'd9885,17'd12116,17'd25675,17'd10991,17'd29790,17'd11398,17'd11526,17'd10479,17'd10022,17'd55615,17'd8248,17'd55616,17'd24871,17'd25683,17'd55617,17'd55618,17'd55619,17'd55620,17'd15697,17'd12594,17'd55425,17'd55621,17'd55622,17'd55623,17'd55624,17'd55625,17'd48714,17'd33511,17'd23731,17'd24249,17'd55626,17'd48047,17'd52971,17'd55627,17'd55329,17'd55628,17'd55329,17'd49390,17'd47239,17'd48522,17'd46201,17'd40825,17'd32185,17'd32016,17'd32016,17'd31352,17'd37513,17'd37513,17'd31035,17'd28853,17'd26062,17'd28481,17'd26903,17'd30586,17'd30735,17'd31353,17'd29379,17'd29246,17'd28726,17'd34767,17'd35023,17'd35023,17'd26781,17'd26901,17'd26901,17'd26901,17'd26781,17'd26782,17'd27515,17'd28723,17'd28369,17'd25177,17'd25438,17'd28369,17'd28598,17'd27513,17'd27767,17'd27639,17'd25949,17'd25833,17'd28602,17'd28597,17'd27512,17'd27637,17'd29103,17'd53557,17'd55629,17'd48706,17'd48993,17'd47735,17'd49280,17'd50467,17'd49484,17'd49389,17'd49289,17'd45261,17'd54749,17'd54940,17'd47530,17'd46434,17'd54840,17'd48258,17'd50068,17'd43157,17'd24745,17'd28722,17'd23566,17'd30128,17'd37386,17'd23387,17'd28849,17'd28718,17'd25438,17'd28717,17'd28254,17'd24896,17'd28974,17'd27637,17'd27511,17'd28369,17'd25567,17'd25317,17'd25180,17'd23916,17'd30879,17'd33794,17'd46966,17'd33649,17'd46678,17'd55630,17'd55631,17'd55632,17'd54755,17'd42439,17'd55633,17'd53569,17'd51726,17'd55634,17'd55635,17'd55636,17'd55637,17'd55638,17'd55639,17'd55640,17'd55641,17'd20509,17'd28053,17'd22573,17'd53730,17'd55642,17'd24141,17'd55643,17'd55644,17'd23276,17'd23973,17'd23108,17'd24645,17'd24647,17'd4683,17'd28536,17'd37153,17'd37029,17'd30637,17'd5160,17'd5335,17'd5160,17'd30638,17'd27935,17'd6219,17'd9091,17'd27696,17'd27696,17'd9933,17'd9933,17'd29593,17'd29593,17'd29593,17'd31888,17'd34658,17'd29740,17'd9091,17'd32073,17'd6220,17'd5919,17'd5009,17'd34791,17'd54673,17'd55645,17'd55646,17'd55555,17'd55647,17'd4199,17'd49599,17'd53580,17'd50176,17'd52011,17'd52011,17'd54499,17'd4201,17'd49400,17'd52765,17'd47083,17'd55648,17'd55649,17'd55558,17'd55463,17'd55650,17'd55651,17'd55652,17'd55653,17'd54971,17'd53799,17'd55164,17'd27944,17'd55471,17'd55562,17'd37444,17'd55654,17'd52613,17'd55655,17'd55656,17'd18513,17'd37167,17'd36748,17'd630,17'd796,17'd796,17'd1121,17'd795,17'd3745,17'd795,17'd52021,17'd1265,17'd55364,17'd236,17'd630,17'd235,17'd628,17'd1402,17'd625,17'd445,17'd3391,17'd228,17'd52615,17'd55657,17'd3071,17'd55079,17'd36454,17'd35058,17'd55366,17'd55367,17'd55658,17'd2384,17'd55084,17'd55659,17'd54425,17'd54786,17'd53366
},
'{
17'd10670,17'd10670,17'd10802,17'd10669,17'd10547,17'd52621,17'd2597,17'd2597,17'd2257,17'd2425,17'd1416,17'd17,17'd22965,17'd1416,17'd17,17'd4089,17'd26,17'd26,17'd26,17'd27,17'd286,17'd27,17'd7060,17'd27444,17'd4430,17'd4430,17'd4091,17'd3255,17'd2941,17'd2942,17'd2785,17'd22615,17'd40,17'd817,17'd51,17'd55660,17'd55661,17'd55662,17'd14750,17'd14750,17'd2791,17'd2791,17'd2790,17'd995,17'd998,17'd33056,17'd2446,17'd21798,17'd55663,17'd20139,17'd55664,17'd55665,17'd55666,17'd55667,17'd16033,17'd10565,17'd10286,17'd10284,17'd10283,17'd14472,17'd20886,17'd20886,17'd12066,17'd15897,17'd54247,17'd54247,17'd23154,17'd12813,17'd15516,17'd23154,17'd17317,17'd16164,17'd14768,17'd32894,17'd18657,17'd16518,17'd11362,17'd17941,17'd28204,17'd55575,17'd17942,17'd15524,17'd15899,17'd24348,17'd24348,17'd14346,17'd49814,17'd55668,17'd55576,17'd55669,17'd54172,17'd55670,17'd55671,17'd55377,17'd55672,17'd55673,17'd55674,17'd55280,17'd55675,17'd55676,17'd55677,17'd55678,17'd55679,17'd55680,17'd55681,17'd55682,17'd55683,17'd55684,17'd55685,17'd55686,17'd55687,17'd5566,17'd55688,17'd55689,17'd6490,17'd55690,17'd55396,17'd55505,17'd55691,17'd55597,17'd55300,17'd55508,17'd55600,17'd55692,17'd55693,17'd55694,17'd55603,17'd26613,17'd20894,17'd53964,17'd27333,17'd55604,17'd53533,17'd19770,17'd15796,17'd55695,17'd55696,17'd16053,17'd55697,17'd15285,17'd53895,17'd17835,17'd12099,17'd26143,17'd12237,17'd11647,17'd21199,17'd21496,17'd20601,17'd12089,17'd18799,17'd12236,17'd12087,17'd14662,17'd16060,17'd23676,17'd24850,17'd55698,17'd55123,17'd18199,17'd55611,17'd18199,17'd55417,17'd55612,17'd55699,17'd18685,17'd15811,17'd14526,17'd15570,17'd12415,17'd27349,17'd29201,17'd30220,17'd50021,17'd34704,17'd34835,17'd31129,17'd32282,17'd32919,17'd47295,17'd55700,17'd31762,17'd31943,17'd50863,17'd55701,17'd55702,17'd52799,17'd52401,17'd51694,17'd51602,17'd51694,17'd34705,17'd34387,17'd33096,17'd32597,17'd37205,17'd28103,17'd25925,17'd16203,17'd19920,17'd13762,17'd13516,17'd12262,17'd11963,17'd11806,17'd12420,17'd12580,17'd12414,17'd13882,17'd13363,17'd11667,17'd11274,17'd19282,17'd11134,17'd9619,17'd15180,17'd10174,17'd9194,17'd10336,17'd9743,17'd16328,17'd9479,17'd9480,17'd17011,17'd22131,17'd11528,17'd17966,17'd16687,17'd42674,17'd11276,17'd18196,17'd55703,17'd8248,17'd15693,17'd18921,17'd54737,17'd55704,17'd55705,17'd55525,17'd55706,17'd55707,17'd55708,17'd55709,17'd55710,17'd55711,17'd55712,17'd55713,17'd55714,17'd55715,17'd55716,17'd35999,17'd55717,17'd55718,17'd51740,17'd41268,17'd55719,17'd50474,17'd55720,17'd45033,17'd48263,17'd41414,17'd47238,17'd48710,17'd40520,17'd34637,17'd30735,17'd35426,17'd31353,17'd44826,17'd44704,17'd26901,17'd28725,17'd25949,17'd28481,17'd27515,17'd26902,17'd26901,17'd28979,17'd34767,17'd55721,17'd55721,17'd46431,17'd26781,17'd26781,17'd26902,17'd26902,17'd26901,17'd28486,17'd30586,17'd27259,17'd28481,17'd33507,17'd33000,17'd25317,17'd29970,17'd28130,17'd27638,17'd30606,17'd27767,17'd28481,17'd26174,17'd25565,17'd28720,17'd28717,17'd28719,17'd27637,17'd38667,17'd55722,17'd55723,17'd55724,17'd47734,17'd48155,17'd48154,17'd49289,17'd54572,17'd49389,17'd43419,17'd45368,17'd55725,17'd49374,17'd46757,17'd53414,17'd55335,17'd48445,17'd53262,17'd33483,17'd24252,17'd24902,17'd23566,17'd32191,17'd29686,17'd29242,17'd28975,17'd25180,17'd27765,17'd31366,17'd28254,17'd24897,17'd28596,17'd25177,17'd28369,17'd25567,17'd28598,17'd25317,17'd24898,17'd24415,17'd23917,17'd31029,17'd46669,17'd41726,17'd52438,17'd52153,17'd55726,17'd55727,17'd55728,17'd46340,17'd55729,17'd51238,17'd55730,17'd55731,17'd55732,17'd55733,17'd54302,17'd55734,17'd55735,17'd55736,17'd55737,17'd55738,17'd55739,17'd22745,17'd22750,17'd55642,17'd55740,17'd55741,17'd23276,17'd55644,17'd23452,17'd23278,17'd7657,17'd24647,17'd4683,17'd28536,17'd37153,17'd37288,17'd25627,17'd5335,17'd5335,17'd25627,17'd30638,17'd5614,17'd6219,17'd32073,17'd27696,17'd27696,17'd9933,17'd27815,17'd29593,17'd29593,17'd31888,17'd27696,17'd55742,17'd7499,17'd32073,17'd6554,17'd6391,17'd5919,17'd29024,17'd55743,17'd55350,17'd55744,17'd55646,17'd55745,17'd55746,17'd55647,17'd55747,17'd54499,17'd49997,17'd52011,17'd52011,17'd53580,17'd38446,17'd55748,17'd55749,17'd37298,17'd55750,17'd55649,17'd55751,17'd55559,17'd55752,17'd55463,17'd55753,17'd55754,17'd55755,17'd55266,17'd55164,17'd55358,17'd55471,17'd55074,17'd37444,17'd53589,17'd55756,17'd50496,17'd55656,17'd36600,17'd37167,17'd6867,17'd630,17'd796,17'd796,17'd54778,17'd1402,17'd3745,17'd795,17'd52021,17'd1265,17'd55757,17'd630,17'd235,17'd448,17'd628,17'd1402,17'd3898,17'd2586,17'd3247,17'd1824,17'd53222,17'd3569,17'd7341,17'd55080,17'd55758,17'd39029,17'd55759,17'd55760,17'd55761,17'd55762,17'd55763,17'd2231,17'd2086,17'd55764,17'd55765
},
'{
17'd54978,17'd10670,17'd10669,17'd10669,17'd10547,17'd10547,17'd2258,17'd2596,17'd2257,17'd2257,17'd1414,17'd1414,17'd1414,17'd2257,17'd2257,17'd1416,17'd653,17'd980,17'd27,17'd27,17'd286,17'd286,17'd7060,17'd27444,17'd27444,17'd4248,17'd4091,17'd3595,17'd3254,17'd2943,17'd2262,17'd1968,17'd660,17'd1554,17'd301,17'd55660,17'd55766,17'd21023,17'd68,17'd15366,17'd65,17'd55767,17'd483,17'd668,17'd1290,17'd54789,17'd55768,17'd38205,17'd4751,17'd49109,17'd17800,17'd55769,17'd55770,17'd34519,17'd39796,17'd15899,17'd11088,17'd10691,17'd10283,17'd24975,17'd12532,17'd12532,17'd10815,17'd11629,17'd20424,17'd12680,17'd11229,17'd54340,17'd11086,17'd34015,17'd18884,17'd21808,17'd16167,17'd55771,17'd55772,17'd15898,17'd16766,17'd17941,17'd27834,17'd24688,17'd16768,17'd16032,17'd14219,17'd16034,17'd16519,17'd17448,17'd31917,17'd55773,17'd55774,17'd55775,17'd55776,17'd55670,17'd55283,17'd55090,17'd55777,17'd55778,17'd55779,17'd55780,17'd55490,17'd55781,17'd55782,17'd55783,17'd55784,17'd55785,17'd55786,17'd2841,17'd55787,17'd55788,17'd55789,17'd55790,17'd55791,17'd55792,17'd55793,17'd55794,17'd55795,17'd55796,17'd55797,17'd55798,17'd55799,17'd55800,17'd55597,17'd55598,17'd55801,17'd55802,17'd55803,17'd55804,17'd55805,17'd55806,17'd21196,17'd26026,17'd26356,17'd20598,17'd22123,17'd19770,17'd17955,17'd55807,17'd55808,17'd55809,17'd55810,17'd55811,17'd55812,17'd24988,17'd11793,17'd11504,17'd12089,17'd55813,17'd55814,17'd55815,17'd55816,17'd23848,17'd24852,17'd15935,17'd14125,17'd13995,17'd12708,17'd55817,17'd22292,17'd55818,17'd55819,17'd55820,17'd17234,17'd17234,17'd18331,17'd55417,17'd55821,17'd55822,17'd53102,17'd14930,17'd13252,17'd12418,17'd27486,17'd28945,17'd29930,17'd36491,17'd36491,17'd34835,17'd33096,17'd38498,17'd33568,17'd30973,17'd47295,17'd55823,17'd32761,17'd36354,17'd55521,17'd53323,17'd53322,17'd55824,17'd55825,17'd55826,17'd51602,17'd53630,17'd35100,17'd33243,17'd34385,17'd29482,17'd39070,17'd23511,17'd16324,17'd11960,17'd13762,17'd14262,17'd14262,17'd11963,17'd11806,17'd11961,17'd12419,17'd12110,17'd12111,17'd12718,17'd11961,17'd13516,17'd11131,17'd12863,17'd24037,17'd9039,17'd9040,17'd9040,17'd9621,17'd10336,17'd22813,17'd17601,17'd9620,17'd9344,17'd18080,17'd15048,17'd19155,17'd20312,17'd17847,17'd12116,17'd34382,17'd55827,17'd19923,17'd7953,17'd22480,17'd15306,17'd55828,17'd55829,17'd55830,17'd55831,17'd55832,17'd13009,17'd55833,17'd55834,17'd55835,17'd55836,17'd55837,17'd55838,17'd22854,17'd55839,17'd39134,17'd55037,17'd55840,17'd55841,17'd53196,17'd55842,17'd55843,17'd55844,17'd55845,17'd55846,17'd39432,17'd46435,17'd46200,17'd32005,17'd30735,17'd29245,17'd29245,17'd29246,17'd44704,17'd44703,17'd33963,17'd27640,17'd26530,17'd27514,17'd27640,17'd27259,17'd26782,17'd33963,17'd33963,17'd35023,17'd33963,17'd33963,17'd33963,17'd26781,17'd26902,17'd26902,17'd26902,17'd26902,17'd28853,17'd28482,17'd40828,17'd40828,17'd28481,17'd27766,17'd28720,17'd28130,17'd25317,17'd28130,17'd26064,17'd25949,17'd25833,17'd28602,17'd28717,17'd27764,17'd25568,17'd25030,17'd34282,17'd55847,17'd47048,17'd47725,17'd48781,17'd49586,17'd43281,17'd49183,17'd48995,17'd48995,17'd48361,17'd53988,17'd48046,17'd51739,17'd48785,17'd48784,17'd48258,17'd48258,17'd44105,17'd25032,17'd29100,17'd23564,17'd29686,17'd29374,17'd29827,17'd23384,17'd24416,17'd29101,17'd28597,17'd31520,17'd29548,17'd33666,17'd27637,17'd25317,17'd27638,17'd27513,17'd27638,17'd25709,17'd24896,17'd24416,17'd23917,17'd34894,17'd34108,17'd41275,17'd55848,17'd54847,17'd55234,17'd55849,17'd53655,17'd55850,17'd55851,17'd55852,17'd47749,17'd55853,17'd55854,17'd55855,17'd55548,17'd55856,17'd55857,17'd55858,17'd55859,17'd55860,17'd55861,17'd22397,17'd22217,17'd55155,17'd23621,17'd22931,17'd23106,17'd55862,17'd55863,17'd7657,17'd24478,17'd6381,17'd4840,17'd4686,17'd28536,17'd31245,17'd5167,17'd37030,17'd30638,17'd30638,17'd27935,17'd5615,17'd6219,17'd32073,17'd27696,17'd9933,17'd31888,17'd31888,17'd27815,17'd27696,17'd32074,17'd27696,17'd50282,17'd6853,17'd6554,17'd5614,17'd29159,17'd42031,17'd55864,17'd39314,17'd55865,17'd55866,17'd4030,17'd55867,17'd55868,17'd49498,17'd52183,17'd52183,17'd38193,17'd38193,17'd55869,17'd49897,17'd55870,17'd38450,17'd55871,17'd55872,17'd55259,17'd55461,17'd55873,17'd55874,17'd55875,17'd55463,17'd55876,17'd55877,17'd55878,17'd55164,17'd24492,17'd54774,17'd55879,17'd32879,17'd55880,17'd55165,17'd40860,17'd55881,17'd55882,17'd53745,17'd36323,17'd36748,17'd18144,17'd1121,17'd55657,17'd1264,17'd1402,17'd1402,17'd447,17'd1545,17'd31726,17'd31726,17'd961,17'd1681,17'd959,17'd1264,17'd1825,17'd5195,17'd5357,17'd5195,17'd795,17'd796,17'd53151,17'd54777,17'd8948,17'd40098,17'd19863,17'd55883,17'd55884,17'd55885,17'd55886,17'd2551,17'd55887,17'd55888,17'd55889,17'd55890
},
'{
17'd54978,17'd10802,17'd10669,17'd10669,17'd10547,17'd10547,17'd2258,17'd2596,17'd2425,17'd2257,17'd1414,17'd1414,17'd2257,17'd2257,17'd2257,17'd1414,17'd289,17'd652,17'd28,17'd28,17'd286,17'd286,17'd7060,17'd27444,17'd27444,17'd4248,17'd4091,17'd3595,17'd3254,17'd2943,17'd2262,17'd13303,17'd660,17'd1697,17'd301,17'd55660,17'd55891,17'd1429,17'd55892,17'd20129,17'd55660,17'd15747,17'd61,17'd668,17'd1290,17'd2443,17'd55893,17'd55894,17'd55895,17'd54337,17'd31263,17'd28199,17'd55896,17'd55371,17'd33220,17'd24350,17'd15765,17'd10286,17'd10690,17'd24975,17'd12531,17'd11362,17'd19621,17'd17317,17'd12531,17'd43747,17'd10111,17'd25124,17'd10108,17'd34938,17'd12532,17'd21808,17'd16167,17'd55897,17'd55898,17'd13468,17'd11231,17'd16766,17'd27834,17'd24688,17'd14768,17'd16030,17'd14347,17'd16169,17'd17320,17'd17448,17'd31917,17'd55773,17'd55899,17'd55900,17'd54705,17'd55901,17'd55902,17'd55903,17'd55904,17'd55905,17'd55906,17'd55907,17'd55490,17'd55908,17'd55909,17'd55910,17'd55911,17'd55912,17'd55913,17'd55914,17'd55915,17'd55916,17'd55917,17'd5281,17'd55918,17'd55919,17'd55920,17'd55921,17'd55922,17'd55923,17'd55105,17'd55504,17'd55924,17'd55925,17'd55799,17'd55926,17'd55927,17'd55928,17'd55929,17'd55930,17'd55931,17'd55932,17'd26613,17'd55933,17'd23673,17'd53381,17'd22123,17'd53177,17'd17955,17'd55807,17'd55934,17'd55310,17'd55935,17'd55936,17'd55937,17'd23677,17'd26143,17'd55938,17'd15172,17'd12700,17'd55021,17'd55815,17'd25269,17'd14245,17'd24852,17'd12850,17'd18799,17'd14125,17'd13128,17'd55939,17'd55940,17'd55413,17'd55941,17'd55416,17'd45933,17'd45933,17'd45933,17'd55417,17'd55942,17'd55943,17'd18562,17'd13642,17'd13760,17'd12856,17'd16557,17'd28572,17'd29930,17'd30220,17'd36491,17'd34381,17'd53250,17'd36936,17'd31590,17'd31127,17'd32919,17'd29329,17'd34827,17'd55944,17'd55945,17'd55946,17'd53393,17'd55947,17'd55825,17'd55826,17'd52401,17'd51694,17'd34705,17'd33243,17'd34385,17'd29647,17'd55948,17'd28107,17'd25671,17'd11960,17'd13762,17'd14262,17'd14262,17'd11807,17'd11806,17'd11960,17'd12580,17'd12109,17'd12419,17'd12718,17'd11960,17'd16326,17'd11275,17'd12863,17'd24037,17'd9188,17'd17237,17'd8569,17'd8880,17'd10176,17'd22645,17'd39977,17'd10335,17'd12117,17'd17964,17'd15569,17'd11135,17'd11401,17'd11671,17'd9479,17'd24040,17'd23684,17'd8578,17'd35371,17'd55949,17'd14533,17'd55950,17'd55951,17'd55952,17'd18094,17'd55953,17'd16082,17'd55954,17'd55955,17'd55956,17'd55957,17'd55958,17'd55959,17'd45272,17'd54057,17'd55960,17'd55961,17'd55962,17'd49581,17'd55963,17'd55964,17'd55039,17'd55965,17'd55966,17'd53649,17'd50159,17'd50903,17'd40218,17'd37908,17'd30735,17'd29245,17'd28980,17'd38537,17'd44703,17'd34767,17'd26782,17'd27259,17'd27515,17'd27515,17'd27640,17'd27259,17'd26782,17'd26782,17'd33963,17'd35023,17'd33963,17'd33963,17'd33963,17'd26781,17'd26902,17'd26782,17'd26782,17'd28725,17'd26903,17'd26530,17'd28481,17'd26062,17'd25949,17'd26062,17'd26064,17'd28594,17'd28130,17'd25435,17'd28602,17'd27766,17'd25949,17'd28598,17'd28719,17'd25029,17'd25568,17'd25180,17'd55967,17'd55968,17'd47237,17'd40363,17'd47735,17'd49576,17'd43541,17'd49288,17'd49289,17'd43419,17'd45742,17'd51476,17'd52586,17'd55969,17'd46102,17'd42299,17'd42597,17'd43017,17'd42148,17'd24416,17'd28722,17'd34137,17'd29686,17'd23386,17'd29689,17'd24090,17'd25179,17'd39591,17'd33000,17'd28480,17'd55970,17'd33666,17'd25178,17'd25317,17'd27513,17'd27513,17'd27638,17'd28717,17'd24896,17'd24416,17'd29534,17'd31828,17'd55971,17'd51164,17'd55972,17'd54754,17'd55973,17'd55974,17'd21702,17'd55975,17'd55976,17'd47362,17'd55977,17'd55978,17'd55979,17'd55980,17'd54759,17'd55981,17'd55982,17'd55983,17'd55056,17'd55984,17'd55985,17'd22924,17'd22739,17'd55155,17'd23620,17'd23623,17'd55986,17'd55987,17'd6839,17'd7658,17'd5912,17'd5323,17'd4840,17'd4841,17'd28536,17'd4842,17'd5167,17'd37030,17'd30638,17'd28185,17'd27935,17'd5614,17'd6219,17'd9091,17'd9933,17'd9933,17'd29593,17'd31888,17'd27815,17'd9933,17'd29740,17'd9091,17'd52270,17'd37434,17'd28185,17'd5336,17'd55988,17'd27697,17'd54673,17'd54960,17'd55989,17'd55866,17'd55990,17'd55991,17'd38570,17'd49498,17'd52183,17'd38569,17'd38193,17'd38193,17'd50588,17'd53428,17'd55992,17'd55993,17'd55994,17'd55995,17'd55259,17'd55461,17'd55996,17'd55997,17'd55998,17'd55559,17'd55876,17'd55999,17'd56000,17'd56001,17'd56002,17'd54685,17'd55879,17'd32722,17'd53743,17'd21322,17'd40860,17'd18757,17'd36181,17'd38715,17'd36323,17'd6867,17'd1943,17'd38856,17'd54778,17'd52615,17'd1402,17'd1402,17'd959,17'd1545,17'd31726,17'd1681,17'd961,17'd1545,17'd2113,17'd1402,17'd1824,17'd5629,17'd5357,17'd3898,17'd2587,17'd629,17'd38856,17'd6405,17'd55564,17'd56003,17'd36453,17'd55883,17'd55884,17'd56004,17'd56005,17'd56006,17'd56007,17'd55888,17'd55889,17'd56008
},
'{
17'd54978,17'd10802,17'd10669,17'd10669,17'd10547,17'd52621,17'd2258,17'd2596,17'd2425,17'd2257,17'd2257,17'd1414,17'd2257,17'd2257,17'd2257,17'd1416,17'd2938,17'd653,17'd28,17'd28,17'd28,17'd287,17'd7061,17'd7060,17'd27444,17'd27444,17'd4248,17'd3595,17'd3254,17'd2940,17'd3253,17'd2939,17'd660,17'd1697,17'd301,17'd15248,17'd1429,17'd1150,17'd56009,17'd56010,17'd56011,17'd56012,17'd61,17'd668,17'd2614,17'd40259,17'd56013,17'd34803,17'd41164,17'd56014,17'd4910,17'd56015,17'd56016,17'd56017,17'd33699,17'd18413,17'd15765,17'd10564,17'd10111,17'd9572,17'd11914,17'd11362,17'd11629,17'd11629,17'd12531,17'd43599,17'd11914,17'd11229,17'd54340,17'd34938,17'd12680,17'd15765,17'd48474,17'd56018,17'd55771,17'd14475,17'd16164,17'd21964,17'd16986,17'd16289,17'd16033,17'd32739,17'd32739,17'd16987,17'd17448,17'd17692,17'd24194,17'd55773,17'd56019,17'd56020,17'd56021,17'd54992,17'd56022,17'd56023,17'd56024,17'd56025,17'd55182,17'd56026,17'd56027,17'd56028,17'd56029,17'd56030,17'd56031,17'd54899,17'd56032,17'd56033,17'd2313,17'd56034,17'd5425,17'd56035,17'd56036,17'd56037,17'd56038,17'd56039,17'd56040,17'd56041,17'd56042,17'd56043,17'd56044,17'd55925,17'd56045,17'd55397,17'd55398,17'd55927,17'd56046,17'd56047,17'd56048,17'd56049,17'd26614,17'd22984,17'd25665,17'd25917,17'd52122,17'd53177,17'd19770,17'd10579,17'd11105,17'd56050,17'd56051,17'd56052,17'd56053,17'd55813,17'd24852,17'd11939,17'd12089,17'd13627,17'd55813,17'd55021,17'd55021,17'd21496,17'd12090,17'd12850,17'd12242,17'd15423,17'd12399,17'd55939,17'd56054,17'd23845,17'd53774,17'd56055,17'd13511,17'd45933,17'd45933,17'd55417,17'd55942,17'd55821,17'd18685,17'd17014,17'd13512,17'd14809,17'd49221,17'd28348,17'd29926,17'd29785,17'd36491,17'd34704,17'd33243,17'd35100,17'd51118,17'd33574,17'd31588,17'd30527,17'd29329,17'd39211,17'd35644,17'd52133,17'd53393,17'd53322,17'd52302,17'd52401,17'd52401,17'd51602,17'd51603,17'd33243,17'd31591,17'd30372,17'd34390,17'd34213,17'd18564,17'd14130,17'd15185,17'd11964,17'd14262,17'd11395,17'd11962,17'd11961,17'd12419,17'd12110,17'd12111,17'd12718,17'd11960,17'd19158,17'd11808,17'd11527,17'd24037,17'd9188,17'd12118,17'd8725,17'd11966,17'd8878,17'd9045,17'd10174,17'd12117,17'd16318,17'd26626,17'd9345,17'd11276,17'd19155,17'd11276,17'd10743,17'd16318,17'd56056,17'd11138,17'd13768,17'd24868,17'd11676,17'd56057,17'd56058,17'd56059,17'd56060,17'd55831,17'd11408,17'd55954,17'd56061,17'd56062,17'd56063,17'd56064,17'd56065,17'd56066,17'd23734,17'd56067,17'd56068,17'd48621,17'd55332,17'd55963,17'd55964,17'd56069,17'd56070,17'd56071,17'd39736,17'd46756,17'd46103,17'd32184,17'd32016,17'd30735,17'd31035,17'd28979,17'd28726,17'd34767,17'd33963,17'd27259,17'd27515,17'd26903,17'd27515,17'd27515,17'd26903,17'd27259,17'd28725,17'd26782,17'd27371,17'd33963,17'd33963,17'd26902,17'd26902,17'd26902,17'd26782,17'd27259,17'd27259,17'd27515,17'd27514,17'd27514,17'd26174,17'd25949,17'd26064,17'd30606,17'd28594,17'd26064,17'd27766,17'd27766,17'd28602,17'd27638,17'd28480,17'd28596,17'd24898,17'd28254,17'd30432,17'd50069,17'd50994,17'd47732,17'd47734,17'd48709,17'd49586,17'd48622,17'd49288,17'd45150,17'd49090,17'd48359,17'd53561,17'd51475,17'd53911,17'd48037,17'd49975,17'd42742,17'd43549,17'd25179,17'd24252,17'd30275,17'd23566,17'd29826,17'd29689,17'd29102,17'd24745,17'd39443,17'd25317,17'd28717,17'd27764,17'd37387,17'd55970,17'd29244,17'd25317,17'd27638,17'd30606,17'd28598,17'd28480,17'd24897,17'd24416,17'd30424,17'd39440,17'd56072,17'd52983,17'd56073,17'd52152,17'd56074,17'd55338,17'd54947,17'd56075,17'd56076,17'd56077,17'd56078,17'd56079,17'd56080,17'd56081,17'd56082,17'd56083,17'd56084,17'd56085,17'd20668,17'd56086,17'd22227,17'd29588,17'd56087,17'd53731,17'd23620,17'd23624,17'd55862,17'd56088,17'd8911,17'd6543,17'd6381,17'd4992,17'd4840,17'd4995,17'd5328,17'd5002,17'd5166,17'd5163,17'd30638,17'd28185,17'd27935,17'd27935,17'd6219,17'd7668,17'd27815,17'd9933,17'd29593,17'd29593,17'd9933,17'd9933,17'd7499,17'd37028,17'd33369,17'd28185,17'd5335,17'd5336,17'd35193,17'd4846,17'd39612,17'd55452,17'd56089,17'd56090,17'd56091,17'd56091,17'd38570,17'd49498,17'd55456,17'd50176,17'd56092,17'd38445,17'd38321,17'd53141,17'd56093,17'd55459,17'd56094,17'd3192,17'd56095,17'd56096,17'd55873,17'd55998,17'd55875,17'd55559,17'd55876,17'd56097,17'd56098,17'd56001,17'd56002,17'd56099,17'd56100,17'd56101,17'd53743,17'd21322,17'd19729,17'd18757,17'd2738,17'd1665,17'd35059,17'd52462,17'd1943,17'd3711,17'd54778,17'd38071,17'd5775,17'd1944,17'd234,17'd1681,17'd1681,17'd1681,17'd961,17'd793,17'd447,17'd3072,17'd5195,17'd5629,17'd4712,17'd1825,17'd795,17'd1120,17'd3711,17'd6405,17'd56102,17'd56103,17'd56104,17'd56105,17'd56106,17'd56107,17'd56108,17'd2382,17'd56109,17'd55888,17'd55889,17'd56110
},
'{
17'd10670,17'd10802,17'd10669,17'd10669,17'd52621,17'd52621,17'd2258,17'd2596,17'd2425,17'd2257,17'd2257,17'd1414,17'd2257,17'd2257,17'd2257,17'd2257,17'd1692,17'd653,17'd652,17'd652,17'd28,17'd287,17'd7061,17'd7060,17'd27444,17'd4430,17'd4091,17'd3595,17'd3254,17'd2943,17'd2262,17'd2939,17'd660,17'd56111,17'd301,17'd55660,17'd56112,17'd56113,17'd56114,17'd56115,17'd56116,17'd15122,17'd14871,17'd64,17'd2614,17'd56117,17'd56013,17'd56118,17'd3115,17'd21173,17'd56119,17'd17673,17'd56120,17'd56121,17'd55371,17'd32738,17'd19384,17'd56122,17'd56123,17'd8064,17'd10562,17'd11362,17'd11362,17'd11629,17'd12532,17'd14472,17'd10111,17'd11914,17'd54340,17'd10814,17'd11914,17'd10944,17'd14100,17'd52932,17'd56124,17'd33549,17'd18060,17'd23156,17'd16986,17'd16164,17'd15902,17'd32894,17'd15385,17'd14766,17'd16290,17'd17208,17'd16029,17'd56125,17'd56126,17'd56021,17'd54888,17'd55184,17'd56127,17'd56128,17'd56129,17'd56130,17'd56131,17'd56132,17'd55379,17'd55490,17'd56029,17'd56133,17'd56134,17'd56135,17'd55494,17'd56136,17'd55290,17'd56137,17'd56138,17'd56139,17'd56140,17'd56141,17'd56142,17'd56143,17'd56144,17'd56145,17'd55006,17'd54546,17'd55798,17'd56045,17'd56146,17'd56147,17'd56148,17'd56149,17'd56150,17'd56151,17'd56152,17'd55805,17'd56153,17'd9855,17'd23330,17'd23673,17'd20598,17'd19147,17'd19770,17'd10579,17'd16784,17'd56154,17'd56155,17'd56156,17'd55936,17'd11646,17'd56157,17'd12088,17'd12088,17'd13627,17'd17831,17'd16429,17'd15553,17'd56158,17'd54275,17'd11937,17'd12243,17'd13505,17'd13357,17'd55607,17'd20307,17'd21976,17'd14255,17'd56159,17'd56160,17'd54043,17'd18331,17'd55612,17'd55942,17'd55942,17'd56161,17'd54825,17'd13134,17'd14525,17'd56162,17'd37206,17'd29642,17'd30073,17'd36491,17'd31773,17'd33243,17'd51432,17'd52305,17'd56163,17'd56164,17'd30675,17'd47107,17'd47296,17'd48747,17'd51692,17'd53323,17'd53323,17'd52868,17'd53473,17'd53473,17'd51602,17'd51603,17'd35100,17'd31591,17'd30371,17'd37205,17'd28103,17'd25925,17'd14130,17'd13520,17'd11964,17'd14262,17'd13762,17'd13135,17'd11961,17'd12419,17'd12419,17'd12419,17'd12718,17'd13761,17'd15185,17'd11274,17'd11527,17'd24037,17'd8875,17'd8727,17'd8572,17'd15429,17'd24368,17'd8886,17'd29637,17'd56165,17'd16318,17'd16318,17'd13887,17'd11277,17'd51697,17'd11135,17'd9480,17'd9038,17'd53253,17'd9048,17'd56166,17'd56167,17'd11676,17'd56168,17'd56169,17'd56170,17'd56171,17'd56172,17'd56173,17'd56174,17'd56175,17'd56176,17'd56177,17'd56178,17'd24228,17'd46452,17'd33950,17'd56179,17'd56180,17'd51313,17'd56181,17'd56182,17'd39893,17'd55845,17'd56183,17'd40214,17'd49272,17'd47925,17'd46425,17'd32185,17'd30735,17'd31035,17'd28486,17'd26901,17'd26781,17'd26781,17'd27371,17'd27515,17'd26174,17'd25833,17'd27515,17'd27515,17'd27515,17'd27259,17'd27259,17'd26782,17'd26782,17'd33963,17'd26781,17'd26902,17'd27027,17'd26902,17'd26782,17'd27259,17'd27640,17'd26903,17'd27515,17'd27514,17'd25949,17'd26064,17'd28594,17'd28594,17'd28602,17'd28481,17'd26530,17'd25949,17'd30606,17'd25709,17'd28596,17'd34283,17'd24897,17'd25030,17'd53557,17'd53117,17'd47048,17'd48046,17'd48707,17'd48446,17'd47538,17'd49091,17'd49288,17'd52170,17'd52676,17'd48152,17'd47934,17'd48146,17'd56184,17'd48258,17'd44589,17'd43156,17'd29825,17'd24898,17'd24415,17'd23733,17'd23566,17'd28976,17'd28849,17'd38407,17'd27511,17'd29970,17'd25709,17'd25568,17'd28596,17'd44117,17'd29702,17'd27511,17'd25317,17'd27638,17'd30606,17'd28598,17'd33803,17'd24898,17'd24416,17'd29527,17'd53781,17'd35155,17'd56185,17'd56186,17'd51991,17'd56187,17'd22317,17'd55976,17'd56188,17'd56189,17'd56190,17'd56191,17'd56192,17'd56193,17'd56194,17'd56195,17'd34146,17'd56196,17'd56197,17'd20669,17'd56198,17'd21898,17'd53502,17'd55155,17'd30483,17'd23791,17'd23105,17'd55987,17'd54957,17'd6543,17'd7324,17'd24649,17'd4992,17'd4683,17'd5152,17'd28536,17'd5329,17'd5163,17'd5163,17'd30638,17'd27935,17'd27935,17'd6554,17'd9091,17'd9933,17'd27815,17'd9933,17'd29592,17'd29593,17'd9933,17'd28184,17'd7499,17'd33042,17'd33369,17'd30638,17'd5335,17'd27571,17'd56199,17'd4690,17'd56200,17'd56201,17'd56202,17'd56091,17'd56091,17'd56090,17'd38570,17'd49599,17'd55455,17'd49805,17'd38445,17'd56203,17'd38447,17'd56204,17'd56205,17'd55556,17'd46588,17'd56206,17'd55259,17'd55461,17'd56207,17'd56208,17'd55998,17'd55559,17'd55876,17'd56209,17'd56210,17'd56211,17'd56212,17'd54685,17'd56213,17'd33047,17'd56214,17'd3066,17'd51670,17'd18757,17'd2738,17'd56215,17'd36902,17'd18144,17'd3711,17'd3711,17'd52698,17'd38071,17'd1944,17'd1120,17'd793,17'd1681,17'd1681,17'd961,17'd961,17'd1546,17'd795,17'd3745,17'd5629,17'd5629,17'd4400,17'd3426,17'd1402,17'd1120,17'd38856,17'd6237,17'd55365,17'd56103,17'd56104,17'd56105,17'd56106,17'd56216,17'd56217,17'd2382,17'd56109,17'd56218,17'd56219,17'd56220
},
'{
17'd10925,17'd10924,17'd10669,17'd10669,17'd52621,17'd52621,17'd2597,17'd2596,17'd2257,17'd2257,17'd1414,17'd1414,17'd2257,17'd2257,17'd2257,17'd22965,17'd56221,17'd2938,17'd652,17'd652,17'd652,17'd28,17'd7061,17'd7061,17'd27444,17'd27444,17'd4248,17'd3595,17'd3254,17'd2940,17'd3253,17'd2939,17'd37,17'd56111,17'd301,17'd55660,17'd56112,17'd56222,17'd56222,17'd56223,17'd56224,17'd55660,17'd14750,17'd64,17'd43332,17'd16266,17'd23491,17'd56118,17'd22112,17'd4907,17'd5397,17'd31417,17'd56225,17'd56226,17'd35624,17'd33062,17'd19256,17'd10693,17'd56227,17'd23326,17'd56228,17'd11629,17'd18412,17'd12532,17'd18412,17'd10815,17'd10562,17'd11914,17'd11477,17'd10814,17'd25124,17'd10692,17'd13466,17'd48299,17'd48642,17'd56229,17'd15524,17'd19384,17'd16410,17'd16410,17'd24348,17'd32894,17'd32098,17'd56230,17'd56231,17'd17208,17'd15767,17'd56232,17'd56126,17'd56233,17'd56234,17'd56234,17'd56235,17'd56236,17'd56237,17'd56130,17'd56238,17'd56239,17'd56240,17'd56241,17'd55676,17'd56242,17'd56243,17'd56244,17'd56245,17'd56246,17'd56033,17'd56247,17'd56248,17'd56249,17'd56250,17'd56251,17'd56252,17'd56253,17'd56254,17'd56040,17'd56255,17'd56256,17'd55926,17'd56045,17'd56257,17'd56258,17'd56259,17'd56148,17'd56149,17'd56260,17'd56261,17'd55931,17'd56262,17'd56263,17'd56264,17'd25665,17'd53381,17'd53313,17'd53698,17'd55118,17'd55515,17'd55695,17'd55410,17'd11106,17'd56265,17'd14794,17'd13631,17'd12397,17'd12088,17'd13627,17'd15420,17'd14511,17'd56266,17'd14919,17'd21199,17'd13627,17'd56267,17'd24699,17'd13506,17'd15555,17'd20169,17'd22126,17'd56268,17'd56269,17'd56270,17'd56271,17'd18199,17'd39214,17'd56272,17'd56272,17'd56161,17'd38238,17'd16915,17'd15811,17'd56273,17'd16684,17'd29201,17'd30074,17'd29785,17'd50021,17'd31591,17'd34047,17'd52305,17'd56163,17'd56274,17'd37065,17'd29066,17'd47010,17'd31763,17'd31590,17'd54279,17'd53323,17'd52869,17'd53473,17'd53473,17'd51694,17'd51603,17'd35100,17'd31591,17'd37985,17'd29481,17'd27235,17'd18200,17'd16203,17'd13520,17'd13762,17'd10989,17'd11395,17'd11962,17'd11806,17'd12420,17'd12419,17'd12419,17'd12110,17'd13761,17'd15185,17'd14673,17'd14518,17'd9619,17'd8875,17'd8409,17'd17481,17'd17481,17'd17481,17'd8728,17'd12263,17'd56275,17'd9335,17'd9193,17'd19415,17'd9619,17'd17599,17'd34038,17'd9620,17'd9041,17'd37604,17'd9048,17'd8423,17'd54048,17'd14142,17'd56276,17'd16213,17'd56277,17'd56278,17'd56279,17'd25008,17'd56280,17'd56281,17'd56282,17'd56283,17'd25162,17'd56284,17'd23735,17'd56285,17'd56286,17'd55962,17'd48521,17'd49182,17'd55845,17'd56287,17'd56182,17'd43830,17'd51162,17'd47627,17'd48256,17'd32184,17'd33163,17'd32016,17'd27027,17'd26902,17'd26902,17'd26902,17'd26782,17'd27883,17'd25949,17'd27766,17'd26174,17'd26174,17'd27514,17'd27514,17'd27640,17'd28725,17'd26782,17'd26902,17'd26781,17'd26901,17'd27027,17'd27027,17'd27027,17'd26782,17'd27259,17'd27640,17'd26903,17'd27514,17'd26530,17'd26062,17'd28720,17'd28130,17'd28594,17'd26064,17'd26530,17'd26530,17'd27767,17'd25567,17'd25178,17'd24417,17'd23561,17'd24744,17'd32668,17'd50562,17'd49977,17'd46953,17'd52822,17'd46321,17'd47446,17'd48153,17'd48362,17'd48622,17'd54841,17'd56288,17'd53561,17'd52504,17'd53911,17'd56289,17'd49975,17'd44589,17'd44359,17'd25438,17'd24744,17'd24415,17'd23918,17'd28976,17'd29689,17'd28008,17'd28719,17'd25435,17'd27765,17'd28480,17'd29976,17'd34283,17'd25029,17'd25177,17'd25317,17'd28130,17'd27638,17'd28594,17'd28597,17'd56290,17'd28254,17'd29688,17'd33794,17'd51151,17'd53415,17'd56291,17'd56292,17'd52754,17'd56293,17'd53495,17'd56188,17'd56294,17'd56295,17'd53788,17'd56296,17'd54949,17'd56297,17'd56298,17'd56299,17'd56300,17'd56301,17'd56302,17'd20970,17'd21441,17'd56303,17'd56304,17'd56305,17'd30483,17'd23791,17'd23105,17'd56088,17'd24793,17'd8143,17'd5322,17'd24649,17'd5607,17'd4995,17'd5152,17'd28418,17'd5329,17'd5002,17'd5002,17'd5160,17'd27935,17'd27935,17'd6554,17'd9091,17'd9933,17'd9933,17'd31888,17'd29593,17'd29593,17'd27696,17'd8780,17'd6219,17'd56306,17'd56307,17'd5159,17'd5335,17'd29429,17'd56308,17'd54862,17'd56201,17'd56309,17'd56309,17'd51404,17'd38706,17'd38850,17'd51664,17'd4201,17'd4200,17'd54499,17'd50836,17'd38321,17'd53141,17'd56310,17'd56311,17'd56312,17'd3363,17'd56313,17'd56314,17'd56315,17'd56316,17'd56317,17'd56318,17'd56319,17'd56320,17'd56320,17'd53740,17'd56321,17'd56322,17'd54511,17'd2360,17'd56323,17'd56324,17'd20861,17'd56325,17'd56102,17'd38715,17'd51940,17'd784,17'd630,17'd1121,17'd52698,17'd628,17'd628,17'd1120,17'd796,17'd630,17'd236,17'd961,17'd961,17'd1545,17'd959,17'd795,17'd3745,17'd5629,17'd3898,17'd3591,17'd56326,17'd52918,17'd4059,17'd53151,17'd54780,17'd23300,17'd20560,17'd56104,17'd56327,17'd56106,17'd34929,17'd56328,17'd2382,17'd56329,17'd56218,17'd56219,17'd56330
},
'{
17'd10925,17'd10924,17'd10669,17'd10669,17'd52621,17'd52621,17'd2597,17'd2596,17'd2257,17'd2257,17'd1414,17'd1414,17'd2257,17'd2257,17'd2257,17'd2257,17'd56331,17'd2938,17'd652,17'd652,17'd652,17'd28,17'd7061,17'd7061,17'd27444,17'd27444,17'd4430,17'd3595,17'd3254,17'd2940,17'd3253,17'd2939,17'd1553,17'd296,17'd817,17'd50,17'd56332,17'd56222,17'd56333,17'd56114,17'd56334,17'd56116,17'd65,17'd304,17'd14873,17'd15631,17'd2271,17'd56335,17'd15881,17'd3610,17'd39951,17'd5071,17'd56336,17'd56337,17'd56338,17'd55371,17'd56339,17'd10565,17'd12682,17'd8687,17'd9439,17'd10427,17'd11362,17'd12532,17'd18412,17'd11362,17'd10691,17'd10562,17'd25124,17'd10942,17'd25124,17'd10112,17'd13470,17'd56340,17'd48563,17'd56341,17'd17811,17'd17694,17'd16410,17'd10429,17'd20585,17'd16168,17'd34937,17'd56342,17'd56230,17'd24013,17'd47971,17'd56343,17'd56344,17'd54888,17'd56345,17'd56346,17'd56241,17'd56240,17'd56347,17'd56348,17'd56349,17'd56350,17'd56026,17'd56351,17'd55676,17'd56352,17'd56353,17'd56354,17'd56355,17'd56356,17'd56357,17'd3157,17'd56358,17'd3320,17'd56359,17'd56360,17'd56361,17'd56362,17'd56363,17'd56364,17'd54358,17'd54103,17'd56365,17'd55798,17'd56257,17'd56146,17'd56366,17'd56367,17'd55398,17'd56368,17'd56369,17'd56048,17'd56370,17'd56371,17'd56372,17'd25133,17'd23673,17'd19910,17'd53698,17'd55118,17'd15796,17'd54187,17'd12385,17'd56373,17'd56051,17'd11107,17'd11249,17'd13631,17'd12240,17'd13627,17'd56374,17'd56375,17'd13631,17'd22640,17'd12984,17'd11647,17'd16902,17'd24026,17'd12243,17'd13877,17'd20899,17'd21200,17'd22468,17'd56376,17'd56377,17'd53706,17'd56378,17'd39214,17'd55612,17'd55612,17'd56161,17'd38238,17'd17475,17'd17726,17'd56379,17'd50521,17'd36347,17'd30974,17'd30221,17'd36491,17'd36214,17'd34037,17'd51118,17'd56380,17'd56381,17'd32436,17'd30370,17'd30831,17'd40133,17'd31762,17'd52798,17'd55613,17'd52799,17'd53545,17'd53473,17'd51694,17'd51603,17'd35100,17'd33095,17'd31597,17'd36211,17'd29336,17'd25528,17'd16203,17'd19920,17'd13762,17'd13516,17'd11964,17'd11962,17'd11806,17'd12420,17'd12419,17'd12420,17'd12110,17'd13761,17'd13520,17'd16068,17'd13886,17'd15048,17'd9038,17'd8409,17'd17126,17'd21208,17'd8248,17'd8574,17'd12424,17'd48326,17'd9188,17'd9193,17'd9337,17'd10743,17'd14928,17'd16680,17'd16328,17'd9621,17'd8731,17'd56382,17'd8735,17'd13528,17'd15444,17'd24050,17'd56383,17'd56277,17'd11001,17'd11145,17'd56384,17'd56385,17'd56386,17'd56387,17'd56388,17'd56389,17'd56390,17'd40680,17'd56391,17'd56392,17'd48152,17'd55332,17'd54572,17'd56069,17'd38794,17'd55627,17'd46955,17'd47725,17'd49275,17'd44827,17'd36690,17'd28486,17'd32016,17'd28725,17'd28725,17'd28725,17'd28853,17'd27259,17'd28482,17'd26064,17'd28723,17'd25949,17'd26530,17'd26530,17'd27883,17'd27259,17'd26782,17'd26902,17'd26902,17'd26901,17'd26901,17'd27027,17'd27027,17'd27027,17'd26782,17'd27259,17'd27640,17'd27514,17'd26530,17'd28482,17'd28602,17'd28600,17'd28600,17'd28720,17'd28481,17'd27640,17'd26530,17'd30734,17'd33484,17'd24745,17'd24090,17'd28601,17'd28851,17'd54394,17'd51828,17'd50158,17'd46953,17'd49388,17'd49279,17'd48153,17'd48360,17'd48535,17'd48362,17'd56393,17'd54204,17'd49580,17'd56394,17'd56395,17'd56396,17'd42300,17'd43979,17'd43022,17'd28254,17'd28718,17'd24090,17'd23384,17'd29377,17'd23563,17'd28595,17'd25567,17'd27766,17'd31055,17'd33803,17'd24898,17'd28718,17'd27512,17'd27882,17'd28484,17'd28130,17'd28594,17'd27638,17'd33000,17'd33803,17'd28254,17'd34621,17'd56397,17'd21848,17'd56398,17'd56291,17'd56399,17'd56400,17'd56401,17'd51815,17'd56402,17'd56294,17'd22340,17'd46854,17'd56403,17'd56404,17'd56405,17'd56406,17'd56407,17'd56408,17'd56409,17'd55450,17'd56410,17'd56411,17'd56412,17'd22218,17'd30483,17'd23620,17'd23106,17'd23276,17'd54957,17'd24149,17'd5912,17'd24798,17'd4992,17'd4993,17'd5152,17'd5327,17'd4842,17'd5002,17'd5005,17'd5002,17'd5160,17'd28185,17'd31717,17'd32073,17'd29740,17'd29593,17'd29593,17'd29593,17'd29593,17'd9933,17'd7668,17'd6220,17'd28185,17'd56413,17'd28307,17'd50175,17'd5335,17'd41889,17'd56414,17'd56415,17'd56309,17'd39019,17'd39617,17'd51404,17'd54004,17'd38706,17'd51664,17'd38446,17'd54227,17'd50749,17'd50749,17'd52605,17'd56416,17'd38062,17'd56417,17'd47083,17'd56418,17'd56419,17'd56314,17'd56420,17'd56421,17'd56422,17'd56317,17'd56319,17'd56320,17'd56423,17'd56424,17'd56211,17'd56322,17'd54419,17'd56425,17'd56426,17'd56427,17'd56428,17'd18865,17'd56102,17'd38715,17'd36323,17'd238,17'd630,17'd1121,17'd54778,17'd628,17'd796,17'd1121,17'd960,17'd630,17'd630,17'd961,17'd961,17'd1546,17'd447,17'd1402,17'd3745,17'd5195,17'd1825,17'd56429,17'd56429,17'd52918,17'd53293,17'd56430,17'd54780,17'd23300,17'd20560,17'd56431,17'd56432,17'd34929,17'd56328,17'd56433,17'd2551,17'd56434,17'd56435,17'd56436,17'd56330
},
'{
17'd10924,17'd10924,17'd10669,17'd10669,17'd52621,17'd3429,17'd2597,17'd1414,17'd1414,17'd1414,17'd1414,17'd1414,17'd1414,17'd2257,17'd2257,17'd2257,17'd27442,17'd1416,17'd289,17'd289,17'd653,17'd28,17'd286,17'd286,17'd27444,17'd27444,17'd4430,17'd3908,17'd290,17'd982,17'd32,17'd34,17'd2428,17'd1699,17'd302,17'd55660,17'd56437,17'd56438,17'd56439,17'd56222,17'd56440,17'd56334,17'd66,17'd305,17'd56441,17'd307,17'd2617,17'd2128,17'd32091,17'd41164,17'd39793,17'd40565,17'd25254,17'd56442,17'd56443,17'd55481,17'd32415,17'd15766,17'd10694,17'd9006,17'd22634,17'd10691,17'd11362,17'd12532,17'd11629,17'd11087,17'd10816,17'd10562,17'd11229,17'd25124,17'd54341,17'd24014,17'd10113,17'd48474,17'd49814,17'd56444,17'd34177,17'd16165,17'd15766,17'd10428,17'd29623,17'd16034,17'd35351,17'd56445,17'd34177,17'd15767,17'd47972,17'd53163,17'd56446,17'd56447,17'd56345,17'd56448,17'd56449,17'd55092,17'd56450,17'd56451,17'd56452,17'd56453,17'd56454,17'd56455,17'd56455,17'd56456,17'd56457,17'd56458,17'd56459,17'd56460,17'd56461,17'd3973,17'd56462,17'd56463,17'd56464,17'd56465,17'd56466,17'd56467,17'd56468,17'd56469,17'd56470,17'd53307,17'd54632,17'd56471,17'd56257,17'd56472,17'd56473,17'd56147,17'd56474,17'd56475,17'd56476,17'd56477,17'd56370,17'd56478,17'd56479,17'd56480,17'd25665,17'd53381,17'd18670,17'd56481,17'd56482,17'd56483,17'd56484,17'd14116,17'd56485,17'd56486,17'd11374,17'd56487,17'd12397,17'd12394,17'd56488,17'd56489,17'd13494,17'd56490,17'd56491,17'd12984,17'd23677,17'd24699,17'd13638,17'd12401,17'd21355,17'd56492,17'd21356,17'd56493,17'd56494,17'd56495,17'd56378,17'd56496,17'd55612,17'd56497,17'd56161,17'd56161,17'd18685,17'd56161,17'd18449,17'd56498,17'd31294,17'd38500,17'd30974,17'd36491,17'd34704,17'd33568,17'd35644,17'd52305,17'd31942,17'd31588,17'd29924,17'd29923,17'd51601,17'd47295,17'd31590,17'd55418,17'd53187,17'd52133,17'd51602,17'd51694,17'd51513,17'd35100,17'd33243,17'd36214,17'd29646,17'd28572,17'd26758,17'd16324,17'd19920,17'd13762,17'd13516,17'd11964,17'd11962,17'd11806,17'd12420,17'd12419,17'd12420,17'd12419,17'd13761,17'd13135,17'd13762,17'd10605,17'd22131,17'd9039,17'd8409,17'd8099,17'd18566,17'd18919,17'd8574,17'd23861,17'd25531,17'd9038,17'd9193,17'd9347,17'd18332,17'd9619,17'd14383,17'd10334,17'd9621,17'd8571,17'd56382,17'd8735,17'd14678,17'd10182,17'd15309,17'd14144,17'd56171,17'd56499,17'd56500,17'd56501,17'd56502,17'd56503,17'd56504,17'd56505,17'd56506,17'd50564,17'd56507,17'd56508,17'd55038,17'd56509,17'd52505,17'd55434,17'd54390,17'd56510,17'd56511,17'd39901,17'd47050,17'd46100,17'd32184,17'd31353,17'd28727,17'd31035,17'd27259,17'd26903,17'd26903,17'd28724,17'd27514,17'd27767,17'd28594,17'd28723,17'd26174,17'd27514,17'd27514,17'd27640,17'd28725,17'd26902,17'd27027,17'd26901,17'd26901,17'd26901,17'd27027,17'd27027,17'd26902,17'd26782,17'd27259,17'd27640,17'd26530,17'd26062,17'd28481,17'd26064,17'd28130,17'd28130,17'd28602,17'd26174,17'd26903,17'd26062,17'd31366,17'd28596,17'd24743,17'd30879,17'd34467,17'd48987,17'd49171,17'd50901,17'd50821,17'd47234,17'd48781,17'd51994,17'd48534,17'd45368,17'd48535,17'd48360,17'd53988,17'd53910,17'd51645,17'd56512,17'd48784,17'd49975,17'd42885,17'd43286,17'd27511,17'd24896,17'd24743,17'd28975,17'd29243,17'd29378,17'd28601,17'd25178,17'd28600,17'd28598,17'd31856,17'd33803,17'd24896,17'd24744,17'd25177,17'd25567,17'd28130,17'd28130,17'd28594,17'd28598,17'd25709,17'd27512,17'd27637,17'd33482,17'd56513,17'd35427,17'd56514,17'd56515,17'd47161,17'd22317,17'd56516,17'd53496,17'd46456,17'd56517,17'd56518,17'd47152,17'd56519,17'd56520,17'd56521,17'd56522,17'd56523,17'd56524,17'd56525,17'd56526,17'd56527,17'd56528,17'd56529,17'd22218,17'd56530,17'd23790,17'd23106,17'd23276,17'd24793,17'd6543,17'd6381,17'd24649,17'd5757,17'd4840,17'd47174,17'd5328,17'd5002,17'd4842,17'd4842,17'd5329,17'd5160,17'd5160,17'd28185,17'd9091,17'd27696,17'd31888,17'd29593,17'd29593,17'd31888,17'd27696,17'd7668,17'd6390,17'd30637,17'd30796,17'd28307,17'd28307,17'd25627,17'd56531,17'd56532,17'd56533,17'd56534,17'd56535,17'd56536,17'd56536,17'd53507,17'd52689,17'd56537,17'd52605,17'd50672,17'd50672,17'd38572,17'd49499,17'd56310,17'd56538,17'd56539,17'd37298,17'd55460,17'd56419,17'd56314,17'd56540,17'd56316,17'd56317,17'd56318,17'd56319,17'd56320,17'd56541,17'd56542,17'd56211,17'd56543,17'd56544,17'd56545,17'd56546,17'd56547,17'd56548,17'd18865,17'd36600,17'd36455,17'd36323,17'd238,17'd235,17'd796,17'd52698,17'd628,17'd235,17'd236,17'd237,17'd236,17'd630,17'd1545,17'd1545,17'd959,17'd3248,17'd3072,17'd3745,17'd3898,17'd3426,17'd56326,17'd4229,17'd56549,17'd53068,17'd38716,17'd6237,17'd23300,17'd38577,17'd55366,17'd56550,17'd56106,17'd56551,17'd24163,17'd56552,17'd56553,17'd56554,17'd56555,17'd56556
},
'{
17'd10924,17'd10924,17'd10669,17'd10669,17'd52621,17'd2258,17'd2257,17'd1414,17'd1414,17'd1414,17'd1415,17'd1414,17'd1414,17'd2257,17'd2257,17'd2257,17'd27442,17'd1416,17'd289,17'd289,17'd653,17'd652,17'd27,17'd286,17'd27444,17'd27444,17'd4430,17'd3908,17'd290,17'd982,17'd32,17'd34,17'd2261,17'd38,17'd1419,17'd51,17'd56557,17'd56438,17'd56558,17'd56333,17'd56559,17'd56332,17'd56560,17'd56560,17'd21023,17'd1000,17'd56561,17'd56562,17'd56118,17'd3273,17'd4907,17'd5233,17'd4754,17'd56563,17'd37051,17'd56564,17'd32892,17'd19256,17'd9703,17'd56565,17'd9573,17'd22634,17'd11629,17'd11629,17'd22284,17'd11915,17'd11087,17'd22284,17'd12066,17'd56566,17'd9298,17'd9004,17'd15006,17'd14100,17'd56567,17'd56568,17'd56569,17'd15386,17'd13469,17'd10428,17'd30205,17'd20585,17'd35351,17'd56570,17'd54886,17'd48080,17'd56571,17'd56572,17'd54172,17'd56573,17'd56345,17'd55280,17'd56574,17'd55283,17'd56575,17'd56576,17'd56577,17'd56578,17'd56579,17'd56580,17'd54703,17'd56581,17'd56582,17'd56239,17'd56583,17'd56584,17'd56585,17'd56586,17'd56587,17'd56588,17'd56589,17'd56590,17'd56591,17'd56592,17'd56593,17'd56594,17'd56595,17'd56596,17'd56597,17'd54716,17'd56257,17'd56598,17'd56598,17'd56258,17'd55397,17'd56599,17'd56600,17'd56601,17'd56602,17'd56478,17'd56603,17'd56604,17'd25133,17'd20302,17'd56605,17'd56606,17'd56482,17'd15548,17'd13987,17'd56607,17'd11246,17'd56485,17'd14117,17'd14118,17'd14249,17'd12397,17'd14249,17'd56608,17'd56609,17'd56610,17'd56611,17'd14510,17'd55813,17'd15172,17'd12711,17'd12712,17'd12989,17'd56492,17'd21357,17'd24850,17'd56612,17'd56613,17'd56614,17'd56615,17'd38367,17'd38367,17'd56616,17'd56616,17'd18448,17'd31772,17'd17726,17'd56498,17'd37855,17'd30528,17'd31767,17'd36937,17'd31773,17'd36490,17'd35644,17'd52305,17'd31943,17'd31128,17'd30971,17'd30218,17'd56617,17'd31286,17'd33568,17'd56618,17'd53103,17'd53320,17'd52302,17'd51694,17'd51513,17'd51603,17'd35100,17'd56619,17'd30220,17'd36347,17'd27737,17'd12254,17'd11959,17'd19158,17'd13516,17'd11964,17'd11963,17'd12861,17'd12857,17'd12419,17'd12420,17'd12419,17'd11960,17'd13135,17'd13762,17'd10605,17'd14928,17'd10174,17'd12264,17'd8248,17'd8580,17'd12426,17'd24710,17'd26038,17'd17472,17'd8874,17'd16318,17'd12117,17'd9343,17'd9478,17'd32916,17'd17601,17'd9045,17'd24711,17'd56620,17'd56621,17'd24715,17'd13772,17'd15816,17'd56622,17'd56623,17'd56624,17'd56625,17'd56626,17'd56627,17'd56628,17'd56629,17'd56630,17'd56631,17'd40960,17'd55536,17'd56632,17'd48442,17'd44929,17'd43541,17'd56633,17'd38794,17'd56634,17'd40674,17'd40363,17'd46756,17'd56635,17'd36690,17'd29246,17'd29245,17'd26901,17'd26903,17'd25707,17'd26903,17'd26903,17'd28482,17'd40828,17'd27638,17'd25566,17'd26174,17'd27883,17'd27640,17'd27371,17'd26782,17'd27027,17'd26901,17'd26901,17'd26901,17'd26901,17'd27027,17'd26902,17'd26782,17'd27371,17'd27640,17'd27515,17'd26174,17'd28602,17'd26064,17'd27638,17'd28598,17'd27638,17'd25949,17'd28252,17'd26174,17'd28594,17'd27512,17'd28718,17'd30879,17'd23732,17'd34883,17'd53331,17'd56636,17'd56637,17'd51738,17'd50995,17'd51740,17'd51557,17'd49581,17'd45368,17'd47344,17'd48049,17'd49388,17'd56638,17'd56639,17'd54060,17'd42742,17'd46753,17'd47629,17'd43022,17'd25178,17'd28595,17'd28601,17'd28852,17'd23563,17'd28008,17'd24896,17'd41730,17'd42749,17'd46549,17'd56290,17'd28719,17'd34283,17'd25030,17'd25709,17'd27765,17'd28130,17'd28130,17'd28594,17'd25567,17'd25177,17'd25178,17'd25178,17'd33801,17'd56640,17'd56641,17'd56642,17'd53493,17'd53840,17'd51642,17'd56643,17'd56644,17'd56645,17'd56646,17'd47544,17'd55978,17'd29005,17'd56647,17'd56648,17'd56649,17'd56650,17'd56651,17'd56652,17'd56653,17'd56198,17'd56654,17'd53502,17'd22391,17'd23620,17'd22931,17'd23276,17'd56655,17'd24309,17'd6702,17'd24798,17'd5323,17'd32552,17'd4840,17'd47174,17'd4841,17'd5329,17'd28418,17'd4842,17'd5329,17'd5160,17'd30333,17'd31717,17'd7499,17'd9933,17'd31888,17'd39164,17'd31243,17'd31888,17'd7668,17'd6391,17'd28185,17'd28536,17'd31716,17'd5003,17'd30637,17'd5162,17'd56656,17'd49705,17'd38849,17'd52449,17'd56535,17'd56310,17'd55748,17'd53507,17'd52689,17'd56657,17'd52605,17'd38195,17'd38572,17'd56658,17'd56659,17'd56660,17'd52525,17'd37565,17'd37162,17'd3192,17'd56661,17'd53738,17'd56540,17'd56316,17'd56316,17'd56317,17'd56319,17'd56320,17'd56662,17'd56663,17'd56424,17'd56543,17'd56544,17'd56664,17'd2380,17'd40097,17'd56665,17'd36599,17'd36600,17'd56215,17'd35059,17'd243,17'd235,17'd796,17'd52698,17'd628,17'd630,17'd237,17'd797,17'd236,17'd630,17'd1545,17'd1545,17'd447,17'd3072,17'd3745,17'd3745,17'd1824,17'd52615,17'd56326,17'd4712,17'd56549,17'd38718,17'd18143,17'd6405,17'd36599,17'd39029,17'd55759,17'd56550,17'd56666,17'd56667,17'd56668,17'd56552,17'd56669,17'd56670,17'd56555,17'd56556
},
'{
17'd10925,17'd11071,17'd3593,17'd3593,17'd52621,17'd2426,17'd2257,17'd1414,17'd1416,17'd1416,17'd1416,17'd1416,17'd1414,17'd2257,17'd2257,17'd2257,17'd2257,17'd2257,17'd17,17'd16,17'd653,17'd652,17'd286,17'd27,17'd27,17'd980,17'd653,17'd289,17'd30,17'd469,17'd32,17'd294,17'd2261,17'd38,17'd1419,17'd56671,17'd56557,17'd56559,17'd56672,17'd56673,17'd56674,17'd56675,17'd56115,17'd56676,17'd55892,17'd839,17'd308,17'd2126,17'd23141,17'd2276,17'd56677,17'd39793,17'd20282,17'd18524,17'd56678,17'd56443,17'd56679,17'd19009,17'd13972,17'd15006,17'd9158,17'd56680,17'd11362,17'd11362,17'd10817,17'd30356,17'd19754,17'd22284,17'd10427,17'd10285,17'd56681,17'd56682,17'd11232,17'd13843,17'd54527,17'd56683,17'd56568,17'd16029,17'd13721,17'd10428,17'd30205,17'd16289,17'd56231,17'd56684,17'd56685,17'd32100,17'd33857,17'd56686,17'd54021,17'd54346,17'd56687,17'd56449,17'd56688,17'd56689,17'd55781,17'd56690,17'd56691,17'd56692,17'd56693,17'd56694,17'd56695,17'd54703,17'd56026,17'd56696,17'd56697,17'd56698,17'd56699,17'd56700,17'd56701,17'd56702,17'd56703,17'd56704,17'd56705,17'd56706,17'd56707,17'd56708,17'd56364,17'd56709,17'd50096,17'd54909,17'd55798,17'd56472,17'd56710,17'd56711,17'd56712,17'd56713,17'd56714,17'd34687,17'd56715,17'd56716,17'd56717,17'd56153,17'd56264,17'd56718,17'd18792,17'd56719,17'd56720,17'd15282,17'd13987,17'd56484,17'd56721,17'd56722,17'd11495,17'd56723,17'd11645,17'd14511,17'd14249,17'd13873,17'd56724,17'd56725,17'd56726,17'd56727,17'd14659,17'd55813,17'd13638,17'd12572,17'd18800,17'd12407,17'd21201,17'd24696,17'd56728,17'd54373,17'd54374,17'd56729,17'd38503,17'd55417,17'd56616,17'd56616,17'd31772,17'd18448,17'd18685,17'd37857,17'd37986,17'd30530,17'd30974,17'd30221,17'd36491,17'd34381,17'd34037,17'd51118,17'd31943,17'd31128,17'd56730,17'd27857,17'd28347,17'd51601,17'd47404,17'd56380,17'd53103,17'd53187,17'd51602,17'd51694,17'd51602,17'd34556,17'd53250,17'd31591,17'd37335,17'd36347,17'd27858,17'd18564,17'd18198,17'd12996,17'd11964,17'd11964,17'd11963,17'd12861,17'd12857,17'd12111,17'd12111,17'd12111,17'd12113,17'd11806,17'd11807,17'd10604,17'd16070,17'd8874,17'd15429,17'd13139,17'd8419,17'd9888,17'd8576,17'd56731,17'd16795,17'd10173,17'd25525,17'd15180,17'd13887,17'd9345,17'd56732,17'd22814,17'd9348,17'd11404,17'd56382,17'd56733,17'd56734,17'd13772,17'd56735,17'd14941,17'd56736,17'd56737,17'd56738,17'd56739,17'd56740,17'd56741,17'd56742,17'd23706,17'd45381,17'd40680,17'd56743,17'd56744,17'd53844,17'd45742,17'd49288,17'd55434,17'd44585,17'd56745,17'd53269,17'd47234,17'd47925,17'd46425,17'd30735,17'd29246,17'd28726,17'd26782,17'd26530,17'd28252,17'd28252,17'd25949,17'd27767,17'd40828,17'd27638,17'd28602,17'd26903,17'd33815,17'd33815,17'd26782,17'd26902,17'd33963,17'd33963,17'd28486,17'd26781,17'd26901,17'd27027,17'd27027,17'd28725,17'd27640,17'd26530,17'd28482,17'd28602,17'd28720,17'd28130,17'd27765,17'd30734,17'd26062,17'd28724,17'd31351,17'd28720,17'd25177,17'd24416,17'd28722,17'd23732,17'd24086,17'd33482,17'd56746,17'd56747,17'd50900,17'd54059,17'd55137,17'd51915,17'd48261,17'd56748,17'd48534,17'd49279,17'd51740,17'd47536,17'd53782,17'd49274,17'd51746,17'd43548,17'd43838,17'd43978,17'd28850,17'd24897,17'd28718,17'd34884,17'd23563,17'd47533,17'd56749,17'd29244,17'd43836,17'd25438,17'd28719,17'd25029,17'd56750,17'd25030,17'd27637,17'd28597,17'd28599,17'd28723,17'd28594,17'd28597,17'd25317,17'd29244,17'd32007,17'd25031,17'd56751,17'd22864,17'd51632,17'd52825,17'd53131,17'd56752,17'd56753,17'd56754,17'd56755,17'd56756,17'd22514,17'd56757,17'd56758,17'd56759,17'd56760,17'd56761,17'd56762,17'd56763,17'd56764,17'd56765,17'd56766,17'd56767,17'd56768,17'd53502,17'd22928,17'd23620,17'd22931,17'd23276,17'd54958,17'd24149,17'd6544,17'd24798,17'd5608,17'd32552,17'd4995,17'd4841,17'd4687,17'd28418,17'd28536,17'd4842,17'd5330,17'd5004,17'd31553,17'd6219,17'd7499,17'd32074,17'd29592,17'd39164,17'd31888,17'd9933,17'd7499,17'd37289,17'd5009,17'd29431,17'd4687,17'd26452,17'd30180,17'd5161,17'd56769,17'd49498,17'd39019,17'd53581,17'd52836,17'd55748,17'd55870,17'd53057,17'd56204,17'd52998,17'd4202,17'd52908,17'd56770,17'd56771,17'd37811,17'd52766,17'd55556,17'd37298,17'd56772,17'd56313,17'd56773,17'd53738,17'd56540,17'd56774,17'd56317,17'd56775,17'd56423,17'd56320,17'd56776,17'd56777,17'd56211,17'd55267,17'd56778,17'd56779,17'd56780,17'd23299,17'd56003,17'd55882,17'd36455,17'd56781,17'd800,17'd244,17'd793,17'd959,17'd1545,17'd629,17'd236,17'd797,17'd236,17'd961,17'd31726,17'd56782,17'd959,17'd1264,17'd1402,17'd3745,17'd1824,17'd52615,17'd52615,17'd3591,17'd50843,17'd5937,17'd38857,17'd5627,17'd6083,17'd40098,17'd39325,17'd56783,17'd56432,17'd56784,17'd56551,17'd56785,17'd56786,17'd56669,17'd56554,17'd56787,17'd56788
},
'{
17'd10925,17'd11071,17'd3593,17'd3593,17'd52621,17'd2258,17'd2257,17'd1414,17'd1416,17'd1416,17'd1416,17'd1416,17'd1414,17'd2257,17'd2257,17'd2257,17'd2425,17'd2425,17'd1416,17'd17,17'd2938,17'd652,17'd27,17'd27,17'd27,17'd980,17'd652,17'd289,17'd30,17'd469,17'd32,17'd294,17'd2261,17'd38,17'd1554,17'd818,17'd56789,17'd56559,17'd56672,17'd56790,17'd56791,17'd56792,17'd56793,17'd56437,17'd56794,17'd56795,17'd56796,17'd56797,17'd16638,17'd55894,17'd3767,17'd21336,17'd5069,17'd3931,17'd56798,17'd3454,17'd56799,17'd56800,17'd16028,17'd15138,17'd9574,17'd56680,17'd10427,17'd10563,17'd9158,17'd10693,17'd10944,17'd16518,17'd10816,17'd13327,17'd56682,17'd9004,17'd9573,17'd16880,17'd24013,17'd56801,17'd49199,17'd34178,17'd14100,17'd10113,17'd30205,17'd17319,17'd17209,17'd56685,17'd56802,17'd48298,17'd56571,17'd52850,17'd56803,17'd56804,17'd56687,17'd56805,17'd56574,17'd56689,17'd56028,17'd56806,17'd56807,17'd56808,17'd55487,17'd56454,17'd56809,17'd56809,17'd56026,17'd55910,17'd56810,17'd56811,17'd56812,17'd56813,17'd56814,17'd56815,17'd56816,17'd56817,17'd56818,17'd56819,17'd56820,17'd56821,17'd56822,17'd56470,17'd53091,17'd55690,17'd55396,17'd56257,17'd56823,17'd56823,17'd56824,17'd56712,17'd56825,17'd56826,17'd56827,17'd56828,17'd56829,17'd56830,17'd56831,17'd56832,17'd56833,17'd10955,17'd56834,17'd15282,17'd13987,17'd13987,17'd56484,17'd56484,17'd11372,17'd56835,17'd56836,17'd13626,17'd17339,17'd13873,17'd56837,17'd56838,17'd14243,17'd56726,17'd14655,17'd12985,17'd12089,17'd12402,17'd12402,17'd12403,17'd23675,17'd56839,17'd56840,17'd56841,17'd56842,17'd56843,17'd56729,17'd55417,17'd56616,17'd31772,17'd56844,17'd18448,17'd55699,17'd18562,17'd37855,17'd30528,17'd31767,17'd30221,17'd36491,17'd34704,17'd33720,17'd51118,17'd56163,17'd31441,17'd56845,17'd28345,17'd28347,17'd40440,17'd56846,17'd32920,17'd55418,17'd53187,17'd52302,17'd51693,17'd51602,17'd34556,17'd35100,17'd31591,17'd36491,17'd29481,17'd27857,17'd23855,17'd19408,17'd15053,17'd16326,17'd11964,17'd11963,17'd12861,17'd12857,17'd12857,17'd12857,17'd12111,17'd12113,17'd11806,17'd11807,17'd14931,17'd19642,17'd15944,17'd8412,17'd9745,17'd8581,17'd21824,17'd13256,17'd56731,17'd39977,17'd16328,17'd10173,17'd13887,17'd13887,17'd15180,17'd56732,17'd17473,17'd9041,17'd15429,17'd56382,17'd56847,17'd22479,17'd19539,17'd16081,17'd23529,17'd56736,17'd56848,17'd56849,17'd56850,17'd56851,17'd56852,17'd56853,17'd56854,17'd23569,17'd50730,17'd56286,17'd56855,17'd54131,17'd54841,17'd54572,17'd56856,17'd56857,17'd56181,17'd41269,17'd47531,17'd48145,17'd45878,17'd30735,17'd28980,17'd26781,17'd43290,17'd26530,17'd25707,17'd25833,17'd28481,17'd40965,17'd27513,17'd30606,17'd28602,17'd27515,17'd27640,17'd43290,17'd26782,17'd26781,17'd33963,17'd33963,17'd26781,17'd28486,17'd26901,17'd26782,17'd28725,17'd27259,17'd27515,17'd28482,17'd27767,17'd27638,17'd25567,17'd28369,17'd25567,17'd30606,17'd27515,17'd28978,17'd25707,17'd28717,17'd24745,17'd28722,17'd23565,17'd30275,17'd32186,17'd50463,17'd56636,17'd51386,17'd52330,17'd47534,17'd56858,17'd48442,17'd48142,17'd55725,17'd46199,17'd45034,17'd49889,17'd48260,17'd56859,17'd46101,17'd42299,17'd44478,17'd45749,17'd28721,17'd25177,17'd24896,17'd24252,17'd34884,17'd28129,17'd56749,17'd28974,17'd29101,17'd29825,17'd25178,17'd24898,17'd24897,17'd28595,17'd28254,17'd28717,17'd27765,17'd27638,17'd28723,17'd27638,17'd28597,17'd28369,17'd25179,17'd34276,17'd30733,17'd51229,17'd41112,17'd56860,17'd52346,17'd51654,17'd53652,17'd35710,17'd35571,17'd56861,17'd56862,17'd56863,17'd56864,17'd56865,17'd56866,17'd56867,17'd56868,17'd56869,17'd56870,17'd56871,17'd56872,17'd56873,17'd56874,17'd22058,17'd22218,17'd22929,17'd56875,17'd23792,17'd56655,17'd54764,17'd7324,17'd26217,17'd5323,17'd5607,17'd4840,17'd4683,17'd4686,17'd4686,17'd28418,17'd28536,17'd5005,17'd25627,17'd5004,17'd30333,17'd6219,17'd29740,17'd35052,17'd29592,17'd39164,17'd31888,17'd27696,17'd7668,17'd5337,17'd37153,17'd50585,17'd4847,17'd53578,17'd30180,17'd5007,17'd55254,17'd38570,17'd53581,17'd56876,17'd55748,17'd55748,17'd56876,17'd53057,17'd49499,17'd49499,17'd56877,17'd4202,17'd4032,17'd56878,17'd56879,17'd55749,17'd56880,17'd37162,17'd56881,17'd40094,17'd56773,17'd53738,17'd56540,17'd56774,17'd56422,17'd53798,17'd56423,17'd56320,17'd56542,17'd53798,17'd56424,17'd55267,17'd56425,17'd56882,17'd56883,17'd37572,17'd18865,17'd56102,17'd56884,17'd56781,17'd1115,17'd622,17'd1122,17'd447,17'd959,17'd54604,17'd235,17'd236,17'd235,17'd793,17'd56782,17'd1545,17'd1264,17'd3072,17'd1825,17'd1824,17'd1824,17'd1825,17'd3426,17'd3591,17'd4400,17'd4558,17'd38857,17'd6238,17'd5933,17'd36747,17'd56885,17'd56886,17'd56887,17'd56888,17'd2733,17'd2550,17'd56889,17'd56669,17'd56554,17'd56787,17'd56788
},
'{
17'd10925,17'd11071,17'd3593,17'd3429,17'd2426,17'd2258,17'd2257,17'd1415,17'd17,17'd17,17'd1416,17'd1416,17'd1414,17'd1414,17'd2257,17'd2257,17'd2425,17'd2425,17'd2257,17'd17,17'd2938,17'd653,17'd27,17'd980,17'd27,17'd980,17'd652,17'd289,17'd30,17'd469,17'd32,17'd984,17'd13303,17'd37,17'd1697,17'd818,17'd56789,17'd56890,17'd56792,17'd56891,17'd56892,17'd56438,17'd56223,17'd56893,17'd20272,17'd1430,17'd842,17'd1845,17'd1988,17'd32564,17'd14197,17'd53441,17'd21030,17'd56894,17'd56895,17'd56896,17'd56897,17'd56898,17'd24687,17'd16880,17'd10565,17'd13602,17'd22634,17'd10112,17'd11232,17'd10428,17'd10944,17'd21964,17'd10943,17'd10817,17'd23326,17'd8218,17'd21969,17'd10429,17'd16032,17'd54527,17'd49303,17'd50191,17'd47867,17'd12959,17'd10565,17'd17319,17'd15643,17'd34177,17'd56899,17'd48563,17'd52932,17'd52850,17'd56900,17'd56901,17'd56902,17'd56903,17'd56904,17'd56905,17'd56241,17'd56906,17'd56907,17'd56349,17'd56908,17'd56909,17'd56910,17'd56911,17'd56912,17'd56690,17'd56913,17'd56914,17'd56915,17'd56916,17'd56917,17'd56816,17'd56816,17'd56918,17'd56919,17'd56920,17'd56921,17'd56922,17'd56923,17'd56924,17'd56925,17'd54103,17'd55503,17'd56926,17'd56823,17'd56927,17'd56928,17'd56929,17'd56713,17'd56930,17'd56931,17'd56932,17'd56829,17'd56933,17'd56479,17'd56934,17'd17827,17'd17708,17'd56935,17'd56720,17'd15282,17'd56936,17'd56936,17'd56936,17'd12695,17'd56937,17'd56723,17'd11644,17'd56938,17'd56939,17'd56940,17'd56941,17'd56942,17'd56943,17'd56944,17'd56945,17'd17831,17'd12089,17'd12402,17'd22294,17'd23845,17'd54821,17'd54922,17'd54460,17'd54645,17'd54731,17'd56729,17'd55417,17'd56616,17'd31772,17'd56946,17'd56272,17'd56947,17'd55822,17'd56948,17'd38500,17'd31448,17'd30677,17'd29785,17'd36491,17'd56949,17'd34380,17'd54044,17'd33574,17'd33733,17'd31768,17'd28230,17'd40440,17'd40133,17'd31287,17'd52867,17'd53187,17'd52402,17'd56950,17'd51602,17'd34705,17'd35100,17'd33095,17'd56951,17'd30373,17'd28229,17'd18084,17'd21671,17'd13883,17'd19158,17'd16326,17'd16204,17'd13135,17'd12113,17'd12857,17'd20313,17'd20313,17'd12113,17'd12113,17'd11962,17'd14810,17'd51697,17'd15807,17'd11966,17'd22298,17'd21209,17'd21209,17'd23343,17'd33404,17'd26760,17'd10026,17'd9743,17'd10174,17'd26626,17'd15180,17'd56732,17'd56952,17'd9194,17'd15429,17'd56382,17'd16804,17'd14678,17'd15696,17'd56953,17'd18574,17'd56954,17'd56955,17'd56956,17'd56957,17'd56958,17'd56959,17'd56960,17'd23365,17'd34894,17'd55328,17'd56961,17'd48142,17'd56962,17'd56182,17'd56963,17'd56964,17'd54841,17'd56965,17'd49784,17'd50158,17'd44477,17'd33309,17'd31035,17'd28979,17'd27371,17'd33815,17'd26530,17'd26174,17'd28602,17'd27513,17'd30734,17'd27513,17'd30606,17'd25949,17'd27514,17'd27259,17'd26782,17'd27371,17'd35023,17'd26781,17'd26781,17'd33963,17'd30586,17'd27027,17'd28725,17'd27259,17'd27515,17'd26062,17'd40965,17'd38671,17'd28598,17'd33000,17'd25709,17'd25567,17'd25949,17'd28978,17'd28724,17'd28594,17'd24898,17'd23917,17'd23566,17'd29376,17'd23565,17'd56966,17'd56967,17'd56968,17'd56969,17'd48253,17'd48046,17'd48047,17'd53910,17'd56970,17'd55841,17'd48700,17'd48781,17'd47535,17'd56971,17'd56972,17'd48445,17'd44589,17'd43838,17'd49273,17'd25317,17'd25178,17'd24744,17'd24252,17'd34884,17'd28367,17'd28485,17'd25177,17'd42749,17'd27511,17'd25030,17'd24745,17'd24744,17'd24896,17'd27512,17'd28597,17'd28594,17'd28594,17'd26064,17'd28598,17'd28597,17'd27511,17'd25031,17'd33644,17'd56973,17'd22161,17'd56974,17'd52896,17'd52174,17'd51562,17'd56975,17'd35710,17'd56861,17'd35295,17'd56976,17'd56977,17'd47351,17'd56978,17'd56979,17'd56521,17'd56980,17'd56981,17'd56982,17'd56983,17'd56984,17'd56410,17'd56985,17'd43725,17'd22218,17'd23621,17'd23623,17'd23106,17'd54958,17'd24644,17'd7324,17'd24649,17'd5757,17'd4683,17'd4683,17'd4840,17'd4687,17'd4841,17'd28536,17'd28418,17'd5004,17'd5004,17'd25627,17'd27935,17'd6219,17'd9091,17'd29740,17'd29593,17'd29593,17'd31888,17'd29740,17'd6391,17'd5166,17'd28778,17'd5154,17'd4526,17'd37433,17'd4848,17'd50918,17'd49705,17'd38706,17'd56535,17'd52836,17'd50380,17'd55748,17'd52524,17'd52764,17'd49499,17'd4204,17'd49898,17'd37810,17'd56986,17'd52766,17'd53000,17'd56987,17'd36895,17'd56988,17'd3192,17'd40094,17'd43874,17'd56989,17'd56540,17'd56774,17'd56316,17'd53798,17'd56662,17'd56541,17'd56776,17'd56542,17'd56211,17'd54511,17'd56990,17'd56991,17'd56992,17'd19997,17'd36599,17'd2904,17'd56993,17'd36323,17'd784,17'd799,17'd226,17'd2587,17'd959,17'd448,17'd451,17'd235,17'd448,17'd1546,17'd1545,17'd1546,17'd795,17'd2249,17'd446,17'd1824,17'd4400,17'd4229,17'd3591,17'd3591,17'd4400,17'd6085,17'd38857,17'd6084,17'd55564,17'd56994,17'd39325,17'd56995,17'd56886,17'd56996,17'd56997,17'd2550,17'd56007,17'd56998,17'd56554,17'd56787,17'd56999
},
'{
17'd10924,17'd11071,17'd3593,17'd3593,17'd3429,17'd2258,17'd2257,17'd1415,17'd17,17'd17,17'd17,17'd17,17'd1414,17'd1414,17'd2257,17'd2257,17'd2257,17'd2425,17'd2257,17'd1415,17'd468,17'd653,17'd980,17'd980,17'd27,17'd980,17'd652,17'd289,17'd30,17'd469,17'd32,17'd984,17'd13303,17'd37,17'd1697,17'd57000,17'd57001,17'd56890,17'd56674,17'd56891,17'd57002,17'd57002,17'd57003,17'd57004,17'd57005,17'd57006,17'd843,17'd492,17'd1987,17'd57007,17'd27831,17'd45187,17'd4752,17'd4444,17'd18282,17'd3933,17'd57008,17'd57009,17'd57010,17'd18060,17'd20585,17'd13722,17'd6931,17'd11232,17'd9159,17'd10428,17'd11231,17'd21649,17'd15765,17'd13471,17'd9701,17'd8536,17'd13213,17'd9574,17'd22631,17'd15900,17'd56232,17'd50005,17'd31743,17'd14099,17'd15766,17'd17207,17'd15768,17'd24013,17'd56899,17'd57011,17'd57012,17'd56343,17'd57013,17'd55484,17'd57014,17'd56903,17'd56904,17'd57015,17'd56241,17'd55909,17'd57016,17'd56238,17'd57017,17'd57018,17'd57019,17'd55779,17'd57020,17'd56690,17'd57021,17'd57022,17'd57023,17'd1037,17'd57024,17'd57025,17'd57026,17'd1325,17'd57027,17'd57028,17'd57029,17'd57030,17'd57031,17'd57032,17'd57033,17'd56255,17'd54816,17'd57034,17'd56711,17'd57035,17'd57036,17'd57037,17'd57038,17'd56713,17'd56826,17'd57039,17'd57040,17'd57041,17'd57042,17'd57043,17'd57044,17'd57045,17'd18314,17'd11103,17'd57046,17'd57047,17'd56936,17'd57047,17'd12693,17'd11372,17'd57048,17'd11497,17'd57049,17'd57050,17'd57051,17'd57052,17'd57053,17'd57053,17'd57054,17'd56726,17'd13631,17'd17593,17'd13638,17'd12098,17'd23845,17'd55413,17'd54459,17'd57055,17'd57056,17'd57057,17'd55416,17'd55417,17'd55699,17'd31772,17'd57058,17'd56947,17'd56947,17'd55822,17'd56948,17'd38500,17'd31448,17'd30677,17'd30073,17'd36491,17'd57059,17'd34380,17'd57060,17'd36213,17'd33576,17'd31285,17'd35376,17'd40440,17'd31286,17'd31941,17'd51272,17'd53187,17'd52648,17'd56950,17'd51602,17'd53630,17'd34705,17'd33095,17'd57061,17'd57062,17'd28572,17'd26758,17'd23168,17'd11959,17'd16442,17'd16326,17'd16204,17'd12996,17'd12113,17'd12857,17'd11961,17'd20313,17'd12113,17'd12113,17'd11963,17'd14673,17'd27488,17'd51696,17'd36205,17'd26380,17'd16688,17'd34040,17'd8580,17'd26039,17'd57063,17'd34541,17'd22812,17'd10174,17'd15430,17'd13887,17'd33237,17'd14383,17'd10174,17'd8725,17'd32121,17'd53710,17'd24369,17'd18333,17'd23181,17'd57064,17'd56954,17'd52805,17'd57065,17'd57066,17'd57067,17'd57068,17'd57069,17'd22854,17'd51232,17'd56508,17'd54745,17'd48353,17'd41104,17'd55842,17'd55842,17'd55627,17'd49089,17'd47537,17'd46952,17'd50825,17'd44590,17'd32496,17'd28486,17'd26901,17'd27883,17'd28482,17'd26174,17'd25949,17'd30606,17'd28599,17'd28598,17'd27638,17'd26064,17'd25949,17'd27515,17'd27259,17'd27371,17'd27371,17'd35023,17'd33963,17'd26781,17'd26902,17'd26902,17'd27258,17'd27258,17'd26903,17'd28481,17'd30734,17'd31055,17'd31055,17'd28597,17'd33000,17'd28597,17'd28723,17'd25707,17'd25707,17'd26064,17'd33484,17'd24742,17'd23918,17'd23923,17'd23387,17'd23733,17'd57070,17'd50069,17'd57071,17'd57072,17'd47534,17'd53561,17'd56855,17'd54745,17'd57073,17'd51740,17'd50572,17'd55137,17'd55437,17'd57074,17'd57075,17'd49975,17'd42885,17'd33156,17'd32658,17'd27882,17'd25178,17'd24745,17'd24252,17'd34884,17'd38407,17'd28719,17'd25317,17'd29970,17'd27512,17'd24897,17'd28718,17'd24417,17'd27637,17'd25709,17'd27765,17'd28720,17'd28720,17'd27638,17'd28598,17'd28597,17'd25438,17'd29533,17'd57076,17'd57077,17'd45765,17'd51632,17'd47068,17'd52004,17'd42440,17'd43841,17'd33161,17'd51379,17'd21693,17'd57078,17'd57079,17'd30162,17'd57080,17'd57081,17'd57082,17'd57083,17'd57084,17'd57085,17'd57086,17'd57087,17'd57088,17'd55247,17'd53793,17'd22565,17'd23621,17'd23623,17'd23276,17'd23455,17'd25223,17'd6702,17'd24649,17'd4688,17'd4995,17'd4995,17'd32552,17'd4687,17'd5328,17'd31716,17'd4842,17'd5004,17'd33368,17'd30333,17'd6390,17'd9091,17'd7499,17'd9933,17'd29593,17'd29593,17'd29740,17'd7499,17'd6391,17'd37029,17'd57089,17'd5155,17'd5155,17'd37432,17'd5007,17'd50918,17'd54227,17'd38850,17'd57090,17'd57091,17'd57092,17'd55748,17'd52606,17'd49600,17'd49499,17'd4204,17'd57093,17'd37701,17'd57094,17'd57095,17'd56987,17'd47178,17'd37036,17'd57096,17'd3192,17'd40094,17'd56773,17'd57097,17'd56540,17'd57098,17'd56316,17'd53798,17'd57099,17'd56662,17'd56775,17'd56663,17'd56211,17'd54511,17'd57100,17'd57101,17'd2732,17'd57102,17'd36454,17'd36600,17'd54688,17'd1115,17'd2418,17'd1257,17'd226,17'd447,17'd1546,17'd237,17'd243,17'd630,17'd235,17'd1545,17'd1545,17'd2113,17'd1825,17'd446,17'd624,17'd4712,17'd4400,17'd3591,17'd3591,17'd4400,17'd6085,17'd5356,17'd57103,17'd6405,17'd56102,17'd55168,17'd56885,17'd2555,17'd57104,17'd57105,17'd57106,17'd57107,17'd56007,17'd56998,17'd56554,17'd57108,17'd56999
},
'{
17'd10924,17'd11071,17'd3593,17'd3429,17'd2258,17'd2597,17'd1414,17'd1415,17'd17,17'd17,17'd17,17'd17,17'd1415,17'd1414,17'd2257,17'd2257,17'd2596,17'd2258,17'd2257,17'd17,17'd2938,17'd653,17'd980,17'd980,17'd3906,17'd980,17'd652,17'd29,17'd809,17'd1129,17'd10671,17'd984,17'd471,17'd1553,17'd1695,17'd57000,17'd57001,17'd57109,17'd56440,17'd57110,17'd56333,17'd57002,17'd1151,17'd57111,17'd57112,17'd57113,17'd1293,17'd77,17'd17188,17'd57114,17'd57115,17'd2802,17'd3768,17'd57116,17'd57117,17'd56798,17'd57118,17'd57119,17'd32097,17'd19129,17'd17319,17'd13471,17'd6931,17'd9006,17'd10694,17'd10694,17'd11231,17'd16986,17'd19384,17'd15517,17'd9573,17'd8536,17'd8366,17'd9158,17'd13844,17'd47673,17'd57120,17'd50094,17'd33857,17'd48474,17'd16028,17'd16519,17'd17322,17'd15260,17'd57121,17'd57122,17'd56343,17'd57123,17'd57124,17'd57125,17'd57126,17'd57127,17'd57128,17'd54802,17'd55380,17'd55908,17'd57129,17'd56131,17'd57130,17'd57131,17'd57132,17'd57133,17'd56450,17'd56450,17'd55091,17'd57134,17'd57135,17'd57136,17'd57137,17'd57138,17'd57139,17'd57140,17'd57141,17'd57142,17'd57143,17'd57144,17'd57145,17'd56363,17'd57146,17'd57147,17'd57148,17'd55107,17'd57149,17'd57150,17'd57151,17'd57152,17'd57153,17'd57154,17'd57155,17'd57156,17'd57157,17'd57158,17'd57159,17'd57160,17'd57161,17'd57162,17'd57163,17'd16052,17'd57164,17'd12080,17'd57047,17'd57047,17'd57165,17'd56936,17'd57166,17'd57167,17'd57168,17'd57169,17'd57170,17'd57052,17'd57171,17'd57172,17'd11931,17'd57173,17'd57174,17'd57175,17'd12088,17'd12095,17'd53896,17'd54729,17'd56839,17'd56840,17'd56841,17'd57176,17'd55416,17'd55417,17'd55699,17'd31772,17'd57177,17'd56497,17'd57178,17'd57179,17'd56948,17'd57180,17'd32926,17'd30974,17'd30677,17'd36937,17'd57181,17'd33096,17'd57182,17'd51432,17'd31288,17'd30677,17'd28460,17'd28103,17'd28571,17'd31588,17'd52305,17'd54279,17'd57183,17'd57184,17'd51602,17'd51603,17'd35100,17'd33095,17'd31597,17'd36353,17'd28945,17'd27736,17'd25671,17'd11959,17'd18917,17'd18806,17'd16204,17'd13135,17'd11958,17'd12857,17'd11961,17'd13363,17'd12113,17'd12113,17'd11963,17'd14673,17'd57185,17'd22814,17'd8730,17'd21209,17'd8422,17'd7953,17'd7948,17'd57186,17'd57187,17'd29478,17'd29478,17'd10173,17'd15430,17'd16318,17'd57188,17'd24998,17'd15430,17'd8724,17'd32121,17'd15188,17'd24369,17'd18333,17'd16338,17'd17488,17'd56954,17'd57189,17'd57190,17'd57191,17'd57192,17'd57193,17'd57194,17'd57195,17'd57196,17'd57197,17'd57073,17'd56288,17'd57198,17'd56510,17'd56964,17'd56071,17'd48792,17'd47535,17'd46436,17'd50908,17'd40826,17'd34637,17'd30586,17'd26782,17'd26530,17'd26062,17'd26174,17'd27766,17'd28598,17'd33000,17'd25567,17'd27765,17'd26064,17'd26174,17'd26903,17'd27640,17'd27640,17'd27640,17'd43290,17'd27371,17'd26782,17'd27027,17'd27258,17'd28978,17'd25707,17'd26064,17'd28599,17'd31366,17'd28717,17'd25709,17'd27882,17'd33000,17'd28594,17'd38538,17'd38538,17'd28723,17'd28717,17'd24897,17'd28722,17'd23386,17'd29686,17'd23387,17'd55228,17'd57199,17'd57200,17'd52076,17'd57197,17'd48046,17'd49374,17'd57201,17'd57202,17'd53561,17'd45607,17'd55438,17'd47934,17'd55723,17'd57203,17'd57204,17'd46753,17'd43979,17'd43978,17'd28600,17'd25709,17'd25178,17'd24897,17'd23561,17'd29240,17'd34283,17'd25177,17'd29970,17'd28850,17'd33951,17'd24896,17'd27763,17'd34283,17'd27511,17'd27765,17'd27638,17'd28130,17'd28130,17'd25567,17'd28597,17'd28369,17'd27511,17'd30432,17'd57205,17'd57206,17'd57207,17'd57208,17'd51814,17'd48275,17'd35155,17'd22512,17'd35295,17'd35156,17'd23042,17'd57209,17'd52826,17'd57210,17'd57211,17'd57212,17'd57213,17'd57214,17'd57215,17'd57216,17'd57217,17'd57218,17'd57219,17'd22057,17'd29588,17'd57220,17'd23620,17'd23623,17'd23276,17'd24793,17'd24149,17'd6381,17'd24649,17'd4688,17'd4995,17'd4995,17'd4688,17'd4687,17'd5327,17'd5328,17'd5005,17'd5004,17'd33368,17'd30638,17'd6220,17'd9091,17'd7499,17'd27815,17'd9933,17'd9933,17'd29740,17'd7499,17'd5615,17'd37433,17'd29430,17'd4526,17'd5155,17'd4527,17'd50835,17'd51931,17'd38446,17'd57221,17'd57090,17'd57222,17'd50380,17'd57090,17'd57090,17'd57223,17'd52998,17'd50177,17'd57224,17'd57225,17'd57226,17'd57227,17'd57228,17'd57229,17'd3364,17'd57230,17'd39785,17'd42642,17'd42642,17'd57231,17'd57232,17'd57098,17'd56316,17'd56663,17'd57233,17'd56542,17'd56775,17'd56211,17'd57234,17'd56544,17'd53362,17'd57235,17'd57236,17'd57102,17'd57237,17'd57238,17'd54688,17'd238,17'd242,17'd798,17'd629,17'd1546,17'd56782,17'd631,17'd238,17'd961,17'd961,17'd56782,17'd1545,17'd232,17'd446,17'd446,17'd2586,17'd2586,17'd1260,17'd3591,17'd4712,17'd5357,17'd50843,17'd53068,17'd38716,17'd18385,17'd23300,17'd56994,17'd39325,17'd57239,17'd57240,17'd39028,17'd57241,17'd57107,17'd57242,17'd57243,17'd57244,17'd57245,17'd57246
},
'{
17'd10924,17'd11071,17'd10669,17'd3593,17'd3429,17'd2597,17'd1414,17'd1415,17'd17,17'd17,17'd17,17'd17,17'd1415,17'd1414,17'd2257,17'd2257,17'd2596,17'd2258,17'd2425,17'd1415,17'd468,17'd2938,17'd980,17'd980,17'd3906,17'd980,17'd652,17'd29,17'd809,17'd469,17'd1130,17'd984,17'd811,17'd659,17'd39,17'd57247,17'd57248,17'd57249,17'd56440,17'd56792,17'd56333,17'd57002,17'd1152,17'd57006,17'd57250,17'd57251,17'd57252,17'd57253,17'd57254,17'd57255,17'd57256,17'd21480,17'd26242,17'd57257,17'd57258,17'd57259,17'd57260,17'd57261,17'd57262,17'd57010,17'd18060,17'd15898,17'd6143,17'd12219,17'd12534,17'd9159,17'd16410,17'd16289,17'd16028,17'd30957,17'd8537,17'd9573,17'd23326,17'd13327,17'd10429,17'd14624,17'd57263,17'd53447,17'd53684,17'd15767,17'd15768,17'd17694,17'd16769,17'd16032,17'd31918,17'd57264,17'd56125,17'd57265,17'd57266,17'd57267,17'd57268,17'd57269,17'd57270,17'd56580,17'd55380,17'd57271,17'd57272,17'd57273,17'd55904,17'd57274,17'd57275,17'd57276,17'd56450,17'd57277,17'd57278,17'd57279,17'd57280,17'd57281,17'd57282,17'd57283,17'd57284,17'd57285,17'd57286,17'd4146,17'd57287,17'd57288,17'd56361,17'd56142,17'd57289,17'd57290,17'd55394,17'd57291,17'd56926,17'd56927,17'd57151,17'd57292,17'd57293,17'd57294,17'd57154,17'd57295,17'd57296,17'd57297,17'd57298,17'd57299,17'd57160,17'd57300,17'd57301,17'd57302,17'd57303,17'd12383,17'd14115,17'd12834,17'd12972,17'd13115,17'd57304,17'd13116,17'd57305,17'd57306,17'd57307,17'd57307,17'd57171,17'd57308,17'd11931,17'd57309,17'd57310,17'd57311,17'd12397,17'd13638,17'd12244,17'd26365,17'd55413,17'd57312,17'd57313,17'd56613,17'd57314,17'd55612,17'd55699,17'd31772,17'd57177,17'd56497,17'd57178,17'd57179,17'd56948,17'd38500,17'd31448,17'd30974,17'd31767,17'd30221,17'd57181,17'd31591,17'd57182,17'd34044,17'd34380,17'd34835,17'd28571,17'd30222,17'd28345,17'd31129,17'd34380,17'd52303,17'd57183,17'd57315,17'd52401,17'd51694,17'd34705,17'd33095,17'd31597,17'd29647,17'd28945,17'd27858,17'd25671,17'd21671,17'd17722,17'd12582,17'd16204,17'd13135,17'd11958,17'd12420,17'd11961,17'd13363,17'd12113,17'd12113,17'd12996,17'd14673,17'd57185,17'd57316,17'd57317,17'd8253,17'd57318,17'd35090,17'd7951,17'd8887,17'd23860,17'd16682,17'd29478,17'd16552,17'd15430,17'd8874,17'd16680,17'd14928,17'd15180,17'd8567,17'd8577,17'd16919,17'd13378,17'd15696,17'd13530,17'd17488,17'd57319,17'd57320,17'd57321,17'd57322,17'd54834,17'd56388,17'd57323,17'd46096,17'd57324,17'd54941,17'd54388,17'd56393,17'd56070,17'd56510,17'd56964,17'd43970,17'd48781,17'd48151,17'd48697,17'd42599,17'd32496,17'd33163,17'd27027,17'd27259,17'd27639,17'd25949,17'd25949,17'd26064,17'd28599,17'd25709,17'd28369,17'd25317,17'd28720,17'd25949,17'd28724,17'd27640,17'd27883,17'd27640,17'd27371,17'd27371,17'd26782,17'd27258,17'd29535,17'd26174,17'd27513,17'd32669,17'd31520,17'd28717,17'd25438,17'd25438,17'd25709,17'd28597,17'd28602,17'd38538,17'd27766,17'd33000,17'd24897,17'd24415,17'd34137,17'd29830,17'd23923,17'd24421,17'd50464,17'd57325,17'd57326,17'd57327,17'd49571,17'd48046,17'd57328,17'd57329,17'd54745,17'd56858,17'd47537,17'd49690,17'd51645,17'd57330,17'd57331,17'd57332,17'd47927,17'd33156,17'd33643,17'd28369,17'd33484,17'd27512,17'd24897,17'd28595,17'd34283,17'd27637,17'd28850,17'd29825,17'd27512,17'd57333,17'd28596,17'd28485,17'd25029,17'd29101,17'd28130,17'd27638,17'd28130,17'd27765,17'd25567,17'd25567,17'd27882,17'd27511,17'd25179,17'd35430,17'd41726,17'd57334,17'd57335,17'd52160,17'd42439,17'd43697,17'd22510,17'd23044,17'd31660,17'd57336,17'd57337,17'd57338,17'd57339,17'd57340,17'd55053,17'd33028,17'd57341,17'd57342,17'd33194,17'd57343,17'd57344,17'd57345,17'd55451,17'd22751,17'd57346,17'd56875,17'd23105,17'd55644,17'd24644,17'd24479,17'd24649,17'd4992,17'd32552,17'd4995,17'd4683,17'd32552,17'd4841,17'd5327,17'd4841,17'd5005,17'd30637,17'd33042,17'd31717,17'd6220,17'd7499,17'd7668,17'd27815,17'd27696,17'd27696,17'd7499,17'd6220,17'd30638,17'd29023,17'd39470,17'd5001,17'd4526,17'd50586,17'd50835,17'd51010,17'd57347,17'd52523,17'd53057,17'd57348,17'd57348,17'd57349,17'd53057,17'd49600,17'd49499,17'd57093,17'd57350,17'd57351,17'd57352,17'd57353,17'd36895,17'd57354,17'd46472,17'd39478,17'd39785,17'd57355,17'd57355,17'd57231,17'd57356,17'd57357,17'd56316,17'd56663,17'd57233,17'd56775,17'd56775,17'd56211,17'd57234,17'd56544,17'd57358,17'd57359,17'd57360,17'd57361,17'd57237,17'd57362,17'd54688,17'd238,17'd451,17'd8014,17'd629,17'd1546,17'd57363,17'd797,17'd243,17'd961,17'd1681,17'd57363,17'd52103,17'd231,17'd625,17'd1119,17'd2586,17'd1119,17'd228,17'd4712,17'd11869,17'd11869,17'd5937,17'd57364,17'd56430,17'd54776,17'd23300,17'd56994,17'd56885,17'd57365,17'd57366,17'd57367,17'd51333,17'd57107,17'd57368,17'd57369,17'd57370,17'd56999,17'd57371
},
'{
17'd10924,17'd11071,17'd10669,17'd3429,17'd2258,17'd2597,17'd1414,17'd17,17'd17,17'd17,17'd16,17'd17,17'd1415,17'd1414,17'd1414,17'd2257,17'd2596,17'd2426,17'd2425,17'd1414,17'd468,17'd2938,17'd1278,17'd980,17'd3906,17'd3906,17'd980,17'd29,17'd809,17'd1129,17'd2259,17'd984,17'd658,17'd473,17'd39,17'd57247,17'd57248,17'd56789,17'd56334,17'd56438,17'd57372,17'd57372,17'd1152,17'd1292,17'd57373,17'd57374,17'd495,17'd20407,17'd20409,17'd57375,17'd57256,17'd2802,17'd57376,17'd57257,17'd57377,17'd57378,17'd37711,17'd57379,17'd32567,17'd57380,17'd19256,17'd16880,17'd8537,17'd5409,17'd12534,17'd9159,17'd16410,17'd19255,17'd19256,17'd23501,17'd9300,17'd9158,17'd24014,17'd24014,17'd9574,17'd14623,17'd57381,17'd57382,17'd53080,17'd34178,17'd15521,17'd24687,17'd17448,17'd15902,17'd16166,17'd57383,17'd57384,17'd57385,17'd57386,17'd57013,17'd54706,17'd57387,17'd57388,17'd57389,17'd55280,17'd55380,17'd55490,17'd57390,17'd57391,17'd57392,17'd57393,17'd57394,17'd56132,17'd57395,17'd57278,17'd57396,17'd57397,17'd57398,17'd57399,17'd57400,17'd57401,17'd57139,17'd57402,17'd57403,17'd3976,17'd57404,17'd57405,17'd57406,17'd56363,17'd57407,17'd57408,17'd57409,17'd57410,17'd57411,17'd57412,17'd57292,17'd57413,17'd57414,17'd57415,17'd57154,17'd57416,17'd57417,17'd57418,17'd57419,17'd57420,17'd57421,17'd57422,17'd57423,17'd17590,17'd57424,17'd12692,17'd12834,17'd12972,17'd12972,17'd57425,17'd57426,17'd57427,17'd57428,17'd57429,17'd57430,17'd57171,17'd57308,17'd57431,17'd57431,17'd12840,17'd57432,17'd18910,17'd13627,17'd12402,17'd53896,17'd57433,17'd57434,17'd53316,17'd53975,17'd54278,17'd17844,17'd18448,17'd55699,17'd57435,17'd38367,17'd57436,17'd57437,17'd57438,17'd57180,17'd35099,17'd31448,17'd30677,17'd30677,17'd57439,17'd34385,17'd35934,17'd51513,17'd35644,17'd34203,17'd29067,17'd28460,17'd28345,17'd29925,17'd33875,17'd51693,17'd57440,17'd57315,17'd52401,17'd51513,17'd35100,17'd33095,17'd36214,17'd29647,17'd28945,17'd27349,17'd23855,17'd16203,17'd18198,17'd18917,17'd12996,17'd13135,17'd11958,17'd12420,17'd13883,17'd11960,17'd11958,17'd12858,17'd16204,17'd14262,17'd26037,17'd22646,17'd57186,17'd7951,17'd57441,17'd57442,17'd25283,17'd57443,17'd26038,17'd29334,17'd16439,17'd34541,17'd15430,17'd9192,17'd14928,17'd14928,17'd15180,17'd8567,17'd8577,17'd16332,17'd8427,17'd19539,17'd13143,17'd57444,17'd57445,17'd57446,17'd56502,17'd57447,17'd57448,17'd57449,17'd57450,17'd51473,17'd57451,17'd57452,17'd48353,17'd54661,17'd57453,17'd57454,17'd56964,17'd40516,17'd56858,17'd52980,17'd44228,17'd33942,17'd33163,17'd27027,17'd26782,17'd27514,17'd27767,17'd25708,17'd28481,17'd27513,17'd33000,17'd28717,17'd28850,17'd25317,17'd28594,17'd25949,17'd26903,17'd27515,17'd27514,17'd27514,17'd27259,17'd28725,17'd28725,17'd26903,17'd26530,17'd40965,17'd39283,17'd46549,17'd27512,17'd25320,17'd29244,17'd25320,17'd25438,17'd28130,17'd25708,17'd25949,17'd28599,17'd28719,17'd24252,17'd30275,17'd28976,17'd29830,17'd23566,17'd57455,17'd51553,17'd57456,17'd50992,17'd55968,17'd53989,17'd54745,17'd57457,17'd57329,17'd53910,17'd51646,17'd57458,17'd51389,17'd51310,17'd57459,17'd48612,17'd44934,17'd44231,17'd38538,17'd28600,17'd25709,17'd33484,17'd27512,17'd28596,17'd28485,17'd25029,17'd29103,17'd41730,17'd27511,17'd33951,17'd57333,17'd27764,17'd27512,17'd25438,17'd25317,17'd28130,17'd28130,17'd27765,17'd25567,17'd28369,17'd28369,17'd33000,17'd25709,17'd25178,17'd35865,17'd33646,17'd46776,17'd52262,17'd52085,17'd34880,17'd57460,17'd21695,17'd33162,17'd54395,17'd57461,17'd57462,17'd57463,17'd57464,17'd57465,17'd57466,17'd27913,17'd57467,17'd57085,17'd57468,17'd57469,17'd20824,17'd42459,17'd28530,17'd22218,17'd56530,17'd56875,17'd23105,17'd57470,17'd23279,17'd7006,17'd5322,17'd5607,17'd4995,17'd4995,17'd4840,17'd4840,17'd5327,17'd5327,17'd4686,17'd5002,17'd33368,17'd33369,17'd6390,17'd9091,17'd7499,17'd8780,17'd8780,17'd7499,17'd9091,17'd9091,17'd6708,17'd37288,17'd57471,17'd5154,17'd44010,17'd55061,17'd56769,17'd51931,17'd54499,17'd49400,17'd52606,17'd57348,17'd57348,17'd57472,17'd57473,17'd57474,17'd49499,17'd57475,17'd57476,17'd57477,17'd52273,17'd57478,17'd57479,17'd57480,17'd36896,17'd57481,17'd39478,17'd39785,17'd3045,17'd57355,17'd57231,17'd57356,17'd57357,17'd56316,17'd57233,17'd57233,17'd56775,17'd56775,17'd56211,17'd56321,17'd57482,17'd57483,17'd2550,17'd57484,17'd57361,17'd57485,17'd57486,17'd239,17'd242,17'd798,17'd8014,17'd629,17'd1545,17'd57487,17'd237,17'd242,17'd961,17'd1681,17'd31250,17'd7681,17'd623,17'd624,17'd3247,17'd2586,17'd3246,17'd3897,17'd4575,17'd3897,17'd4712,17'd3591,17'd53149,17'd3222,17'd56215,17'd39481,17'd39176,17'd39325,17'd57488,17'd57489,17'd55269,17'd51333,17'd57107,17'd57368,17'd57490,17'd57370,17'd57491,17'd57492
},
'{
17'd10924,17'd11071,17'd10669,17'd3429,17'd2258,17'd2597,17'd1414,17'd17,17'd17,17'd17,17'd16,17'd16,17'd1415,17'd1414,17'd1414,17'd2257,17'd2596,17'd2426,17'd57493,17'd1414,17'd30,17'd1692,17'd2938,17'd1278,17'd1278,17'd980,17'd652,17'd29,17'd809,17'd1129,17'd2259,17'd984,17'd658,17'd473,17'd39,17'd661,17'd819,17'd50,17'd56334,17'd56438,17'd57002,17'd1151,17'd1152,17'd1292,17'd57373,17'd57252,17'd1154,17'd57494,17'd1565,17'd57495,17'd16639,17'd2960,17'd2450,17'd57257,17'd57496,17'd57497,17'd16974,17'd57498,17'd34804,17'd57499,17'd57500,17'd13601,17'd8538,17'd5837,17'd9703,17'd9440,17'd10565,17'd20585,17'd13844,17'd23837,17'd13972,17'd9702,17'd13327,17'd9439,17'd9702,17'd13842,17'd57501,17'd53163,17'd53685,17'd50191,17'd15642,17'd15523,17'd22980,17'd16169,17'd16031,17'd48735,17'd57502,17'd57503,17'd49303,17'd57504,17'd57505,17'd57506,17'd57507,17'd57508,17'd57509,17'd57510,17'd57511,17'd56128,17'd57512,17'd57513,17'd57514,17'd57515,17'd57516,17'd56579,17'd56579,17'd57517,17'd57518,17'd57519,17'd57140,17'd57283,17'd57520,17'd57521,17'd57522,17'd57523,17'd57524,17'd57525,17'd57526,17'd57527,17'd57528,17'd57529,17'd56145,17'd55006,17'd57530,17'd55925,17'd56927,17'd57413,17'd57531,17'd57413,17'd57532,17'd57533,17'd57038,17'd57534,17'd57535,17'd57536,17'd57419,17'd57537,17'd57538,17'd57539,17'd16188,17'd12550,17'd13743,17'd57540,17'd12834,17'd12972,17'd57541,17'd12974,17'd57542,17'd57543,17'd57428,17'd57306,17'd57544,17'd57545,17'd57546,17'd57546,17'd57547,17'd57310,17'd13869,17'd11785,17'd12093,17'd12244,17'd57548,17'd57549,17'd52864,17'd57550,17'd57551,17'd17844,17'd18448,17'd55699,17'd57435,17'd56497,17'd57552,17'd55943,17'd57553,17'd57180,17'd35099,17'd31767,17'd30677,17'd30677,17'd57554,17'd54732,17'd36076,17'd51513,17'd50863,17'd31288,17'd29330,17'd28460,17'd35372,17'd30220,17'd34833,17'd51602,17'd57183,17'd57184,17'd51693,17'd52134,17'd35100,17'd33095,17'd36214,17'd30220,17'd28945,17'd29071,17'd23855,17'd23168,17'd11959,17'd15053,17'd18917,17'd13135,17'd11958,17'd11958,17'd11958,17'd11960,17'd15053,17'd15053,17'd19158,17'd11396,17'd20610,17'd49324,17'd9047,17'd8105,17'd57555,17'd9351,17'd57318,17'd10994,17'd26039,17'd8884,17'd35515,17'd36778,17'd23859,17'd9189,17'd14383,17'd14928,17'd15180,17'd17237,17'd24862,17'd22133,17'd57556,17'd11815,17'd13143,17'd23186,17'd57557,17'd57558,17'd57559,17'd57560,17'd57561,17'd57562,17'd57563,17'd57564,17'd57197,17'd57565,17'd54131,17'd49182,17'd57453,17'd57566,17'd57567,17'd52428,17'd47934,17'd57568,17'd46425,17'd32496,17'd30586,17'd26902,17'd27259,17'd28482,17'd27767,17'd25565,17'd27513,17'd28599,17'd28717,17'd25177,17'd29103,17'd28850,17'd28594,17'd25949,17'd27515,17'd26903,17'd27515,17'd27514,17'd26903,17'd33792,17'd31351,17'd25708,17'd57569,17'd39283,17'd31856,17'd28480,17'd25568,17'd25320,17'd25320,17'd25178,17'd28369,17'd28721,17'd25565,17'd27638,17'd28719,17'd24744,17'd31033,17'd23566,17'd29830,17'd48257,17'd23566,17'd52887,17'd50899,17'd50899,17'd51554,17'd57570,17'd57571,17'd57572,17'd57573,17'd57574,17'd52822,17'd55438,17'd47534,17'd51645,17'd53911,17'd57575,17'd42885,17'd43695,17'd31351,17'd27766,17'd25317,17'd25438,17'd33484,17'd27512,17'd27764,17'd33951,17'd25568,17'd29101,17'd28850,17'd27512,17'd48036,17'd57333,17'd56290,17'd25709,17'd25317,17'd27765,17'd27765,17'd28130,17'd27765,17'd25567,17'd28369,17'd25317,17'd31366,17'd25177,17'd25032,17'd30277,17'd57576,17'd21705,17'd51922,17'd51238,17'd34617,17'd50274,17'd31832,17'd49991,17'd47071,17'd57577,17'd51319,17'd57578,17'd57579,17'd57580,17'd57581,17'd57582,17'd57583,17'd57584,17'd57585,17'd57586,17'd22209,17'd57587,17'd22743,17'd53731,17'd56530,17'd57588,17'd57589,17'd23455,17'd8911,17'd7162,17'd24798,17'd5608,17'd42910,17'd4995,17'd32552,17'd4840,17'd47174,17'd5327,17'd4687,17'd5002,17'd33368,17'd31717,17'd9091,17'd9091,17'd7499,17'd8780,17'd7668,17'd9091,17'd32073,17'd6390,17'd5763,17'd37432,17'd57590,17'd41459,17'd5001,17'd34333,17'd54003,17'd51177,17'd49897,17'd49296,17'd49104,17'd57348,17'd57591,17'd57592,17'd57593,17'd49707,17'd57594,17'd57595,17'd57225,17'd57596,17'd57597,17'd57598,17'd57599,17'd57600,17'd46589,17'd39175,17'd57601,17'd40557,17'd57602,17'd3045,17'd57231,17'd57356,17'd57357,17'd56316,17'd57603,17'd57233,17'd53798,17'd53798,17'd56211,17'd57604,17'd57605,17'd57606,17'd57607,17'd23813,17'd20862,17'd53593,17'd56781,17'd238,17'd451,17'd8014,17'd57608,17'd448,17'd55757,17'd632,17'd238,17'd243,17'd243,17'd57609,17'd31250,17'd1114,17'd625,17'd2392,17'd3391,17'd3895,17'd4085,17'd57610,17'd6582,17'd3246,17'd3591,17'd1825,17'd3390,17'd54240,17'd57611,17'd55758,17'd57612,17'd57613,17'd57614,17'd57615,17'd20708,17'd40560,17'd56433,17'd55368,17'd57490,17'd57370,17'd57616,17'd57617
},
'{
17'd10802,17'd10669,17'd3429,17'd3752,17'd2597,17'd1414,17'd17,17'd17,17'd18,17'd18,17'd18,17'd3905,17'd17,17'd1415,17'd1414,17'd2258,17'd1688,17'd1688,17'd57618,17'd2597,17'd2936,17'd2257,17'd468,17'd653,17'd980,17'd57619,17'd652,17'd288,17'd30,17'd1129,17'd469,17'd657,17'd472,17'd659,17'd474,17'd1131,17'd57620,17'd49,17'd57621,17'd56114,17'd56892,17'd57622,17'd57623,17'd1292,17'd57373,17'd57624,17'd57625,17'd57626,17'd1433,17'd57627,17'd57628,17'd21956,17'd2628,17'd57257,17'd4271,17'd4272,17'd57629,17'd39633,17'd55896,17'd57630,17'd21965,17'd12958,17'd10694,17'd7418,17'd13471,17'd15766,17'd10113,17'd9301,17'd57631,17'd12958,17'd9703,17'd9574,17'd22634,17'd12533,17'd7418,17'd8539,17'd52283,17'd52851,17'd53370,17'd55577,17'd57632,17'd47572,17'd17207,17'd57633,17'd22631,17'd32100,17'd57634,17'd57635,17'd57636,17'd56232,17'd53950,17'd55776,17'd57637,17'd57638,17'd57639,17'd57640,17'd57641,17'd56240,17'd57642,17'd56025,17'd57643,17'd57644,17'd57645,17'd56239,17'd57646,17'd57647,17'd57648,17'd57649,17'd57398,17'd57650,17'd57651,17'd57652,17'd57653,17'd57654,17'd57655,17'd57656,17'd57657,17'd57658,17'd57659,17'd57660,17'd57661,17'd57662,17'd6790,17'd55596,17'd57663,17'd57664,17'd57665,17'd57666,17'd57667,17'd57668,17'd57669,17'd57416,17'd57670,17'd57671,17'd57672,17'd57419,17'd57673,17'd57674,17'd57675,17'd15664,17'd57676,17'd11775,17'd12834,17'd57540,17'd57677,17'd13345,17'd57678,17'd57679,17'd12839,17'd57680,17'd57546,17'd57681,17'd57680,17'd57682,17'd57428,17'd57683,17'd57174,17'd57684,17'd12235,17'd57685,17'd55120,17'd53386,17'd57686,17'd57687,17'd54042,17'd18199,17'd55417,17'd55612,17'd55612,17'd57177,17'd57688,17'd55821,17'd31135,17'd57689,17'd35099,17'd32933,17'd30678,17'd30528,17'd36491,17'd33568,17'd52305,17'd50863,17'd51118,17'd31942,17'd31285,17'd28571,17'd29482,17'd36937,17'd34833,17'd52304,17'd52303,17'd52303,17'd52304,17'd52134,17'd35100,17'd31591,17'd34704,17'd30220,17'd28944,17'd28229,17'd23511,17'd23855,17'd12579,17'd17603,17'd18917,17'd15053,17'd11806,17'd12857,17'd12857,17'd12857,17'd13520,17'd13520,17'd17478,17'd25280,17'd21205,17'd15298,17'd35797,17'd57690,17'd8424,17'd12727,17'd24216,17'd15056,17'd57691,17'd22473,17'd12425,17'd8570,17'd24999,17'd15944,17'd11809,17'd33722,17'd15180,17'd17237,17'd11405,17'd57692,17'd10343,17'd24555,17'd55833,17'd57693,17'd57694,17'd57695,17'd57696,17'd57697,17'd57698,17'd57699,17'd57700,17'd57701,17'd57702,17'd54289,17'd48534,17'd56745,17'd57703,17'd57704,17'd57705,17'd40675,17'd46841,17'd46100,17'd33942,17'd36542,17'd27258,17'd28724,17'd27515,17'd26062,17'd25949,17'd26064,17'd28598,17'd27882,17'd28596,17'd25179,17'd25320,17'd28850,17'd28720,17'd26062,17'd27640,17'd27640,17'd26530,17'd25833,17'd33642,17'd28483,17'd27765,17'd33484,17'd33803,17'd28480,17'd28480,17'd27512,17'd25177,17'd25568,17'd25568,17'd27882,17'd25435,17'd28721,17'd25317,17'd28254,17'd24252,17'd31033,17'd23736,17'd32191,17'd37117,17'd29975,17'd30578,17'd57706,17'd57707,17'd57708,17'd57709,17'd57710,17'd57572,17'd57711,17'd57712,17'd51155,17'd57458,17'd47534,17'd50994,17'd57713,17'd53846,17'd41864,17'd42437,17'd31351,17'd25833,17'd28720,17'd25173,17'd24080,17'd25568,17'd28719,17'd27764,17'd27512,17'd28850,17'd39591,17'd25177,17'd57333,17'd33951,17'd28719,17'd28717,17'd28369,17'd27765,17'd27638,17'd28594,17'd28594,17'd28720,17'd27765,17'd27882,17'd25709,17'd31365,17'd39292,17'd57714,17'd38172,17'd57715,17'd57716,17'd57717,17'd43556,17'd50274,17'd31344,17'd57718,17'd35456,17'd57719,17'd57720,17'd35321,17'd57721,17'd57722,17'd57723,17'd27913,17'd56981,17'd26818,17'd57724,17'd57725,17'd20671,17'd57726,17'd56303,17'd22219,17'd57727,17'd22222,17'd23445,17'd23793,17'd23454,17'd6839,17'd24149,17'd5912,17'd24649,17'd6067,17'd4682,17'd4683,17'd4995,17'd47174,17'd4841,17'd5002,17'd4842,17'd5612,17'd6218,17'd6219,17'd9091,17'd10380,17'd10380,17'd10238,17'd7178,17'd5615,17'd5762,17'd5329,17'd57089,17'd57728,17'd49597,17'd55061,17'd55255,17'd52522,17'd57729,17'd49400,17'd51094,17'd55157,17'd57730,17'd57731,17'd57732,17'd49401,17'd57733,17'd57734,17'd57225,17'd57735,17'd57736,17'd57737,17'd57738,17'd45909,17'd57739,17'd39025,17'd39322,17'd57740,17'd57741,17'd44141,17'd57355,17'd57097,17'd57097,17'd57357,17'd56208,17'd57603,17'd57742,17'd57743,17'd56211,17'd56424,17'd55267,17'd53362,17'd2383,17'd35767,17'd57744,17'd52534,17'd31249,17'd792,17'd244,17'd793,17'd234,17'd8014,17'd238,17'd449,17'd450,17'd2418,17'd784,17'd450,17'd57609,17'd57745,17'd231,17'd229,17'd5371,17'd8185,17'd5940,17'd4559,17'd6581,17'd3391,17'd229,17'd228,17'd1825,17'd4228,17'd6405,17'd57746,17'd57747,17'd57748,17'd57749,17'd57750,17'd57751,17'd57752,17'd40560,17'd2381,17'd57753,17'd57754,17'd57755,17'd57756,17'd57757
},
'{
17'd10802,17'd10669,17'd3429,17'd3752,17'd2597,17'd2596,17'd1415,17'd17,17'd18,17'd18,17'd18,17'd3905,17'd17,17'd17,17'd1414,17'd2258,17'd1688,17'd1688,17'd57618,17'd2258,17'd2936,17'd2258,17'd290,17'd289,17'd652,17'd34669,17'd652,17'd288,17'd30,17'd1129,17'd982,17'd657,17'd472,17'd659,17'd986,17'd1131,17'd57000,17'd57758,17'd57759,17'd56674,17'd57002,17'd57622,17'd57372,17'd1292,17'd57113,17'd57760,17'd57761,17'd57762,17'd1296,17'd1566,17'd57375,17'd2133,17'd57763,17'd57257,17'd4271,17'd57764,17'd18642,17'd35489,17'd36186,17'd57765,17'd15523,17'd9575,17'd10694,17'd7418,17'd57766,17'd15766,17'd9301,17'd8067,17'd57767,17'd57631,17'd10113,17'd15517,17'd22119,17'd22633,17'd7418,17'd4611,17'd57768,17'd57769,17'd53522,17'd54254,17'd57382,17'd57770,17'd20585,17'd57771,17'd14219,17'd15767,17'd57635,17'd57772,17'd55483,17'd55483,17'd55577,17'd57773,17'd56574,17'd57774,17'd57775,17'd57776,17'd57509,17'd55583,17'd57276,17'd55777,17'd57777,17'd57778,17'd57779,17'd57780,17'd57781,17'd57782,17'd57783,17'd57784,17'd57785,17'd57786,17'd57282,17'd57787,17'd57788,17'd1602,17'd57789,17'd57790,17'd57143,17'd57791,17'd57792,17'd57793,17'd57794,17'd55595,17'd41333,17'd54631,17'd57795,17'd57796,17'd57667,17'd57797,17'd57666,17'd57798,17'd57799,17'd57800,17'd57670,17'd57535,17'd57801,17'd57802,17'd57803,17'd57804,17'd57805,17'd12832,17'd12227,17'd12691,17'd12692,17'd57540,17'd57806,17'd57677,17'd12694,17'd13232,17'd57807,17'd57808,17'd13234,17'd13234,17'd57809,17'd57810,17'd57811,17'd57812,17'd57813,17'd57814,17'd57815,17'd15675,17'd25404,17'd24850,17'd14126,17'd57816,17'd53775,17'd54278,17'd38503,17'd55612,17'd17844,17'd57177,17'd56946,17'd55942,17'd57817,17'd57689,17'd35099,17'd32933,17'd32926,17'd32926,17'd31773,17'd33568,17'd51272,17'd35239,17'd31589,17'd31127,17'd31440,17'd29645,17'd30220,17'd34704,17'd36936,17'd52134,17'd52304,17'd52134,17'd52304,17'd51513,17'd35100,17'd31591,17'd34704,17'd30220,17'd28461,17'd28229,17'd28107,17'd23855,17'd12108,17'd17474,17'd18197,17'd15053,17'd11806,17'd12857,17'd47110,17'd12112,17'd13520,17'd14379,17'd14382,17'd12583,17'd20610,17'd15298,17'd57818,17'd57819,17'd57820,17'd57821,17'd57822,17'd54046,17'd57823,17'd35930,17'd24711,17'd24368,17'd25677,17'd10174,17'd9479,17'd24998,17'd16553,17'd8724,17'd24863,17'd57824,17'd24549,17'd8588,17'd57825,17'd57826,17'd57827,17'd57828,17'd42262,17'd57829,17'd57830,17'd57831,17'd57832,17'd57833,17'd57834,17'd48451,17'd45368,17'd57835,17'd57836,17'd57837,17'd55138,17'd57838,17'd46435,17'd44358,17'd32496,17'd30735,17'd28853,17'd28724,17'd26174,17'd28481,17'd26062,17'd30606,17'd28597,17'd25177,17'd24896,17'd25031,17'd25179,17'd28850,17'd28594,17'd26062,17'd27515,17'd27640,17'd26530,17'd28602,17'd28721,17'd28484,17'd25177,17'd27512,17'd25568,17'd27512,17'd28719,17'd25568,17'd25709,17'd28480,17'd28717,17'd29970,17'd28600,17'd25317,17'd25178,17'd24416,17'd24086,17'd35865,17'd32008,17'd23217,17'd37386,17'd35865,17'd57839,17'd50648,17'd57840,17'd57841,17'd57842,17'd57843,17'd57844,17'd57845,17'd57846,17'd51155,17'd47638,17'd47339,17'd46554,17'd46202,17'd42299,17'd44478,17'd33478,17'd25707,17'd25708,17'd28594,17'd24079,17'd24080,17'd25177,17'd28719,17'd33803,17'd25709,17'd25317,17'd28369,17'd33484,17'd33803,17'd27512,17'd28717,17'd28369,17'd28130,17'd28720,17'd28720,17'd26064,17'd26064,17'd28598,17'd27765,17'd27882,17'd27882,17'd25951,17'd25569,17'd57847,17'd57848,17'd51633,17'd57849,17'd57850,17'd34617,17'd32665,17'd37534,17'd57851,17'd57852,17'd57853,17'd46773,17'd48997,17'd57854,17'd57855,17'd57856,17'd57582,17'd57857,17'd57858,17'd57859,17'd57860,17'd57861,17'd57862,17'd57863,17'd57864,17'd23626,17'd22222,17'd23445,17'd23972,17'd23454,17'd23974,17'd7324,17'd5323,17'd24649,17'd6067,17'd4682,17'd4683,17'd42910,17'd47174,17'd4686,17'd5002,17'd4842,17'd5158,17'd6218,17'd6219,17'd7499,17'd10380,17'd57865,17'd57866,17'd7178,17'd5614,17'd5333,17'd4686,17'd29595,17'd4998,17'd49597,17'd57867,17'd51931,17'd57868,17'd57869,17'd51012,17'd52355,17'd56205,17'd57730,17'd57870,17'd57871,17'd57872,17'd36738,17'd57873,17'd57874,17'd57875,17'd57876,17'd57877,17'd57878,17'd57879,17'd57880,17'd57881,17'd57882,17'd57883,17'd45182,17'd57741,17'd39623,17'd57884,17'd57097,17'd57357,17'd56208,17'd57603,17'd57742,17'd57743,17'd57743,17'd56211,17'd54511,17'd57885,17'd35205,17'd57886,17'd57887,17'd34510,17'd2419,17'd239,17'd244,17'd3100,17'd1122,17'd451,17'd36902,17'd955,17'd792,17'd24496,17'd35059,17'd450,17'd57609,17'd57888,17'd3098,17'd4880,17'd8185,17'd16382,17'd16382,17'd4714,17'd9123,17'd4729,17'd3246,17'd3246,17'd1824,17'd54163,17'd6405,17'd57889,17'd57747,17'd57890,17'd57891,17'd57892,17'd3219,17'd56548,17'd57106,17'd57359,17'd57893,17'd57894,17'd57895,17'd24161,17'd53800
},
'{
17'd10802,17'd10669,17'd3429,17'd3752,17'd2597,17'd1414,17'd17,17'd16,17'd18,17'd1128,17'd1128,17'd3905,17'd17,17'd17,17'd1414,17'd2425,17'd1831,17'd1831,17'd57618,17'd2426,17'd2596,17'd2425,17'd56331,17'd1692,17'd652,17'd2938,17'd653,17'd28,17'd468,17'd31,17'd982,17'd657,17'd57896,17'd473,17'd986,17'd40,17'd57000,17'd57897,17'd57621,17'd56674,17'd57002,17'd56892,17'd1151,17'd1152,17'd57898,17'd57899,17'd1156,17'd57762,17'd57900,17'd21025,17'd57495,17'd57901,17'd57902,17'd57903,17'd57904,17'd57905,17'd57906,17'd37050,17'd57907,17'd57119,17'd57908,17'd13844,17'd9703,17'd9440,17'd6300,17'd13972,17'd9301,17'd8067,17'd57631,17'd52027,17'd13470,17'd15898,17'd13471,17'd13722,17'd6143,17'd7582,17'd47975,17'd57909,17'd57910,17'd54350,17'd53685,17'd57911,17'd13721,17'd48297,17'd14768,17'd48189,17'd57013,17'd57634,17'd57912,17'd49303,17'd48819,17'd54172,17'd55093,17'd57913,17'd57914,17'd56806,17'd57639,17'd55782,17'd55579,17'd57915,17'd57916,17'd57917,17'd57918,17'd57919,17'd57920,17'd57646,17'd57921,17'd57922,17'd1321,17'd57923,17'd57924,17'd57282,17'd57140,17'd57925,17'd57926,17'd57927,17'd57928,17'd57929,17'd57930,17'd55791,17'd5712,17'd55393,17'd53307,17'd54031,17'd57931,17'd56710,17'd57932,17'd57933,17'd57666,17'd57798,17'd57934,17'd57935,17'd57936,17'd57937,17'd57938,17'd57939,17'd57940,17'd57804,17'd57941,17'd57675,17'd15664,17'd11491,17'd12079,17'd57942,17'd57806,17'd57943,17'd57944,17'd57945,17'd12387,17'd57807,17'd57946,17'd57947,17'd57948,17'd57949,17'd57949,17'd13118,17'd57950,17'd57309,17'd57814,17'd57951,17'd57685,17'd21976,17'd22988,17'd14663,17'd53541,17'd57952,17'd57953,17'd55612,17'd17844,17'd56497,17'd56946,17'd55942,17'd31135,17'd57689,17'd35099,17'd32597,17'd32926,17'd32926,17'd57061,17'd33095,17'd50863,17'd35239,17'd31589,17'd30973,17'd29330,17'd28686,17'd30073,17'd34835,17'd53250,17'd51513,17'd34044,17'd34044,17'd52134,17'd34044,17'd33882,17'd56619,17'd34704,17'd30220,17'd28686,17'd28818,17'd27121,17'd18200,17'd12108,17'd12106,17'd12719,17'd11958,17'd12857,17'd12857,17'd47110,17'd12999,17'd15185,17'd14379,17'd14382,17'd25280,17'd21205,17'd15298,17'd57818,17'd7950,17'd19781,17'd57954,17'd57955,17'd12589,17'd57956,17'd37334,17'd21987,17'd15429,17'd8569,17'd8873,17'd9345,17'd34204,17'd17964,17'd8724,17'd11405,17'd57692,17'd10748,17'd26042,17'd16452,17'd57693,17'd57694,17'd57957,17'd57958,17'd57959,17'd57960,17'd57961,17'd57962,17'd57963,17'd57964,17'd48261,17'd52505,17'd57965,17'd56857,17'd57966,17'd52428,17'd50995,17'd49275,17'd43424,17'd32343,17'd28486,17'd28725,17'd26903,17'd26062,17'd27767,17'd26064,17'd28598,17'd25709,17'd28254,17'd28595,17'd32007,17'd25179,17'd29244,17'd27765,17'd28602,17'd26174,17'd25708,17'd28720,17'd25567,17'd27882,17'd25568,17'd28719,17'd28254,17'd25568,17'd27512,17'd27512,17'd25568,17'd28717,17'd33484,17'd25438,17'd29825,17'd28369,17'd27512,17'd24417,17'd30879,17'd23566,17'd29828,17'd37117,17'd37117,17'd23923,17'd33950,17'd57967,17'd52161,17'd50899,17'd57968,17'd57969,17'd57970,17'd57971,17'd57845,17'd57571,17'd49374,17'd54059,17'd51475,17'd50266,17'd57972,17'd42597,17'd43695,17'd35012,17'd26174,17'd28602,17'd28598,17'd25709,17'd25709,17'd25709,17'd28480,17'd28480,17'd28369,17'd25317,17'd28717,17'd28480,17'd33484,17'd28717,17'd28369,17'd28484,17'd28600,17'd28720,17'd28723,17'd28602,17'd30606,17'd38671,17'd27765,17'd29103,17'd31034,17'd25436,17'd57973,17'd32190,17'd34615,17'd54207,17'd57974,17'd35293,17'd57975,17'd54662,17'd48914,17'd48712,17'd57976,17'd57977,17'd45886,17'd57978,17'd49893,17'd57979,17'd57980,17'd57981,17'd57982,17'd57983,17'd57984,17'd57985,17'd57986,17'd35047,17'd29154,17'd22392,17'd23624,17'd22222,17'd23445,17'd23972,17'd23454,17'd8911,17'd7658,17'd5912,17'd24649,17'd5145,17'd4839,17'd4995,17'd5153,17'd5327,17'd4686,17'd5005,17'd4842,17'd5331,17'd6218,17'd6220,17'd7668,17'd10380,17'd10238,17'd50283,17'd6853,17'd5336,17'd33692,17'd42910,17'd47470,17'd55350,17'd55061,17'd57867,17'd57987,17'd52604,17'd38195,17'd52764,17'd52450,17'd56538,17'd57988,17'd57989,17'd57990,17'd4205,17'd57991,17'd50082,17'd57992,17'd57993,17'd47377,17'd57994,17'd55872,17'd57879,17'd57880,17'd53584,17'd57995,17'd57996,17'd57881,17'd42472,17'd43461,17'd57997,17'd57998,17'd56774,17'd56208,17'd57742,17'd57999,17'd58000,17'd58000,17'd56211,17'd54511,17'd58001,17'd58002,17'd1807,17'd38714,17'd58003,17'd18386,17'd450,17'd1681,17'd3100,17'd1122,17'd238,17'd58004,17'd635,17'd635,17'd635,17'd621,17'd634,17'd31726,17'd1114,17'd1401,17'd5372,17'd5630,17'd14586,17'd16256,17'd9123,17'd5776,17'd4713,17'd4575,17'd3897,17'd4558,17'd18143,17'd6405,17'd55078,17'd58005,17'd57891,17'd58006,17'd58007,17'd58008,17'd58009,17'd58010,17'd58011,17'd58012,17'd57894,17'd58013,17'd58014,17'd53800
},
'{
17'd10669,17'd10669,17'd3429,17'd3752,17'd2596,17'd1414,17'd17,17'd16,17'd18,17'd1128,17'd1128,17'd1128,17'd3905,17'd17,17'd1414,17'd2257,17'd1831,17'd1831,17'd12194,17'd2426,17'd2597,17'd2258,17'd58015,17'd1692,17'd653,17'd2938,17'd653,17'd29,17'd809,17'd31,17'd982,17'd984,17'd57896,17'd58016,17'd986,17'd14599,17'd477,17'd478,17'd57759,17'd56674,17'd56333,17'd56892,17'd1151,17'd1152,17'd1562,17'd57899,17'd58017,17'd58018,17'd58019,17'd1435,17'd21331,17'd58020,17'd58021,17'd58022,17'd57257,17'd57764,17'd58023,17'd58024,17'd36753,17'd56564,17'd58025,17'd15523,17'd23837,17'd13972,17'd6301,17'd9300,17'd9301,17'd8066,17'd8372,17'd13467,17'd13466,17'd23837,17'd13845,17'd13846,17'd6143,17'd9440,17'd48301,17'd58026,17'd58027,17'd58028,17'd58029,17'd58030,17'd14624,17'd14219,17'd14626,17'd48189,17'd56900,17'd58031,17'd48820,17'd57013,17'd55668,17'd57773,17'd58032,17'd58033,17'd58034,17'd56696,17'd58035,17'd56912,17'd55579,17'd56913,17'd58036,17'd58037,17'd58038,17'd58039,17'd58040,17'd57646,17'd58041,17'd58042,17'd58043,17'd58044,17'd58045,17'd58046,17'd58047,17'd58048,17'd58049,17'd58050,17'd58051,17'd58052,17'd58053,17'd58054,17'd58055,17'd58056,17'd56255,17'd42216,17'd58057,17'd58058,17'd57414,17'd57932,17'd58059,17'd58059,17'd58060,17'd58061,17'd58062,17'd58063,17'd58064,17'd58065,17'd57940,17'd57803,17'd58066,17'd57805,17'd12226,17'd12690,17'd58067,17'd57806,17'd58068,17'd57943,17'd57677,17'd58069,17'd57945,17'd12387,17'd57807,17'd58070,17'd58071,17'd58071,17'd57946,17'd58072,17'd11781,17'd57950,17'd57813,17'd58073,17'd12235,17'd13507,17'd53973,17'd58074,17'd53467,17'd58075,17'd58076,17'd56272,17'd17844,17'd56497,17'd56947,17'd55942,17'd58077,17'd57180,17'd32926,17'd32597,17'd30528,17'd32597,17'd57061,17'd33095,17'd50863,17'd35239,17'd35093,17'd31287,17'd30072,17'd28686,17'd30073,17'd34835,17'd53250,17'd51603,17'd35100,17'd34044,17'd52134,17'd51603,17'd53250,17'd56619,17'd34704,17'd30220,17'd28686,17'd28818,17'd27121,17'd18084,17'd12254,17'd17348,17'd17603,17'd11958,17'd12420,17'd12857,17'd12105,17'd12999,17'd15185,17'd14264,17'd14382,17'd25280,17'd21205,17'd15298,17'd23341,17'd16566,17'd15949,17'd58078,17'd58079,17'd16077,17'd25412,17'd23342,17'd21987,17'd11404,17'd8724,17'd8720,17'd9344,17'd33083,17'd15430,17'd8724,17'd24713,17'd15947,17'd24551,17'd55125,17'd16452,17'd58080,17'd58081,17'd58082,17'd58083,17'd58084,17'd56178,17'd58085,17'd58086,17'd58087,17'd58088,17'd54131,17'd49090,17'd57965,17'd57837,17'd58089,17'd58090,17'd47049,17'd46203,17'd44590,17'd33163,17'd26781,17'd28725,17'd27515,17'd28481,17'd27513,17'd30606,17'd31055,17'd25709,17'd28596,17'd28718,17'd25032,17'd25179,17'd25320,17'd27882,17'd28720,17'd32658,17'd28721,17'd27765,17'd28717,17'd27512,17'd25029,17'd25029,17'd28254,17'd28719,17'd25568,17'd25568,17'd28719,17'd28480,17'd27882,17'd28850,17'd27511,17'd25178,17'd24744,17'd29100,17'd34137,17'd29686,17'd37117,17'd37117,17'd36987,17'd29099,17'd58091,17'd56285,17'd57196,17'd58092,17'd58093,17'd58094,17'd50645,17'd58095,17'd57844,17'd53989,17'd58096,17'd58097,17'd56639,17'd50566,17'd55335,17'd44699,17'd49273,17'd27766,17'd28602,17'd28594,17'd28597,17'd31366,17'd25709,17'd25709,17'd33484,17'd25709,17'd28484,17'd25317,17'd33484,17'd28480,17'd25709,17'd27882,17'd28130,17'd28600,17'd28130,17'd28720,17'd28723,17'd28602,17'd27513,17'd30734,17'd25567,17'd41730,17'd33318,17'd31521,17'd39450,17'd43842,17'd34616,17'd46455,17'd52251,17'd34881,17'd58098,17'd48279,17'd58099,17'd58100,17'd58101,17'd58102,17'd58103,17'd24097,17'd58104,17'd58105,17'd58106,17'd58107,17'd58108,17'd58109,17'd33685,17'd58110,17'd58111,17'd22057,17'd29424,17'd30483,17'd23624,17'd23445,17'd23445,17'd23453,17'd23454,17'd24149,17'd6702,17'd24649,17'd24798,17'd5145,17'd4682,17'd5153,17'd5153,17'd4841,17'd4686,17'd4842,17'd5004,17'd6218,17'd8303,17'd7499,17'd8780,17'd10380,17'd50283,17'd52094,17'd53214,17'd5335,17'd4845,17'd30485,17'd58112,17'd49704,17'd56532,17'd49997,17'd57987,17'd58113,17'd56877,17'd49297,17'd52186,17'd52766,17'd58114,17'd57989,17'd58115,17'd57991,17'd57991,17'd58116,17'd58117,17'd58118,17'd58119,17'd58120,17'd53737,17'd39025,17'd39025,17'd58121,17'd57882,17'd58122,17'd58123,17'd53584,17'd42472,17'd42642,17'd58124,17'd56421,17'd58125,17'd57742,17'd57999,17'd58000,17'd58000,17'd58126,17'd54419,17'd58001,17'd58127,17'd58128,17'd35906,17'd58129,17'd36323,17'd238,17'd1681,17'd609,17'd1257,17'd800,17'd58130,17'd636,17'd454,17'd636,17'd955,17'd452,17'd31726,17'd232,17'd445,17'd1946,17'd3073,17'd5631,17'd16256,17'd5776,17'd7365,17'd4730,17'd5789,17'd5373,17'd5937,17'd54779,17'd6237,17'd55078,17'd57889,17'd58006,17'd58131,17'd50002,17'd3218,17'd3067,17'd2900,17'd35904,17'd58132,17'd58133,17'd58013,17'd58134,17'd58135
},
'{
17'd52621,17'd3429,17'd3429,17'd3752,17'd2596,17'd1414,17'd16,17'd18,17'd1128,17'd11,17'd11,17'd1128,17'd3905,17'd17,17'd1414,17'd2257,17'd2597,17'd2258,17'd52621,17'd52621,17'd3752,17'd2258,17'd58015,17'd56331,17'd2938,17'd2938,17'd653,17'd652,17'd289,17'd31,17'd982,17'd1130,17'd57896,17'd58016,17'd986,17'd15362,17'd816,17'd478,17'd57759,17'd56675,17'd58136,17'd56892,17'd1151,17'd57372,17'd58137,17'd58138,17'd58139,17'd58018,17'd58019,17'd1298,17'd58140,17'd58141,17'd1991,17'd21640,17'd34171,17'd57764,17'd58023,17'd58142,17'd58143,17'd58144,17'd58145,17'd58146,17'd15645,17'd13469,17'd58147,17'd8538,17'd9007,17'd9704,17'd13842,17'd14100,17'd14100,17'd58148,17'd13328,17'd9440,17'd6143,17'd13846,17'd9704,17'd48300,17'd58027,17'd54094,17'd54254,17'd53447,17'd56340,17'd14624,17'd15641,17'd48080,17'd57123,17'd55668,17'd58149,17'd57013,17'd55576,17'd58150,17'd58151,17'd58152,17'd58034,17'd58153,17'd56696,17'd56132,17'd56132,17'd56239,17'd58154,17'd58155,17'd58156,17'd58157,17'd58158,17'd58159,17'd56909,17'd58160,17'd55784,17'd58161,17'd58162,17'd58163,17'd58164,17'd58165,17'd58166,17'd58167,17'd58168,17'd58169,17'd58170,17'd58171,17'd58172,17'd58173,17'd58174,17'd41925,17'd58175,17'd55504,17'd56711,17'd58176,17'd58177,17'd58178,17'd58059,17'd58060,17'd58179,17'd58180,17'd58181,17'd58182,17'd58183,17'd57940,17'd58184,17'd57941,17'd58185,17'd12226,17'd14501,17'd58186,17'd58068,17'd58187,17'd58068,17'd58188,17'd57944,17'd57945,17'd58189,17'd58190,17'd58191,17'd58192,17'd58193,17'd58194,17'd12554,17'd12839,17'd13118,17'd57813,17'd57684,17'd12706,17'd20305,17'd23844,17'd52950,17'd56159,17'd55416,17'd56947,17'd56161,17'd56616,17'd56616,17'd39661,17'd58077,17'd58195,17'd58196,17'd58195,17'd32597,17'd37985,17'd57061,17'd33095,17'd50863,17'd35239,17'd35093,17'd30973,17'd29067,17'd28686,17'd30073,17'd34381,17'd33243,17'd35100,17'd33243,17'd34044,17'd51513,17'd51432,17'd33243,17'd56619,17'd34704,17'd30220,17'd29481,17'd28572,17'd26629,17'd18084,17'd12254,17'd17348,17'd12106,17'd12420,17'd12420,17'd12857,17'd12105,17'd12999,17'd15185,17'd14264,17'd11522,17'd25280,17'd26037,17'd15298,17'd10607,17'd8253,17'd14390,17'd53835,17'd15572,17'd15689,17'd22648,17'd11138,17'd9196,17'd17481,17'd8725,17'd9044,17'd9346,17'd16065,17'd15430,17'd8725,17'd24713,17'd15947,17'd24551,17'd18924,17'd12870,17'd23186,17'd58197,17'd58198,17'd58199,17'd58200,17'd58201,17'd58202,17'd58203,17'd58204,17'd58205,17'd45368,17'd57835,17'd56857,17'd44820,17'd48359,17'd47044,17'd48524,17'd58206,17'd43020,17'd27372,17'd26782,17'd28725,17'd27514,17'd27767,17'd27513,17'd28599,17'd33484,17'd29244,17'd24896,17'd24417,17'd30126,17'd29533,17'd29976,17'd25177,17'd25317,17'd29970,17'd29101,17'd25177,17'd25029,17'd25029,17'd25029,17'd25029,17'd27637,17'd28719,17'd25568,17'd27512,17'd28719,17'd25177,17'd29101,17'd29103,17'd25030,17'd24744,17'd24415,17'd34137,17'd29374,17'd23216,17'd23216,17'd36987,17'd29830,17'd23920,17'd53556,17'd50563,17'd58207,17'd58208,17'd58209,17'd58210,17'd58211,17'd58212,17'd57574,17'd49571,17'd54132,17'd56639,17'd56512,17'd50264,17'd48258,17'd45036,17'd33643,17'd28720,17'd28720,17'd27638,17'd28597,17'd33000,17'd28597,17'd33000,17'd28597,17'd27765,17'd27765,17'd27882,17'd33484,17'd31366,17'd28597,17'd25567,17'd28600,17'd25435,17'd28720,17'd28720,17'd28723,17'd26064,17'd30734,17'd27638,17'd28597,17'd28484,17'd33483,17'd38978,17'd32351,17'd58213,17'd33946,17'd58214,17'd46456,17'd58215,17'd58216,17'd58217,17'd58218,17'd58219,17'd58220,17'd58221,17'd58222,17'd58223,17'd58224,17'd58225,17'd58226,17'd58227,17'd58228,17'd58229,17'd20672,17'd58230,17'd22383,17'd55058,17'd58231,17'd23621,17'd23624,17'd23445,17'd23625,17'd23453,17'd23278,17'd6543,17'd7324,17'd53352,17'd53352,17'd6067,17'd5145,17'd4996,17'd4995,17'd4686,17'd4841,17'd28418,17'd5335,17'd6219,17'd9091,17'd7668,17'd9933,17'd7499,17'd36586,17'd31717,17'd28185,17'd5330,17'd4686,17'd57728,17'd47470,17'd4369,17'd49805,17'd38445,17'd52604,17'd37562,17'd57594,17'd57731,17'd58232,17'd58233,17'd37564,17'd49003,17'd58234,17'd57734,17'd56771,17'd58235,17'd58236,17'd47083,17'd58237,17'd58238,17'd58239,17'd57881,17'd57741,17'd58121,17'd58122,17'd41309,17'd42040,17'd58240,17'd42642,17'd57997,17'd56315,17'd56208,17'd58125,17'd53798,17'd58241,17'd58000,17'd57234,17'd56212,17'd57482,17'd57242,17'd58242,17'd24495,17'd38457,17'd36322,17'd35059,17'd243,17'd961,17'd1122,17'd799,17'd955,17'd58243,17'd455,17'd455,17'd635,17'd955,17'd1540,17'd31250,17'd427,17'd2392,17'd2097,17'd6889,17'd5631,17'd58244,17'd5029,17'd4714,17'd6581,17'd5789,17'd37708,17'd56549,17'd6238,17'd6237,17'd55078,17'd57889,17'd58245,17'd58246,17'd58247,17'd40999,17'd39324,17'd21783,17'd58248,17'd58249,17'd58250,17'd58251,17'd58252,17'd58253
},
'{
17'd52621,17'd3429,17'd3429,17'd2597,17'd2257,17'd1414,17'd17,17'd18,17'd1128,17'd11,17'd11,17'd1128,17'd3905,17'd3905,17'd1416,17'd2257,17'd2597,17'd2258,17'd3429,17'd10547,17'd3429,17'd3752,17'd58254,17'd58015,17'd468,17'd2938,17'd653,17'd652,17'd29,17'd30,17'd291,17'd1130,17'd57896,17'd15118,17'd986,17'd15362,17'd815,17'd298,17'd58255,17'd58256,17'd57110,17'd57002,17'd1151,17'd57372,17'd58137,17'd57899,17'd58257,17'd57762,17'd1158,17'd1298,17'd1565,17'd58258,17'd57628,17'd58021,17'd58259,17'd58260,17'd58023,17'd57378,17'd58261,17'd58262,17'd58263,17'd58264,17'd58265,17'd13844,17'd7582,17'd7750,17'd8538,17'd9704,17'd13842,17'd14099,17'd48300,17'd58266,17'd58267,17'd58268,17'd7418,17'd13846,17'd58268,17'd58269,17'd52851,17'd53522,17'd58270,17'd54254,17'd57012,17'd58271,17'd47865,17'd48080,17'd56343,17'd53685,17'd58149,17'd57504,17'd58272,17'd58150,17'd58273,17'd55907,17'd58274,17'd58275,17'd56239,17'd57516,17'd57390,17'd58276,17'd58277,17'd58278,17'd58279,17'd58280,17'd58281,17'd56696,17'd58282,17'd58283,17'd1460,17'd58284,17'd57398,17'd58285,17'd57283,17'd58286,17'd58287,17'd58288,17'd58289,17'd4796,17'd58290,17'd58291,17'd58292,17'd58293,17'd54906,17'd44522,17'd51104,17'd54545,17'd55505,17'd58294,17'd58177,17'd58178,17'd58295,17'd58177,17'd58177,17'd58060,17'd58296,17'd58297,17'd58298,17'd58299,17'd58300,17'd58301,17'd58302,17'd58303,17'd58304,17'd13621,17'd58305,17'd58187,17'd58306,17'd58306,17'd58188,17'd58307,17'd13346,17'd13116,17'd58190,17'd58308,17'd58309,17'd58310,17'd57807,17'd12696,17'd12978,17'd13625,17'd56943,17'd13242,17'd12849,17'd12244,17'd24986,17'd58311,17'd57551,17'd56497,17'd56161,17'd56161,17'd56161,17'd39661,17'd58312,17'd58195,17'd58313,17'd58196,17'd32766,17'd36214,17'd58314,17'd33243,17'd50863,17'd35239,17'd35093,17'd32283,17'd34551,17'd28686,17'd29785,17'd34381,17'd33243,17'd53250,17'd33095,17'd34047,17'd51432,17'd35100,17'd33095,17'd54732,17'd31773,17'd29646,17'd29481,17'd28572,17'd27737,17'd26758,17'd23855,17'd19407,17'd17474,17'd16321,17'd12419,17'd12420,17'd12259,17'd11957,17'd19158,17'd14264,17'd11396,17'd25280,17'd26037,17'd15298,17'd12264,17'd8253,17'd16078,17'd58315,17'd53635,17'd12727,17'd18203,17'd25679,17'd8578,17'd9349,17'd8726,17'd9621,17'd9743,17'd25408,17'd15430,17'd8724,17'd13257,17'd58316,17'd22478,17'd25537,17'd12870,17'd58317,17'd58318,17'd58319,17'd58320,17'd58321,17'd58322,17'd58323,17'd58324,17'd58325,17'd58326,17'd54841,17'd56857,17'd45606,17'd55332,17'd48621,17'd54748,17'd46326,17'd41864,17'd52336,17'd27146,17'd26902,17'd28725,17'd25949,17'd30606,17'd28598,17'd31520,17'd27512,17'd29976,17'd24417,17'd24742,17'd28851,17'd34276,17'd25180,17'd27512,17'd25177,17'd25320,17'd25178,17'd25029,17'd28974,17'd24898,17'd25030,17'd28254,17'd27637,17'd25177,17'd28719,17'd27512,17'd25177,17'd29244,17'd29244,17'd25178,17'd24745,17'd24090,17'd23918,17'd23923,17'd23216,17'd30425,17'd29973,17'd29975,17'd23386,17'd29528,17'd53556,17'd56285,17'd58327,17'd58328,17'd50645,17'd58329,17'd50814,17'd58330,17'd54941,17'd58331,17'd58332,17'd57330,17'd58333,17'd48258,17'd43017,17'd43550,17'd28600,17'd28594,17'd28594,17'd25567,17'd28597,17'd28597,17'd28597,17'd33000,17'd27765,17'd28130,17'd25567,17'd25709,17'd25709,17'd28597,17'd28597,17'd28130,17'd25435,17'd28723,17'd28723,17'd28723,17'd25566,17'd28602,17'd27638,17'd25567,17'd27765,17'd28484,17'd29533,17'd58334,17'd52752,17'd43427,17'd47839,17'd58335,17'd58336,17'd58337,17'd58338,17'd58339,17'd58340,17'd44242,17'd44832,17'd58341,17'd36011,17'd58342,17'd58343,17'd58344,17'd58345,17'd58346,17'd58347,17'd58348,17'd20821,17'd58349,17'd22745,17'd29021,17'd22391,17'd56875,17'd58350,17'd23445,17'd23972,17'd23107,17'd23279,17'd7658,17'd7324,17'd53352,17'd53352,17'd5145,17'd38442,17'd30486,17'd4683,17'd4686,17'd28418,17'd30180,17'd27935,17'd9091,17'd9091,17'd27696,17'd9933,17'd32073,17'd31717,17'd30638,17'd5160,17'd4845,17'd5155,17'd47660,17'd39938,17'd52183,17'd54499,17'd52688,17'd58351,17'd58352,17'd58353,17'd49105,17'd58354,17'd58355,17'd58356,17'd58357,17'd3847,17'd57991,17'd56659,17'd58358,17'd58359,17'd58360,17'd58361,17'd58362,17'd58363,17'd57881,17'd58364,17'd58123,17'd45780,17'd41309,17'd44266,17'd42472,17'd57355,17'd57097,17'd58365,17'd58366,17'd58125,17'd53798,17'd58241,17'd58000,17'd56321,17'd56002,17'd58367,17'd58368,17'd1662,17'd58369,17'd58129,17'd36455,17'd36748,17'd630,17'd793,17'd234,17'd244,17'd955,17'd58370,17'd455,17'd455,17'd635,17'd792,17'd245,17'd31100,17'd954,17'd1810,17'd3073,17'd4714,17'd35060,17'd58244,17'd11335,17'd7537,17'd6094,17'd5789,17'd37821,17'd58371,17'd6238,17'd6237,17'd55078,17'd57889,17'd58372,17'd9245,17'd51580,17'd58373,17'd58374,17'd52360,17'd57606,17'd58375,17'd58250,17'd58376,17'd58377,17'd58378
},
'{
17'd3429,17'd3429,17'd2597,17'd2597,17'd2257,17'd1414,17'd17,17'd18,17'd1128,17'd11,17'd10,17'd1128,17'd3905,17'd3905,17'd17,17'd1414,17'd2597,17'd2258,17'd3429,17'd10547,17'd3429,17'd3752,17'd57618,17'd57493,17'd1692,17'd468,17'd2938,17'd653,17'd29,17'd809,17'd291,17'd32,17'd57896,17'd15118,17'd58016,17'd986,17'd41,17'd819,17'd58379,17'd58380,17'd56792,17'd57002,17'd57372,17'd57372,17'd58381,17'd1562,17'd58382,17'd57626,17'd58383,17'd58384,17'd58385,17'd1713,17'd58386,17'd58387,17'd57763,17'd3769,17'd4445,17'd58388,17'd58389,17'd58390,17'd58144,17'd58145,17'd58391,17'd21965,17'd8538,17'd5409,17'd7582,17'd13469,17'd13842,17'd14623,17'd48300,17'd58392,17'd58393,17'd8539,17'd9159,17'd8537,17'd5410,17'd58394,17'd58395,17'd58396,17'd53608,17'd58397,17'd53370,17'd48078,17'd47865,17'd47972,17'd57012,17'd48821,17'd55773,17'd58398,17'd58399,17'd58400,17'd55185,17'd58401,17'd58402,17'd58403,17'd58404,17'd58405,17'd58159,17'd56579,17'd58406,17'd55905,17'd58279,17'd58407,17'd56350,17'd57516,17'd58159,17'd58408,17'd58409,17'd58410,17'd57135,17'd58411,17'd58412,17'd58413,17'd57285,17'd58414,17'd58415,17'd58416,17'd58417,17'd58418,17'd58419,17'd58420,17'd58421,17'd58422,17'd51023,17'd54102,17'd56043,17'd58423,17'd58179,17'd58178,17'd58295,17'd58424,17'd58424,17'd58177,17'd58425,17'd58426,17'd58298,17'd58299,17'd58427,17'd58428,17'd58429,17'd58430,17'd58431,17'd14791,17'd58432,17'd58305,17'd58433,17'd58434,17'd58435,17'd58188,17'd58436,17'd58437,17'd58438,17'd58439,17'd58440,17'd58441,17'd58442,17'd58443,17'd58443,17'd58444,17'd58445,17'd57049,17'd12558,17'd18189,17'd22294,17'd53182,17'd55819,17'd57953,17'd56161,17'd55699,17'd56161,17'd39661,17'd58312,17'd58446,17'd58447,17'd58447,17'd58448,17'd58446,17'd31597,17'd33243,17'd51118,17'd35239,17'd35644,17'd34704,17'd28686,17'd29645,17'd30220,17'd34381,17'd33243,17'd53250,17'd54926,17'd33243,17'd35100,17'd53250,17'd33095,17'd54732,17'd31773,17'd29646,17'd29481,17'd28572,17'd28104,17'd26758,17'd23855,17'd14807,17'd16321,17'd16321,17'd12419,17'd12857,17'd11957,17'd11962,17'd19158,17'd14264,17'd11396,17'd10990,17'd25928,17'd33083,17'd8409,17'd16566,17'd19536,17'd58449,17'd10862,17'd14938,17'd8254,17'd8250,17'd8417,17'd17126,17'd8409,17'd8881,17'd8874,17'd25814,17'd15430,17'd8724,17'd13257,17'd58316,17'd8586,17'd10864,17'd23528,17'd58450,17'd58451,17'd58452,17'd58453,17'd58454,17'd58455,17'd58456,17'd58457,17'd50261,17'd48251,17'd57837,17'd56857,17'd58458,17'd51557,17'd55438,17'd48523,17'd46203,17'd44590,17'd33154,17'd27146,17'd27258,17'd28724,17'd26062,17'd30606,17'd28597,17'd49481,17'd25029,17'd25032,17'd28601,17'd23916,17'd34467,17'd28368,17'd25032,17'd28596,17'd27764,17'd24897,17'd24898,17'd24896,17'd24896,17'd24898,17'd25030,17'd28254,17'd27637,17'd25568,17'd27764,17'd27637,17'd25320,17'd29976,17'd25032,17'd24744,17'd34467,17'd31502,17'd30128,17'd23216,17'd41273,17'd30425,17'd29973,17'd29686,17'd31502,17'd29527,17'd58459,17'd52887,17'd58460,17'd58461,17'd58462,17'd58463,17'd58464,17'd57573,17'd58465,17'd54203,17'd54575,17'd50152,17'd48258,17'd43155,17'd44359,17'd28130,17'd27765,17'd28130,17'd28130,17'd28597,17'd28597,17'd25567,17'd28597,17'd25567,17'd28130,17'd28130,17'd25567,17'd25709,17'd25709,17'd25567,17'd25567,17'd28720,17'd28720,17'd33333,17'd26402,17'd33970,17'd33970,17'd33009,17'd30456,17'd27765,17'd29970,17'd27882,17'd34276,17'd45746,17'd41729,17'd21695,17'd58466,17'd58467,17'd58468,17'd58469,17'd25182,17'd58470,17'd58471,17'd58472,17'd44123,17'd58473,17'd58474,17'd58475,17'd58476,17'd58477,17'd58107,17'd58478,17'd57585,17'd20820,17'd58479,17'd21594,17'd58480,17'd56304,17'd23268,17'd57588,17'd57589,17'd23973,17'd23972,17'd58481,17'd8289,17'd24477,17'd5322,17'd5144,17'd5145,17'd5144,17'd38442,17'd5153,17'd4683,17'd5328,17'd28418,17'd25627,17'd27935,17'd9091,17'd32074,17'd9933,17'd29740,17'd37152,17'd31891,17'd5160,17'd5329,17'd4847,17'd34657,17'd55645,17'd39016,17'd53580,17'd50672,17'd58113,17'd37562,17'd49898,17'd57094,17'd58356,17'd3542,17'd58482,17'd58483,17'd58484,17'd3847,17'd58485,17'd57591,17'd58486,17'd55556,17'd58487,17'd57601,17'd58488,17'd40095,17'd58489,17'd58490,17'd41154,17'd58491,17'd58492,17'd44266,17'd42472,17'd57355,17'd57097,17'd56207,17'd58125,17'd58125,17'd58241,17'd58126,17'd56321,17'd55267,17'd2070,17'd32402,17'd58493,17'd58494,17'd58495,17'd58129,17'd56215,17'd3071,17'd235,17'd447,17'd429,17'd245,17'd955,17'd454,17'd455,17'd637,17'd592,17'd634,17'd1093,17'd233,17'd1680,17'd7210,17'd14178,17'd16256,17'd35060,17'd58496,17'd11336,17'd9544,17'd6891,17'd4730,17'd5939,17'd58497,17'd6238,17'd6237,17'd58498,17'd57889,17'd58372,17'd55166,17'd50496,17'd37819,17'd2900,17'd58499,17'd58500,17'd58501,17'd58250,17'd58502,17'd58376,17'd58378
},
'{
17'd3429,17'd3429,17'd2597,17'd2597,17'd2257,17'd1414,17'd17,17'd18,17'd1128,17'd11,17'd10,17'd11,17'd3905,17'd3905,17'd17,17'd1416,17'd2257,17'd2426,17'd3429,17'd12195,17'd52621,17'd3429,17'd58503,17'd12194,17'd290,17'd468,17'd468,17'd653,17'd29,17'd289,17'd2599,17'd2259,17'd16011,17'd15118,17'd58016,17'd58504,17'd15497,17'd58505,17'd48,17'd58380,17'd56674,17'd56672,17'd57002,17'd57372,17'd58506,17'd78,17'd58382,17'd58507,17'd58508,17'd58509,17'd58510,17'd18518,17'd58511,17'd16639,17'd57763,17'd58512,17'd4445,17'd57497,17'd58513,17'd58514,17'd58262,17'd58515,17'd58025,17'd58516,17'd9007,17'd5409,17'd8537,17'd13469,17'd13842,17'd58394,17'd58392,17'd58026,17'd58517,17'd7751,17'd12534,17'd8537,17'd6463,17'd58267,17'd57769,17'd53448,17'd53523,17'd58518,17'd58519,17'd58520,17'd48079,17'd47971,17'd52932,17'd49200,17'd49303,17'd57502,17'd58399,17'd58521,17'd55900,17'd58522,17'd56023,17'd58523,17'd58524,17'd58525,17'd55378,17'd55378,17'd58406,17'd58526,17'd58279,17'd58527,17'd56807,17'd58528,17'd58282,17'd58529,17'd1459,17'd58530,17'd58531,17'd58532,17'd58533,17'd58534,17'd58535,17'd58536,17'd58537,17'd58538,17'd58539,17'd58540,17'd58541,17'd58542,17'd58543,17'd58544,17'd54266,17'd54908,17'd58545,17'd56712,17'd58546,17'd58547,17'd58548,17'd58549,17'd58424,17'd58177,17'd58425,17'd58550,17'd58551,17'd58552,17'd58553,17'd58554,17'd58555,17'd58556,17'd58557,17'd14240,17'd58558,17'd58559,17'd58433,17'd58434,17'd58560,17'd58435,17'd58561,17'd58436,17'd57304,17'd58562,17'd58563,17'd58564,17'd58565,17'd58566,17'd12838,17'd12696,17'd12839,17'd57168,17'd58567,17'd13501,17'd21980,17'd53465,17'd53468,17'd58568,17'd55417,17'd55699,17'd18685,17'd39661,17'd58312,17'd58446,17'd58447,17'd58447,17'd58448,17'd58446,17'd31597,17'd33243,17'd51118,17'd35644,17'd34380,17'd34381,17'd29645,17'd29645,17'd30220,17'd34381,17'd33882,17'd33243,17'd58314,17'd54732,17'd33882,17'd53250,17'd34833,17'd54732,17'd31773,17'd29646,17'd29481,17'd29336,17'd27857,17'd26758,17'd23855,17'd19407,17'd17348,17'd16321,17'd12419,17'd12857,17'd11957,17'd11962,17'd19158,17'd11521,17'd14673,17'd11524,17'd25812,17'd33083,17'd14675,17'd12265,17'd58569,17'd56734,17'd22479,17'd15442,17'd25152,17'd16691,17'd10028,17'd12867,17'd11404,17'd10027,17'd10175,17'd25814,17'd17123,17'd8724,17'd13257,17'd58570,17'd19648,17'd18454,17'd58571,17'd58572,17'd58573,17'd58574,17'd58575,17'd58576,17'd58577,17'd58578,17'd58579,17'd58580,17'd58581,17'd56857,17'd44696,17'd46545,17'd51313,17'd48908,17'd46664,17'd48526,17'd43288,17'd27372,17'd27258,17'd29535,17'd28724,17'd28481,17'd28594,17'd27882,17'd28485,17'd24898,17'd24416,17'd29100,17'd24249,17'd23731,17'd29688,17'd24745,17'd28974,17'd28485,17'd34283,17'd24745,17'd24897,17'd24898,17'd25030,17'd25030,17'd28254,17'd25178,17'd25029,17'd28254,17'd25178,17'd25180,17'd24745,17'd24416,17'd34467,17'd23732,17'd30579,17'd23389,17'd36426,17'd41273,17'd23389,17'd23217,17'd29530,17'd35430,17'd35430,17'd56973,17'd50464,17'd58582,17'd58583,17'd57564,17'd58584,17'd58585,17'd57702,17'd58586,17'd58587,17'd54205,17'd53846,17'd42742,17'd43978,17'd25435,17'd28597,17'd25567,17'd28130,17'd27765,17'd33000,17'd28597,17'd25567,17'd33000,17'd27765,17'd27765,17'd27765,17'd28597,17'd25709,17'd25709,17'd25567,17'd27765,17'd28594,17'd28594,17'd30456,17'd26402,17'd33970,17'd33970,17'd33009,17'd30456,17'd28600,17'd43022,17'd25178,17'd50364,17'd36009,17'd31660,17'd58588,17'd58589,17'd58590,17'd58591,17'd58592,17'd58593,17'd58594,17'd58595,17'd58596,17'd58597,17'd58598,17'd30467,17'd58599,17'd58600,17'd58601,17'd58602,17'd57584,17'd58603,17'd58604,17'd58605,17'd58606,17'd22922,17'd56087,17'd23268,17'd57588,17'd57589,17'd23973,17'd23107,17'd23798,17'd7493,17'd24478,17'd6381,17'd5144,17'd6067,17'd4997,17'd38442,17'd42910,17'd5327,17'd31552,17'd30180,17'd28185,17'd6554,17'd32073,17'd29740,17'd9933,17'd9091,17'd31891,17'd30333,17'd5335,17'd27697,17'd4526,17'd39938,17'd58607,17'd55745,17'd50672,17'd58608,17'd58609,17'd37293,17'd58234,17'd58610,17'd37159,17'd58611,17'd20704,17'd58612,17'd36446,17'd58613,17'd58234,17'd50380,17'd56205,17'd58614,17'd58120,17'd58362,17'd58615,17'd58616,17'd58617,17'd58618,17'd41154,17'd58491,17'd3046,17'd58619,17'd43461,17'd57355,17'd53738,17'd56207,17'd58620,17'd58125,17'd58241,17'd58126,17'd56321,17'd57604,17'd58621,17'd58622,17'd58002,17'd58623,17'd38578,17'd53745,17'd18385,17'd53151,17'd1121,17'd447,17'd429,17'd1540,17'd792,17'd636,17'd455,17'd637,17'd453,17'd1540,17'd17915,17'd607,17'd1667,17'd2097,17'd16256,17'd58624,17'd58496,17'd58625,17'd7705,17'd7705,17'd6258,17'd13933,17'd37957,17'd58626,17'd5627,17'd6237,17'd58498,17'd58627,17'd58628,17'd55166,17'd50496,17'd41157,17'd58629,17'd58499,17'd58500,17'd58501,17'd58630,17'd58631,17'd58377,17'd58378
},
'{
17'd2258,17'd2258,17'd2597,17'd2597,17'd2257,17'd1416,17'd3905,17'd18,17'd11,17'd11,17'd11,17'd11,17'd19,17'd18,17'd17,17'd1416,17'd2257,17'd2258,17'd3429,17'd52621,17'd10669,17'd3429,17'd3429,17'd57618,17'd57493,17'd1416,17'd468,17'd468,17'd29,17'd289,17'd290,17'd982,17'd12505,17'd6730,17'd15878,17'd473,17'd296,17'd661,17'd48,17'd57759,17'd56675,17'd56792,17'd57002,17'd57372,17'd1152,17'd1001,17'd58632,17'd1155,17'd58383,17'd58509,17'd58633,17'd21024,17'd58511,17'd58634,17'd21640,17'd58635,17'd58260,17'd58636,17'd58637,17'd58389,17'd56896,17'd58638,17'd58639,17'd58640,17'd13469,17'd7750,17'd7418,17'd9440,17'd9704,17'd58394,17'd58641,17'd58642,17'd58643,17'd58644,17'd8538,17'd7750,17'd7582,17'd8688,17'd58392,17'd58645,17'd58646,17'd58518,17'd58647,17'd58648,17'd48079,17'd47865,17'd47972,17'd48387,17'd53080,17'd48819,17'd57384,17'd54251,17'd58649,17'd58273,17'd56026,17'd58650,17'd56130,17'd58651,17'd55182,17'd58652,17'd58653,17'd58654,17'd58655,17'd58656,17'd58657,17'd58658,17'd58282,17'd58659,17'd58277,17'd58660,17'd58661,17'd58662,17'd58663,17'd58664,17'd58665,17'd58666,17'd3988,17'd58667,17'd58668,17'd58669,17'd58418,17'd55790,17'd58670,17'd58671,17'd54715,17'd53090,17'd41177,17'd58672,17'd58673,17'd58179,17'd58295,17'd58548,17'd58674,17'd58675,17'd58676,17'd58425,17'd58677,17'd58552,17'd58553,17'd58554,17'd58678,17'd58679,17'd58680,17'd13489,17'd58681,17'd58682,17'd58683,17'd58433,17'd58560,17'd58560,17'd58433,17'd58684,17'd58685,17'd58686,17'd58687,17'd58563,17'd58688,17'd58689,17'd58442,17'd58443,17'd12696,17'd58690,17'd12697,17'd58691,17'd12709,17'd23845,17'd58692,17'd56495,17'd45814,17'd56161,17'd55699,17'd28349,17'd58693,17'd58195,17'd58694,17'd58695,17'd58448,17'd58448,17'd32598,17'd32931,17'd36782,17'd51432,17'd34380,17'd34835,17'd37205,17'd29482,17'd30220,17'd34381,17'd33881,17'd33095,17'd56951,17'd31597,17'd33882,17'd33095,17'd54732,17'd57061,17'd36491,17'd36211,17'd29481,17'd28572,17'd28229,17'd24991,17'd20452,17'd14807,17'd16321,17'd16321,17'd12420,17'd12113,17'd11957,17'd19157,17'd13762,17'd11522,17'd14673,17'd10604,17'd10606,17'd15298,17'd11404,17'd12265,17'd58569,17'd10997,17'd10030,17'd14012,17'd22134,17'd17016,17'd8250,17'd8248,17'd17481,17'd8410,17'd10175,17'd15944,17'd17472,17'd8569,17'd32923,17'd58696,17'd18687,17'd11143,17'd15447,17'd58697,17'd58698,17'd58699,17'd58700,17'd58701,17'd58702,17'd58703,17'd58204,17'd58704,17'd58581,17'd56857,17'd58705,17'd58089,17'd41269,17'd47636,17'd49378,17'd41864,17'd33154,17'd34637,17'd28978,17'd27260,17'd28252,17'd27513,17'd28130,17'd27764,17'd27763,17'd24416,17'd28722,17'd23731,17'd31033,17'd23917,17'd29688,17'd32007,17'd25030,17'd24897,17'd24896,17'd24898,17'd25030,17'd25030,17'd25030,17'd25180,17'd27637,17'd25029,17'd27637,17'd25180,17'd25032,17'd24416,17'd34467,17'd24249,17'd24086,17'd23923,17'd22328,17'd23038,17'd22679,17'd23218,17'd23216,17'd30128,17'd38980,17'd50733,17'd50733,17'd56973,17'd52161,17'd58207,17'd58706,17'd58707,17'd58708,17'd58709,17'd58710,17'd58711,17'd56747,17'd53263,17'd50068,17'd43156,17'd32996,17'd31055,17'd28597,17'd27765,17'd28369,17'd27882,17'd25567,17'd25567,17'd28599,17'd27638,17'd28720,17'd27638,17'd25567,17'd25567,17'd27882,17'd27882,17'd44118,17'd39597,17'd30456,17'd58712,17'd33174,17'd33970,17'd26661,17'd26402,17'd33333,17'd26402,17'd25566,17'd39591,17'd30733,17'd35865,17'd42000,17'd50987,17'd42602,17'd58713,17'd58714,17'd58715,17'd58716,17'd58717,17'd58718,17'd58719,17'd58720,17'd58721,17'd58722,17'd58723,17'd58724,17'd58725,17'd58726,17'd56408,17'd58347,17'd58348,17'd20974,17'd58727,17'd29423,17'd58728,17'd57220,17'd30483,17'd57588,17'd57589,17'd23972,17'd24147,17'd10881,17'd58729,17'd4680,17'd24796,17'd6067,17'd5144,17'd4997,17'd38442,17'd42910,17'd4995,17'd5152,17'd5005,17'd5336,17'd31717,17'd7177,17'd9934,17'd9091,17'd37152,17'd33369,17'd5160,17'd5161,17'd4846,17'd49804,17'd55452,17'd55868,17'd49897,17'd38707,17'd38448,17'd37562,17'd58352,17'd58730,17'd58731,17'd36448,17'd3542,17'd3543,17'd58732,17'd58733,17'd3847,17'd57094,17'd58734,17'd55993,17'd58735,17'd57230,17'd58736,17'd42473,17'd58737,17'd39786,17'd44738,17'd58491,17'd58491,17'd58492,17'd58619,17'd58738,17'd58738,17'd58365,17'd58739,17'd58125,17'd56422,17'd58740,17'd58741,17'd56321,17'd54419,17'd58742,17'd55567,17'd58743,17'd58369,17'd58003,17'd58004,17'd3071,17'd960,17'd1545,17'd782,17'd609,17'd211,17'd1547,17'd248,17'd251,17'd462,17'd2420,17'd1093,17'd2778,17'd1962,17'd6407,17'd1946,17'd16256,17'd35060,17'd31899,17'd31899,17'd11061,17'd9414,17'd58744,17'd13933,17'd58745,17'd58497,17'd6238,17'd54780,17'd58746,17'd6405,17'd54514,17'd9245,17'd56665,17'd23299,17'd58747,17'd56991,17'd57358,17'd58501,17'd2359,17'd58748,17'd58749,17'd58750
},
'{
17'd2258,17'd2258,17'd2597,17'd2597,17'd1414,17'd1414,17'd17,17'd18,17'd11,17'd11,17'd11,17'd11,17'd19,17'd18,17'd17,17'd1416,17'd2257,17'd2258,17'd3429,17'd52621,17'd10802,17'd3593,17'd52621,17'd12195,17'd2426,17'd1414,17'd468,17'd468,17'd29,17'd289,17'd290,17'd3429,17'd3751,17'd6730,17'd15878,17'd58016,17'd986,17'd816,17'd57758,17'd58751,17'd58256,17'd56792,17'd56892,17'd56892,17'd1292,17'd1152,17'd493,17'd58752,17'd58383,17'd58509,17'd58633,17'd1565,17'd1849,17'd1990,17'd58753,17'd2961,17'd3769,17'd4445,17'd57497,17'd58754,17'd58755,17'd58756,17'd58757,17'd58758,17'd23501,17'd8537,17'd46366,17'd9440,17'd9704,17'd58394,17'd58759,17'd58760,17'd58761,17'd51948,17'd8066,17'd4611,17'd4767,17'd8688,17'd58762,17'd58763,17'd58764,17'd58765,17'd58647,17'd57382,17'd58030,17'd47971,17'd48299,17'd47971,17'd53080,17'd56125,17'd58766,17'd57635,17'd58400,17'd55185,17'd55674,17'd55182,17'd58767,17'd58768,17'd57921,17'd58408,17'd57396,17'd57779,17'd58769,17'd58279,17'd58770,17'd58771,17'd57132,17'd58772,17'd1459,17'd57022,17'd57778,17'd58773,17'd58774,17'd57520,17'd58775,17'd58666,17'd58776,17'd58777,17'd58778,17'd58779,17'd58052,17'd58780,17'd58781,17'd58782,17'd58783,17'd58784,17'd54908,17'd58785,17'd56929,17'd58786,17'd57798,17'd58548,17'd58674,17'd58548,17'd58787,17'd58425,17'd58788,17'd58789,17'd58790,17'd58791,17'd58678,17'd58792,17'd58793,17'd58794,17'd58795,17'd58796,17'd58797,17'd58433,17'd58560,17'd58560,17'd58798,17'd58434,17'd58433,17'd58799,17'd58800,17'd58801,17'd58802,17'd58565,17'd58566,17'd58566,17'd58566,17'd57427,17'd58803,17'd58804,17'd14512,17'd23676,17'd57312,17'd58805,17'd55316,17'd55612,17'd55699,17'd28349,17'd58806,17'd58195,17'd58694,17'd58695,17'd58448,17'd32600,17'd32598,17'd32931,17'd34047,17'd34047,17'd33574,17'd34381,17'd29481,17'd29482,17'd30220,17'd34835,17'd33881,17'd56619,17'd56951,17'd31597,17'd33096,17'd56619,17'd54732,17'd57061,17'd30220,17'd30373,17'd36347,17'd28572,17'd28229,17'd24991,17'd20452,17'd12108,17'd17348,17'd16321,17'd12420,17'd12113,17'd11957,17'd15810,17'd13762,17'd16068,17'd14810,17'd13886,17'd11528,17'd16065,17'd15429,17'd12265,17'd17852,17'd54118,17'd13529,17'd13770,17'd19036,17'd22133,17'd13648,17'd8579,17'd21987,17'd8410,17'd9042,17'd10174,17'd17472,17'd8724,17'd58807,17'd58696,17'd58808,17'd58809,17'd58810,17'd58811,17'd58812,17'd58813,17'd58814,17'd58815,17'd58816,17'd58817,17'd58325,17'd58818,17'd58458,17'd45982,17'd58819,17'd58820,17'd51076,17'd48523,17'd49679,17'd42599,17'd32343,17'd30586,17'd29535,17'd42147,17'd38538,17'd28598,17'd25317,17'd28596,17'd29240,17'd23916,17'd30275,17'd23920,17'd24086,17'd23731,17'd23916,17'd28851,17'd24745,17'd24897,17'd24898,17'd24897,17'd24897,17'd24897,17'd24897,17'd24897,17'd24897,17'd24898,17'd25180,17'd24895,17'd24416,17'd24249,17'd24086,17'd23733,17'd29827,17'd23216,17'd22678,17'd22332,17'd32827,17'd23217,17'd29828,17'd23567,17'd58821,17'd56751,17'd58822,17'd50730,17'd51307,17'd58823,17'd51232,17'd58824,17'd58825,17'd58709,17'd58826,17'd52076,17'd58827,17'd50361,17'd43017,17'd43978,17'd28594,17'd31055,17'd28597,17'd27765,17'd28369,17'd27882,17'd25567,17'd25567,17'd28599,17'd28594,17'd28594,17'd27638,17'd25567,17'd28597,17'd27882,17'd27882,17'd25951,17'd39597,17'd30456,17'd30456,17'd33970,17'd32364,17'd26661,17'd26402,17'd26402,17'd33510,17'd33510,17'd32353,17'd33801,17'd36288,17'd46949,17'd21695,17'd58828,17'd58829,17'd58830,17'd58831,17'd58832,17'd58833,17'd58834,17'd58835,17'd44719,17'd24750,17'd58836,17'd58837,17'd58838,17'd58839,17'd58840,17'd58841,17'd57086,17'd58842,17'd58479,17'd58843,17'd58844,17'd22062,17'd57220,17'd23620,17'd56875,17'd57589,17'd55986,17'd24307,17'd7493,17'd7659,17'd5322,17'd5322,17'd6067,17'd4997,17'd4997,17'd5144,17'd42910,17'd5152,17'd31716,17'd5004,17'd27935,17'd6554,17'd7177,17'd10238,17'd32073,17'd31891,17'd30333,17'd5160,17'd34921,17'd50081,17'd55351,17'd58845,17'd57347,17'd38707,17'd58846,17'd58847,17'd58848,17'd58849,17'd58850,17'd58851,17'd36448,17'd36448,17'd3543,17'd58852,17'd58853,17'd49298,17'd58854,17'd58610,17'd56987,17'd58855,17'd45064,17'd3046,17'd22602,17'd58856,17'd58857,17'd44963,17'd58491,17'd3046,17'd44016,17'd42919,17'd58858,17'd57231,17'd55996,17'd55996,17'd56422,17'd53739,17'd58859,17'd53668,17'd55267,17'd54511,17'd58860,17'd58861,17'd58862,17'd38714,17'd53593,17'd54688,17'd3222,17'd960,17'd52103,17'd232,17'd233,17'd39949,17'd1547,17'd19102,17'd591,17'd182,17'd211,17'd17915,17'd1539,17'd1380,17'd2905,17'd3073,17'd35060,17'd58863,17'd28066,17'd33051,17'd58864,17'd58865,17'd14858,17'd37709,17'd58866,17'd58867,17'd6238,17'd58868,17'd58869,17'd5774,17'd58870,17'd9245,17'd58871,17'd40560,17'd52532,17'd36042,17'd53362,17'd58872,17'd58873,17'd58874,17'd58377,17'd58750
},
'{
17'd2258,17'd2258,17'd2597,17'd2597,17'd1414,17'd1414,17'd17,17'd18,17'd11,17'd10,17'd10,17'd11,17'd19,17'd18,17'd17,17'd17,17'd2257,17'd2425,17'd2258,17'd52621,17'd10802,17'd10669,17'd10669,17'd58503,17'd12194,17'd2257,17'd1416,17'd1416,17'd29,17'd289,17'd290,17'd982,17'd12505,17'd4086,17'd16011,17'd16392,17'd473,17'd1131,17'd819,17'd58255,17'd58256,17'd56674,17'd56892,17'd56892,17'd1430,17'd1292,17'd1001,17'd1431,17'd58019,17'd58509,17'd1298,17'd58875,17'd58876,17'd57114,17'd57256,17'd2278,17'd29901,17'd58877,17'd58878,17'd58637,17'd58879,17'd3934,17'd58880,17'd58881,17'd57500,17'd9300,17'd13471,17'd13471,17'd13845,17'd48301,17'd58762,17'd58760,17'd3787,17'd52203,17'd8068,17'd8539,17'd8688,17'd4464,17'd58882,17'd58642,17'd3634,17'd58883,17'd58270,17'd54350,17'd57120,17'd52710,17'd47973,17'd47865,17'd52850,17'd53080,17'd49199,17'd48820,17'd55774,17'd55900,17'd56241,17'd58159,17'd58884,17'd58767,17'd58885,17'd58886,17'd57648,17'd57779,17'd58887,17'd58888,17'd58889,17'd58890,17'd58891,17'd58892,17'd57275,17'd58893,17'd56583,17'd58894,17'd58895,17'd58285,17'd58896,17'd58897,17'd58898,17'd58899,17'd58900,17'd58901,17'd58902,17'd58419,17'd58903,17'd56362,17'd58904,17'd58905,17'd54908,17'd58906,17'd58907,17'd57037,17'd57292,17'd58908,17'd58674,17'd58548,17'd58909,17'd58910,17'd58911,17'd58912,17'd58790,17'd58791,17'd58913,17'd58914,17'd58915,17'd58916,17'd58917,17'd58918,17'd58919,17'd58797,17'd58433,17'd58434,17'd58920,17'd58921,17'd58922,17'd58923,17'd58924,17'd58925,17'd58926,17'd58927,17'd13116,17'd58928,17'd58189,17'd12977,17'd12696,17'd58929,17'd58567,17'd13129,17'd21201,17'd58930,17'd58931,17'd38503,17'd55699,17'd39825,17'd58806,17'd58932,17'd58933,17'd58934,17'd58933,17'd32443,17'd32441,17'd32927,17'd33730,17'd33882,17'd33574,17'd36937,17'd29481,17'd29482,17'd29785,17'd31289,17'd33730,17'd58935,17'd57181,17'd37985,17'd34385,17'd36214,17'd31597,17'd30371,17'd30220,17'd30373,17'd28571,17'd27857,17'd27737,17'd23511,17'd20452,17'd12579,17'd12580,17'd16321,17'd12420,17'd12113,17'd11963,17'd15810,17'd13762,17'd16068,17'd13138,17'd10477,17'd15688,17'd18080,17'd15429,17'd54046,17'd14266,17'd58936,17'd58937,17'd7793,17'd18921,17'd16919,17'd53836,17'd8418,17'd8413,17'd8410,17'd9042,17'd17480,17'd17123,17'd8569,17'd58807,17'd58696,17'd58938,17'd58809,17'd58939,17'd58940,17'd58941,17'd58942,17'd58943,17'd58944,17'd58945,17'd58946,17'd50358,17'd47434,17'd58458,17'd58947,17'd58948,17'd54573,17'd47044,17'd46662,17'd46102,17'd44478,17'd27372,17'd27027,17'd42147,17'd33156,17'd28253,17'd25567,17'd27511,17'd34283,17'd29100,17'd24087,17'd29099,17'd30127,17'd23920,17'd24086,17'd23917,17'd24252,17'd28718,17'd24417,17'd25030,17'd24897,17'd24897,17'd24898,17'd24898,17'd24897,17'd24897,17'd25032,17'd32007,17'd24416,17'd24249,17'd31033,17'd31502,17'd30579,17'd23215,17'd32830,17'd23573,17'd30276,17'd23389,17'd23217,17'd23388,17'd38980,17'd58949,17'd58950,17'd58707,17'd58706,17'd50730,17'd57455,17'd40680,17'd58951,17'd57833,17'd58952,17'd50734,17'd56746,17'd58953,17'd50154,17'd43425,17'd29970,17'd31366,17'd32669,17'd25567,17'd27765,17'd25567,17'd28597,17'd25567,17'd25567,17'd28598,17'd28594,17'd28594,17'd28594,17'd25567,17'd27882,17'd34127,17'd30903,17'd33814,17'd25951,17'd30456,17'd26402,17'd32364,17'd32364,17'd26402,17'd26402,17'd58954,17'd26531,17'd32689,17'd37512,17'd37511,17'd45875,17'd21848,17'd52073,17'd58955,17'd51835,17'd58715,17'd58956,17'd58957,17'd58958,17'd58959,17'd58960,17'd58961,17'd58962,17'd58963,17'd58964,17'd53212,17'd58965,17'd58966,17'd56764,17'd57585,17'd20513,17'd58967,17'd58968,17'd58969,17'd58970,17'd57727,17'd23622,17'd23623,17'd23105,17'd23452,17'd23457,17'd24308,17'd24477,17'd5322,17'd5322,17'd5145,17'd38058,17'd33992,17'd4999,17'd5155,17'd34791,17'd28418,17'd25627,17'd27935,17'd6390,17'd7499,17'd9091,17'd31717,17'd33369,17'd25627,17'd5329,17'd5157,17'd58971,17'd56415,17'd58972,17'd58973,17'd58846,17'd58847,17'd58974,17'd58975,17'd58976,17'd50285,17'd3542,17'd36448,17'd36448,17'd58851,17'd58977,17'd58978,17'd49192,17'd58357,17'd58355,17'd57480,17'd58979,17'd44962,17'd41900,17'd58980,17'd44017,17'd58981,17'd58982,17'd58491,17'd58492,17'd42919,17'd58983,17'd58984,17'd58985,17'd58739,17'd55996,17'd56774,17'd58986,17'd58741,17'd53668,17'd56322,17'd2208,17'd58987,17'd58988,17'd58989,17'd927,17'd2419,17'd450,17'd960,17'd52103,17'd1114,17'd607,17'd2778,17'd211,17'd1547,17'd247,17'd50187,17'd965,17'd2255,17'd1097,17'd260,17'd1667,17'd412,17'd2098,17'd5030,17'd28066,17'd28066,17'd27949,17'd58990,17'd9414,17'd6891,17'd58991,17'd58992,17'd53293,17'd58993,17'd58994,17'd58994,17'd3568,17'd58870,17'd2389,17'd19360,17'd22098,17'd58995,17'd58996,17'd58997,17'd58998,17'd58999,17'd1926,17'd58631,17'd59000
},
'{
17'd2258,17'd2258,17'd2597,17'd2597,17'd1414,17'd1414,17'd16,17'd16,17'd19,17'd10,17'd10,17'd10,17'd19,17'd18,17'd16,17'd17,17'd1414,17'd2257,17'd2258,17'd3429,17'd10802,17'd10669,17'd10669,17'd54978,17'd12195,17'd2597,17'd1414,17'd1416,17'd29,17'd289,17'd290,17'd469,17'd12505,17'd4086,17'd16011,17'd16392,17'd659,17'd15497,17'd298,17'd58255,17'd58256,17'd59001,17'd56791,17'd56892,17'd57003,17'd1430,17'd1152,17'd494,17'd58507,17'd1157,17'd1297,17'd1434,17'd58876,17'd16968,17'd59002,17'd59003,17'd59004,17'd59005,17'd57258,17'd57497,17'd59006,17'd59007,17'd3455,17'd59008,17'd57908,17'd16170,17'd59009,17'd13846,17'd7582,17'd8371,17'd58762,17'd58760,17'd59010,17'd3787,17'd52111,17'd3954,17'd4291,17'd59011,17'd58393,17'd58760,17'd3634,17'd53449,17'd58270,17'd58518,17'd53370,17'd57012,17'd52710,17'd59012,17'd56572,17'd53232,17'd55483,17'd57504,17'd54251,17'd56804,17'd55184,17'd59013,17'd59014,17'd59015,17'd59016,17'd59017,17'd58654,17'd59018,17'd57918,17'd59019,17'd59020,17'd59021,17'd57022,17'd59022,17'd59023,17'd59024,17'd58887,17'd59025,17'd59026,17'd56812,17'd58896,17'd59027,17'd57025,17'd2322,17'd59028,17'd59029,17'd59030,17'd59031,17'd59032,17'd56037,17'd59033,17'd59034,17'd59035,17'd59036,17'd59037,17'd56929,17'd57150,17'd59038,17'd59039,17'd58674,17'd59040,17'd59041,17'd59041,17'd58787,17'd59042,17'd59043,17'd59044,17'd59045,17'd59046,17'd58915,17'd59047,17'd59048,17'd59049,17'd59050,17'd58434,17'd59051,17'd58921,17'd59052,17'd59053,17'd59054,17'd59055,17'd59056,17'd59057,17'd58562,17'd59058,17'd59059,17'd59060,17'd59059,17'd59061,17'd12554,17'd59062,17'd19151,17'd54192,17'd56493,17'd59063,17'd55416,17'd56497,17'd39825,17'd59064,17'd32129,17'd59065,17'd59066,17'd58933,17'd59067,17'd32441,17'd35236,17'd33096,17'd33096,17'd33409,17'd36491,17'd29481,17'd29482,17'd29785,17'd31289,17'd33096,17'd58314,17'd59068,17'd37985,17'd36214,17'd31597,17'd30371,17'd29647,17'd29482,17'd28944,17'd28818,17'd27857,17'd26629,17'd23855,17'd12108,17'd12579,17'd12580,17'd16321,17'd12420,17'd11806,17'd12861,17'd11395,17'd11522,17'd16068,17'd13138,17'd10477,17'd25675,17'd18080,17'd15429,17'd22133,17'd24552,17'd59069,17'd59070,17'd59071,17'd15442,17'd55523,17'd23519,17'd10028,17'd25147,17'd8412,17'd10176,17'd17480,17'd17472,17'd9046,17'd32923,17'd8889,17'd58938,17'd10864,17'd59072,17'd59073,17'd59074,17'd59075,17'd59076,17'd59077,17'd59078,17'd59079,17'd49781,17'd47434,17'd59080,17'd59081,17'd59082,17'd48261,17'd50067,17'd57713,17'd52678,17'd47927,17'd30586,17'd26782,17'd43838,17'd44230,17'd44229,17'd28369,17'd29244,17'd23561,17'd28722,17'd23733,17'd23387,17'd23736,17'd30127,17'd31033,17'd30431,17'd34467,17'd24743,17'd23561,17'd24745,17'd24896,17'd24896,17'd24895,17'd25032,17'd24895,17'd24895,17'd30126,17'd28851,17'd24415,17'd24086,17'd30127,17'd30579,17'd32351,17'd41273,17'd41419,17'd23573,17'd22330,17'd30277,17'd32191,17'd23736,17'd40680,17'd56751,17'd58950,17'd59083,17'd59083,17'd53192,17'd51160,17'd58949,17'd58583,17'd59084,17'd59085,17'd59086,17'd50562,17'd53487,17'd53486,17'd43977,17'd28717,17'd31856,17'd31055,17'd27765,17'd25567,17'd25567,17'd28597,17'd25567,17'd27765,17'd27638,17'd28720,17'd28594,17'd28594,17'd25567,17'd27882,17'd34127,17'd30903,17'd33814,17'd33814,17'd39597,17'd26661,17'd26287,17'd32364,17'd26661,17'd59087,17'd59088,17'd59089,17'd59090,17'd59091,17'd22680,17'd22164,17'd47746,17'd59092,17'd59093,17'd59094,17'd59095,17'd59096,17'd24428,17'd59097,17'd59098,17'd59099,17'd59100,17'd59101,17'd48719,17'd59102,17'd59103,17'd59104,17'd56408,17'd59105,17'd59106,17'd59107,17'd59108,17'd59109,17'd29882,17'd57220,17'd23622,17'd23624,17'd23624,17'd23105,17'd56088,17'd8911,17'd24478,17'd24476,17'd5322,17'd6381,17'd38442,17'd59110,17'd33992,17'd4999,17'd41459,17'd34791,17'd5005,17'd30638,17'd31717,17'd6219,17'd7499,17'd6554,17'd33369,17'd31553,17'd5329,17'd27697,17'd50081,17'd54862,17'd52272,17'd59111,17'd56877,17'd58847,17'd58974,17'd58975,17'd58849,17'd59112,17'd58851,17'd59113,17'd36448,17'd36893,17'd58851,17'd36590,17'd58978,17'd58850,17'd50285,17'd59114,17'd59115,17'd58122,17'd41309,17'd59116,17'd59117,17'd46789,17'd59118,17'd58982,17'd59119,17'd44266,17'd42919,17'd58738,17'd57356,17'd59120,17'd58739,17'd56421,17'd58986,17'd58986,17'd58741,17'd53668,17'd56322,17'd58621,17'd59121,17'd35205,17'd59122,17'd59123,17'd800,17'd1681,17'd52021,17'd52021,17'd427,17'd954,17'd1539,17'd408,17'd39949,17'd59124,17'd49713,17'd2255,17'd408,17'd41316,17'd1666,17'd5957,17'd14178,17'd5631,17'd28066,17'd27949,17'd31562,17'd37168,17'd59125,17'd10395,17'd13933,17'd5938,17'd58626,17'd57103,17'd59126,17'd5774,17'd59127,17'd59128,17'd59129,17'd58372,17'd58009,17'd58010,17'd58499,17'd57358,17'd59130,17'd35057,17'd2070,17'd59131,17'd58631,17'd59132
},
'{
17'd2258,17'd2258,17'd2597,17'd2597,17'd1414,17'd1414,17'd17,17'd18,17'd11,17'd10,17'd10,17'd10,17'd19,17'd18,17'd16,17'd16,17'd1416,17'd2257,17'd2597,17'd3429,17'd3101,17'd2593,17'd2935,17'd14188,17'd57618,17'd2258,17'd2257,17'd2257,17'd289,17'd289,17'd30,17'd1129,17'd10924,17'd16392,17'd59133,17'd57896,17'd659,17'd15362,17'd58505,17'd48,17'd58256,17'd59001,17'd56791,17'd56892,17'd57003,17'd57003,17'd1292,17'd1001,17'd1154,17'd1156,17'd1157,17'd59134,17'd20409,17'd1987,17'd55893,17'd2131,17'd58387,17'd16393,17'd59135,17'd57497,17'd59136,17'd59137,17'd58262,17'd58515,17'd59138,17'd59139,17'd16882,17'd13846,17'd5410,17'd8066,17'd59140,17'd58759,17'd57769,17'd57769,17'd3787,17'd4770,17'd4125,17'd4291,17'd58393,17'd58517,17'd3634,17'd3478,17'd59141,17'd58270,17'd53232,17'd56686,17'd59142,17'd59142,17'd57910,17'd59143,17'd55483,17'd57504,17'd54251,17'd58150,17'd54803,17'd56029,17'd57647,17'd56024,17'd58278,17'd59144,17'd57518,17'd57918,17'd59018,17'd59145,17'd58527,17'd59146,17'd59147,17'd59148,17'd59149,17'd56810,17'd57391,17'd59150,17'd59151,17'd59152,17'd1037,17'd58896,17'd59153,17'd2501,17'd2855,17'd59154,17'd59155,17'd59156,17'd59157,17'd5283,17'd59158,17'd59159,17'd59160,17'd59161,17'd59162,17'd56045,17'd57153,17'd59163,17'd58675,17'd58674,17'd59164,17'd59165,17'd59166,17'd59167,17'd59042,17'd59168,17'd59169,17'd59045,17'd59170,17'd59171,17'd58793,17'd59172,17'd59173,17'd59174,17'd58922,17'd59175,17'd59176,17'd59177,17'd59178,17'd59179,17'd59180,17'd59055,17'd58924,17'd58800,17'd59057,17'd59181,17'd59182,17'd59183,17'd59060,17'd12553,17'd59184,17'd59185,17'd14920,17'd21049,17'd59186,17'd55123,17'd38367,17'd39661,17'd30978,17'd30977,17'd59187,17'd59067,17'd59188,17'd59187,17'd59189,17'd58448,17'd33093,17'd33093,17'd33727,17'd29646,17'd30373,17'd29482,17'd30073,17'd31289,17'd31591,17'd58314,17'd57439,17'd30678,17'd37985,17'd30371,17'd29785,17'd30220,17'd29482,17'd36347,17'd28460,17'd28104,17'd27121,17'd12255,17'd23168,17'd16203,17'd14130,17'd11960,17'd11961,17'd12861,17'd18805,17'd11520,17'd11522,17'd11523,17'd10605,17'd22296,17'd25675,17'd34382,17'd31759,17'd11279,17'd24369,17'd59190,17'd59191,17'd59192,17'd14391,17'd55124,17'd23519,17'd8580,17'd25147,17'd8412,17'd16440,17'd17848,17'd17472,17'd9046,17'd32923,17'd8889,17'd24046,17'd59193,17'd58939,17'd59194,17'd59195,17'd59196,17'd59197,17'd59198,17'd59199,17'd59200,17'd59201,17'd59202,17'd59203,17'd59204,17'd56748,17'd51646,17'd47237,17'd50070,17'd51746,17'd47927,17'd30586,17'd28853,17'd46753,17'd43155,17'd43836,17'd28850,17'd25179,17'd34884,17'd23918,17'd29530,17'd32191,17'd29829,17'd29376,17'd23920,17'd29534,17'd32659,17'd24742,17'd24252,17'd24252,17'd24742,17'd24742,17'd24252,17'd24742,17'd35159,17'd32659,17'd30431,17'd23731,17'd23564,17'd29376,17'd29530,17'd23217,17'd39131,17'd34458,17'd34458,17'd22678,17'd22329,17'd30277,17'd23569,17'd31341,17'd40680,17'd58821,17'd52815,17'd59205,17'd52668,17'd46427,17'd39133,17'd59206,17'd58461,17'd59207,17'd59208,17'd59209,17'd52967,17'd53486,17'd43291,17'd27511,17'd28480,17'd31366,17'd28597,17'd27765,17'd25567,17'd25567,17'd25567,17'd28598,17'd27638,17'd28720,17'd28720,17'd28594,17'd27765,17'd28369,17'd27882,17'd34127,17'd38812,17'd32689,17'd33814,17'd33510,17'd26402,17'd59210,17'd59210,17'd59211,17'd32848,17'd59212,17'd59213,17'd59214,17'd31350,17'd22159,17'd22011,17'd51633,17'd47836,17'd47149,17'd58469,17'd59215,17'd59216,17'd59217,17'd59218,17'd59219,17'd26179,17'd59220,17'd59221,17'd59222,17'd59223,17'd59224,17'd59225,17'd56651,17'd59226,17'd58348,17'd20973,17'd59227,17'd22056,17'd29588,17'd57220,17'd23622,17'd23105,17'd57589,17'd23973,17'd55863,17'd7493,17'd24478,17'd24476,17'd4837,17'd5145,17'd4997,17'd59110,17'd33992,17'd4999,17'd41459,17'd34791,17'd4848,17'd37030,17'd31717,17'd9091,17'd6219,17'd31717,17'd31553,17'd30637,17'd5161,17'd34921,17'd49896,17'd59228,17'd59111,17'd59229,17'd59230,17'd58974,17'd59231,17'd4033,17'd36738,17'd49192,17'd59232,17'd59233,17'd36448,17'd36893,17'd58731,17'd59234,17'd58978,17'd58852,17'd59235,17'd36742,17'd45652,17'd59236,17'd59237,17'd59238,17'd46990,17'd46990,17'd52837,17'd45065,17'd41309,17'd44016,17'd43189,17'd57231,17'd59239,17'd59240,17'd56421,17'd59239,17'd58986,17'd59241,17'd53668,17'd53668,17'd56002,17'd59242,17'd59243,17'd59244,17'd24953,17'd31099,17'd593,17'd210,17'd57888,17'd59245,17'd953,17'd642,17'd935,17'd2778,17'd40412,17'd39949,17'd2255,17'd262,17'd41005,17'd426,17'd1823,17'd2905,17'd2098,17'd5777,17'd32082,17'd28315,17'd31729,17'd27949,17'd12923,17'd8187,17'd4883,17'd51761,17'd56549,17'd38718,17'd58993,17'd3568,17'd59128,17'd59128,17'd59246,17'd58245,17'd2388,17'd58010,17'd59247,17'd57358,17'd59130,17'd59248,17'd2070,17'd59249,17'd58631,17'd57617
},
'{
17'd2258,17'd2258,17'd2597,17'd2597,17'd2257,17'd1414,17'd17,17'd16,17'd19,17'd10,17'd10,17'd10,17'd19,17'd18,17'd16,17'd16,17'd1416,17'd2257,17'd2596,17'd3429,17'd2935,17'd2593,17'd2935,17'd3251,17'd58503,17'd2426,17'd2425,17'd2257,17'd289,17'd289,17'd30,17'd469,17'd12505,17'd16392,17'd59133,17'd59133,17'd472,17'd15362,17'd477,17'd59250,17'd59251,17'd59001,17'd56672,17'd56791,17'd57003,17'd57003,17'd1292,17'd1001,17'd1294,17'd1155,17'd58509,17'd1298,17'd18518,17'd59252,17'd56335,17'd59253,17'd59254,17'd59255,17'd59256,17'd59257,17'd59258,17'd58879,17'd59259,17'd59260,17'd59261,17'd59262,17'd16522,17'd59263,17'd5090,17'd4611,17'd58644,17'd58759,17'd58395,17'd54095,17'd3634,17'd59264,17'd4290,17'd59265,17'd58393,17'd58517,17'd3634,17'd3478,17'd59266,17'd59267,17'd59143,17'd53370,17'd56686,17'd59268,17'd54173,17'd59269,17'd53685,17'd57504,17'd59270,17'd59271,17'd56020,17'd55907,17'd57646,17'd58524,17'd57917,17'd59272,17'd59273,17'd59274,17'd59275,17'd57918,17'd59276,17'd59277,17'd59278,17'd59279,17'd59149,17'd59280,17'd59281,17'd59282,17'd59283,17'd57023,17'd59284,17'd59285,17'd59286,17'd59287,17'd59288,17'd59289,17'd59290,17'd59291,17'd59292,17'd59293,17'd59294,17'd59295,17'd58544,17'd53172,17'd54445,17'd55798,17'd56824,17'd58176,17'd58908,17'd58549,17'd59296,17'd59297,17'd59298,17'd59165,17'd59042,17'd59168,17'd59299,17'd59300,17'd59301,17'd59170,17'd59302,17'd59303,17'd59304,17'd59305,17'd59306,17'd59176,17'd59307,17'd59177,17'd59308,17'd59309,17'd59310,17'd59311,17'd59312,17'd59313,17'd59314,17'd59315,17'd59316,17'd59317,17'd59318,17'd13492,17'd13117,17'd57308,17'd14799,17'd20444,17'd59319,17'd58931,17'd57953,17'd39661,17'd31772,17'd57817,17'd59320,17'd32288,17'd32289,17'd32288,17'd30680,17'd58196,17'd32933,17'd34385,17'd34698,17'd29646,17'd30373,17'd29482,17'd30073,17'd34835,17'd56619,17'd58314,17'd57554,17'd30678,17'd37985,17'd30371,17'd30220,17'd29482,17'd28944,17'd50213,17'd28460,17'd26629,17'd24991,17'd12255,17'd23168,17'd16203,17'd14130,17'd11960,17'd11961,17'd12861,17'd13885,17'd16069,17'd23337,17'd25280,17'd10476,17'd10606,17'd17839,17'd18080,17'd31759,17'd59321,17'd59322,17'd54929,17'd59323,17'd59324,17'd53549,17'd59325,17'd11533,17'd10028,17'd21987,17'd26260,17'd26633,17'd26498,17'd23859,17'd8569,17'd32923,17'd58696,17'd59326,17'd59193,17'd58939,17'd59327,17'd59328,17'd59329,17'd59330,17'd59331,17'd59199,17'd59332,17'd59333,17'd48251,17'd59334,17'd59335,17'd48353,17'd52822,17'd47238,17'd50070,17'd51746,17'd43838,17'd27027,17'd27258,17'd43548,17'd53262,17'd38156,17'd41730,17'd29976,17'd28852,17'd23565,17'd32191,17'd23217,17'd23215,17'd29686,17'd23565,17'd24249,17'd35159,17'd28851,17'd30126,17'd24416,17'd24416,17'd24252,17'd29100,17'd24090,17'd24249,17'd24249,17'd31033,17'd30275,17'd29242,17'd23387,17'd32191,17'd36426,17'd22859,17'd23573,17'd22332,17'd32827,17'd23389,17'd23215,17'd37511,17'd38980,17'd34112,17'd56751,17'd58824,17'd59206,17'd59336,17'd46550,17'd59337,17'd59338,17'd50645,17'd58460,17'd59339,17'd48895,17'd43291,17'd43157,17'd39443,17'd27512,17'd27512,17'd27882,17'd25567,17'd27765,17'd25567,17'd25567,17'd27765,17'd27638,17'd28594,17'd28720,17'd28720,17'd28594,17'd25567,17'd27882,17'd27511,17'd33345,17'd38812,17'd32689,17'd40379,17'd59340,17'd26402,17'd31845,17'd59211,17'd32848,17'd59341,17'd59342,17'd59343,17'd59344,17'd45379,17'd21847,17'd56755,17'd59345,17'd51238,17'd59346,17'd59347,17'd58717,17'd59348,17'd59349,17'd59350,17'd59351,17'd59352,17'd59353,17'd59354,17'd59355,17'd59356,17'd59357,17'd59358,17'd58228,17'd28051,17'd59359,17'd20974,17'd59360,17'd21898,17'd58231,17'd57346,17'd56875,17'd23105,17'd57589,17'd23452,17'd23974,17'd7658,17'd24477,17'd5322,17'd5145,17'd38442,17'd38058,17'd38058,17'd33992,17'd33841,17'd41459,17'd4684,17'd5162,17'd36887,17'd31717,17'd36586,17'd6554,17'd30638,17'd5004,17'd5005,17'd5157,17'd50586,17'd4370,17'd59361,17'd59362,17'd59363,17'd59230,17'd59364,17'd4033,17'd59365,17'd58613,17'd58850,17'd59232,17'd59235,17'd36448,17'd37159,17'd59366,17'd59367,17'd36446,17'd58977,17'd36449,17'd51576,17'd53285,17'd43737,17'd59237,17'd53285,17'd35056,17'd59368,17'd59369,17'd59370,17'd59371,17'd42919,17'd58738,17'd57356,17'd56421,17'd56421,17'd59239,17'd59239,17'd53739,17'd59241,17'd53668,17'd55358,17'd2070,17'd32247,17'd59372,17'd1662,17'd1086,17'd432,17'd244,17'd7681,17'd57888,17'd1544,17'd953,17'd970,17'd641,17'd646,17'd408,17'd59373,17'd802,17'd261,17'd3899,17'd1666,17'd5957,17'd1946,17'd5631,17'd33050,17'd27707,17'd28315,17'd31101,17'd36905,17'd38460,17'd6094,17'd58991,17'd38717,17'd38718,17'd54163,17'd39326,17'd59128,17'd5354,17'd59128,17'd59374,17'd59375,17'd19237,17'd22262,17'd59376,17'd53362,17'd59377,17'd59378,17'd57604,17'd59379,17'd58376,17'd57617
},
'{
17'd2258,17'd2258,17'd2597,17'd2597,17'd2257,17'd1414,17'd17,17'd18,17'd11,17'd10,17'd808,17'd10,17'd19,17'd18,17'd16,17'd16,17'd1416,17'd1414,17'd2596,17'd3752,17'd2935,17'd2593,17'd2593,17'd3251,17'd59380,17'd12194,17'd2425,17'd2257,17'd289,17'd289,17'd30,17'd1129,17'd11071,17'd12504,17'd59133,17'd59133,17'd472,17'd59381,17'd987,17'd46,17'd59382,17'd59001,17'd56672,17'd56791,17'd57003,17'd57003,17'd57006,17'd1293,17'd1002,17'd59383,17'd58509,17'd1298,17'd21024,17'd59384,17'd2127,17'd32733,17'd34170,17'd59385,17'd59386,17'd57117,17'd57378,17'd59006,17'd59387,17'd59388,17'd59389,17'd4455,17'd22461,17'd6134,17'd5410,17'd4767,17'd48301,17'd58759,17'd53018,17'd53448,17'd3789,17'd3476,17'd59390,17'd4123,17'd58393,17'd58882,17'd59391,17'd3477,17'd3790,17'd59267,17'd54350,17'd53607,17'd53607,17'd59143,17'd53523,17'd59269,17'd53685,17'd57504,17'd59392,17'd59271,17'd56021,17'd56351,17'd56132,17'd59393,17'd59394,17'd59395,17'd56914,17'd57391,17'd59396,17'd58771,17'd59397,17'd59398,17'd56584,17'd59399,17'd59400,17'd58651,17'd58893,17'd59401,17'd56355,17'd58662,17'd59402,17'd59403,17'd59404,17'd59405,17'd59406,17'd59407,17'd59408,17'd59409,17'd59410,17'd59411,17'd59294,17'd59412,17'd59413,17'd53695,17'd59414,17'd59415,17'd56045,17'd59416,17'd58059,17'd59417,17'd59418,17'd59418,17'd59418,17'd59165,17'd59042,17'd59168,17'd59299,17'd59300,17'd59419,17'd59420,17'd59421,17'd59422,17'd59423,17'd59304,17'd59309,17'd59424,17'd59425,17'd59425,17'd59426,17'd59427,17'd59428,17'd59429,17'd59180,17'd59430,17'd59431,17'd59432,17'd59433,17'd59315,17'd59434,17'd59183,17'd12977,17'd11781,17'd58567,17'd55312,17'd54922,17'd59435,17'd59436,17'd56947,17'd56616,17'd56844,17'd30977,17'd58077,17'd59320,17'd59320,17'd58693,17'd59189,17'd32597,17'd37985,17'd30221,17'd29646,17'd29482,17'd29198,17'd30073,17'd34381,17'd54732,17'd58935,17'd37985,17'd30678,17'd30678,17'd30372,17'd29482,17'd30373,17'd36347,17'd29336,17'd28104,17'd26629,17'd24856,17'd24030,17'd23168,17'd15184,17'd11960,17'd13883,17'd11806,17'd12861,17'd11666,17'd10736,17'd11808,17'd11398,17'd11132,17'd10164,17'd9740,17'd13887,17'd24712,17'd59437,17'd59322,17'd59438,17'd59439,17'd59440,17'd16568,17'd59441,17'd16690,17'd8580,17'd21987,17'd24368,17'd16440,17'd26498,17'd15684,17'd8724,17'd21823,17'd58696,17'd59326,17'd59193,17'd59442,17'd59443,17'd59444,17'd59445,17'd59446,17'd59447,17'd59448,17'd59449,17'd59450,17'd59082,17'd59451,17'd59452,17'd48451,17'd48046,17'd48523,17'd49978,17'd48445,17'd47629,17'd27258,17'd32006,17'd41864,17'd50154,17'd38282,17'd33318,17'd25032,17'd29243,17'd23566,17'd37117,17'd30425,17'd23217,17'd29374,17'd34137,17'd23731,17'd34467,17'd24742,17'd30126,17'd35159,17'd29534,17'd23917,17'd30879,17'd28722,17'd24086,17'd23732,17'd23733,17'd29242,17'd23386,17'd32191,17'd29973,17'd41419,17'd22859,17'd22333,17'd30276,17'd41273,17'd23217,17'd32008,17'd31828,17'd38980,17'd51160,17'd59453,17'd59454,17'd52815,17'd59337,17'd59455,17'd59456,17'd58825,17'd58461,17'd58327,17'd50465,17'd52888,17'd38282,17'd31034,17'd25320,17'd27637,17'd25568,17'd27511,17'd28369,17'd27765,17'd28597,17'd28598,17'd27638,17'd27638,17'd28720,17'd28723,17'd28720,17'd28130,17'd28597,17'd25709,17'd28850,17'd38812,17'd38812,17'd59457,17'd26531,17'd59340,17'd59340,17'd59458,17'd59459,17'd32848,17'd59212,17'd59460,17'd31360,17'd42161,17'd33944,17'd51379,17'd56641,17'd59461,17'd59462,17'd59463,17'd59464,17'd59465,17'd59466,17'd59467,17'd59468,17'd59469,17'd59470,17'd59471,17'd59472,17'd59473,17'd59474,17'd59475,17'd59476,17'd59477,17'd59478,17'd59479,17'd20974,17'd22055,17'd55451,17'd22739,17'd23620,17'd23106,17'd55644,17'd23275,17'd55862,17'd8289,17'd24476,17'd4680,17'd5322,17'd5145,17'd33532,17'd47470,17'd33992,17'd33838,17'd41891,17'd5155,17'd4846,17'd5161,17'd36887,17'd6554,17'd37152,17'd31891,17'd30333,17'd5004,17'd5005,17'd4846,17'd58971,17'd55456,17'd59480,17'd59229,17'd59481,17'd36445,17'd59482,17'd59483,17'd49708,17'd59112,17'd58850,17'd59232,17'd20704,17'd36893,17'd37159,17'd58610,17'd59367,17'd58484,17'd58977,17'd59484,17'd59368,17'd3047,17'd39323,17'd45781,17'd46990,17'd50286,17'd48553,17'd47267,17'd59370,17'd59236,17'd58619,17'd59485,17'd59486,17'd53797,17'd59487,17'd56774,17'd56774,17'd53739,17'd59241,17'd57234,17'd59488,17'd58999,17'd59489,17'd59490,17'd59491,17'd25783,17'd462,17'd20008,17'd41316,17'd1114,17'd1256,17'd1243,17'd1243,17'd9942,17'd409,17'd41316,17'd17787,17'd261,17'd426,17'd260,17'd1823,17'd2740,17'd7027,17'd27094,17'd29037,17'd29610,17'd27708,17'd31101,17'd27949,17'd11061,17'd6095,17'd5939,17'd38717,17'd38718,17'd4228,17'd59492,17'd4396,17'd4554,17'd59128,17'd59493,17'd59494,17'd19237,17'd59495,17'd53063,17'd57100,17'd59377,17'd59378,17'd59488,17'd56322,17'd58376,17'd57617
},
'{
17'd2426,17'd2258,17'd2258,17'd2597,17'd2257,17'd1414,17'd17,17'd16,17'd19,17'd10,17'd808,17'd10,17'd19,17'd18,17'd16,17'd16,17'd1416,17'd1414,17'd1414,17'd2597,17'd2935,17'd2593,17'd2782,17'd3101,17'd59496,17'd10547,17'd2426,17'd2425,17'd809,17'd289,17'd468,17'd1129,17'd11072,17'd11888,17'd59133,17'd59133,17'd295,17'd814,17'd59497,17'd45,17'd59498,17'd59001,17'd59499,17'd56791,17'd57003,17'd59500,17'd57006,17'd57113,17'd59501,17'd1294,17'd1157,17'd1298,17'd58385,17'd59502,17'd2126,17'd2271,17'd59503,17'd59504,17'd2279,17'd16148,17'd59505,17'd59006,17'd59506,17'd59507,17'd59508,17'd59509,17'd59510,17'd21966,17'd5410,17'd5090,17'd58267,17'd58392,17'd57501,17'd59511,17'd53449,17'd4771,17'd3300,17'd4128,17'd59512,17'd59513,17'd53234,17'd3301,17'd3790,17'd59514,17'd58270,17'd53608,17'd53607,17'd58765,17'd53523,17'd58397,17'd54020,17'd58272,17'd54614,17'd58649,17'd59515,17'd59516,17'd56912,17'd59517,17'd57778,17'd59283,17'd57778,17'd59274,17'd59518,17'd59519,17'd59279,17'd59520,17'd56584,17'd59521,17'd59522,17'd57779,17'd59523,17'd59524,17'd58661,17'd59525,17'd59526,17'd59284,17'd59527,17'd879,17'd59528,17'd3988,17'd59529,17'd59530,17'd59531,17'd59532,17'd59533,17'd59534,17'd59535,17'd59536,17'd59537,17'd59538,17'd56044,17'd57153,17'd57668,17'd58424,17'd59297,17'd59418,17'd59539,17'd59297,17'd59540,17'd59541,17'd59542,17'd59543,17'd59544,17'd59545,17'd59546,17'd59547,17'd59548,17'd59423,17'd59549,17'd59178,17'd59425,17'd59550,17'd59551,17'd59552,17'd59553,17'd59554,17'd59555,17'd59556,17'd59430,17'd59557,17'd59558,17'd59559,17'd59560,17'd59561,17'd59562,17'd59563,17'd57053,17'd13501,17'd57433,17'd59564,17'd58568,17'd56497,17'd56616,17'd56844,17'd31135,17'd58806,17'd32130,17'd59320,17'd57553,17'd58312,17'd30678,17'd30372,17'd30372,17'd36211,17'd29482,17'd29198,17'd30073,17'd34704,17'd58935,17'd54732,17'd32597,17'd30678,17'd30678,17'd29785,17'd29482,17'd28944,17'd50213,17'd29336,17'd28103,17'd27121,17'd25925,17'd25671,17'd16203,17'd15184,17'd11960,17'd13883,17'd11806,17'd13253,17'd14262,17'd11808,17'd11668,17'd11399,17'd11133,17'd9739,17'd27003,17'd8874,17'd11967,17'd15947,17'd54737,17'd59565,17'd59566,17'd59567,17'd10748,17'd59568,17'd9197,17'd8419,17'd25147,17'd24368,17'd24212,17'd26498,17'd29637,17'd8569,17'd22474,17'd58696,17'd59569,17'd25537,17'd59570,17'd59443,17'd59571,17'd59572,17'd59573,17'd59574,17'd59575,17'd59576,17'd59450,17'd59577,17'd59204,17'd59578,17'd48451,17'd49690,17'd47627,17'd46203,17'd42597,17'd43837,17'd31351,17'd42437,17'd51746,17'd50154,17'd43553,17'd33483,17'd28977,17'd29972,17'd23387,17'd36426,17'd39131,17'd23389,17'd30128,17'd29099,17'd30879,17'd29100,17'd24090,17'd23916,17'd30431,17'd31033,17'd23732,17'd23732,17'd23733,17'd29376,17'd23566,17'd29530,17'd29374,17'd37117,17'd30425,17'd41419,17'd45037,17'd23573,17'd22681,17'd30276,17'd23389,17'd23215,17'd29974,17'd31655,17'd31341,17'd51160,17'd53192,17'd58824,17'd39133,17'd46550,17'd59579,17'd59580,17'd59581,17'd59582,17'd57199,17'd50647,17'd38406,17'd39443,17'd25320,17'd28596,17'd27637,17'd25438,17'd25438,17'd28369,17'd25567,17'd28597,17'd28598,17'd28594,17'd28594,17'd28720,17'd28723,17'd28720,17'd28130,17'd25709,17'd28717,17'd28850,17'd59583,17'd38812,17'd59457,17'd59212,17'd59341,17'd59458,17'd59211,17'd31211,17'd32848,17'd59342,17'd59584,17'd39596,17'd43843,17'd21845,17'd59585,17'd59586,17'd51921,17'd59587,17'd59588,17'd59589,17'd59590,17'd59591,17'd59592,17'd59593,17'd59594,17'd59595,17'd59596,17'd59597,17'd59598,17'd59599,17'd59600,17'd59601,17'd59602,17'd59603,17'd59604,17'd20974,17'd21286,17'd22922,17'd53731,17'd56875,17'd23106,17'd55644,17'd23275,17'd59605,17'd7658,17'd6381,17'd24796,17'd5322,17'd4681,17'd38058,17'd47470,17'd33841,17'd33841,17'd41891,17'd4526,17'd5157,17'd5161,17'd37434,17'd6390,17'd31717,17'd31553,17'd5004,17'd5002,17'd5005,17'd4847,17'd49895,17'd4200,17'd59362,17'd59229,17'd58849,17'd59482,17'd59606,17'd59606,17'd49298,17'd58484,17'd58731,17'd59232,17'd59607,17'd36893,17'd53001,17'd59608,17'd57351,17'd58850,17'd59609,17'd20857,17'd47084,17'd59610,17'd3047,17'd59611,17'd59612,17'd59613,17'd59614,17'd46697,17'd59370,17'd44266,17'd42328,17'd59615,17'd57357,17'd57357,17'd57357,17'd59239,17'd53739,17'd58986,17'd58741,17'd56321,17'd58999,17'd53868,17'd59616,17'd56328,17'd20398,17'd1087,17'd1822,17'd3100,17'd208,17'd59617,17'd1262,17'd1823,17'd1823,17'd8315,17'd8812,17'd426,17'd59618,17'd426,17'd259,17'd425,17'd192,17'd2575,17'd6721,17'd29169,17'd29610,17'd27708,17'd31101,17'd31101,17'd33051,17'd8507,17'd37445,17'd51671,17'd38717,17'd38857,17'd38857,17'd59619,17'd4865,17'd4865,17'd59620,17'd58627,17'd59621,17'd22778,17'd59495,17'd59622,17'd57100,17'd59377,17'd59378,17'd59623,17'd56322,17'd58377,17'd59624
},
'{
17'd291,17'd59625,17'd2258,17'd2597,17'd2257,17'd1414,17'd16,17'd3905,17'd1128,17'd10,17'd808,17'd10,17'd11,17'd11,17'd19,17'd16,17'd17,17'd1414,17'd2257,17'd2597,17'd2422,17'd2784,17'd2935,17'd3101,17'd3251,17'd37047,17'd10546,17'd52621,17'd30,17'd468,17'd289,17'd290,17'd3752,17'd10924,17'd59133,17'd15878,17'd16392,17'd659,17'd14599,17'd58505,17'd58255,17'd59626,17'd59627,17'd56792,17'd56438,17'd56438,17'd57006,17'd1293,17'd1293,17'd57252,17'd59628,17'd59628,17'd1432,17'd59629,17'd56797,17'd17555,17'd59630,17'd59631,17'd3274,17'd58877,17'd18282,17'd59258,17'd59632,17'd59633,17'd59634,17'd59635,17'd59636,17'd59637,17'd20887,17'd5410,17'd4464,17'd4123,17'd59638,17'd59639,17'd59640,17'd59641,17'd59642,17'd3781,17'd59390,17'd4462,17'd59643,17'd4466,17'd3141,17'd3635,17'd59644,17'd59645,17'd58270,17'd53608,17'd58270,17'd53756,17'd54093,17'd57773,17'd55775,17'd55776,17'd59646,17'd55381,17'd58152,17'd57132,17'd56697,17'd59647,17'd59648,17'd59649,17'd56697,17'd57391,17'd59650,17'd59651,17'd59652,17'd59653,17'd59399,17'd59654,17'd58042,17'd59655,17'd59656,17'd59657,17'd59026,17'd59658,17'd59404,17'd59659,17'd1187,17'd59660,17'd59661,17'd59662,17'd59663,17'd59664,17'd59665,17'd59666,17'd59667,17'd59668,17'd53614,17'd54445,17'd59669,17'd59670,17'd58546,17'd58059,17'd58548,17'd59671,17'd59672,17'd59418,17'd59673,17'd59674,17'd59675,17'd59676,17'd59677,17'd59678,17'd59545,17'd59679,17'd59680,17'd59681,17'd59682,17'd59683,17'd59550,17'd59684,17'd59685,17'd59686,17'd59687,17'd59688,17'd59689,17'd59690,17'd59691,17'd59692,17'd59432,17'd59433,17'd59693,17'd59694,17'd59695,17'd59696,17'd58072,17'd59697,17'd59698,17'd59699,17'd59700,17'd57953,17'd56616,17'd30078,17'd30978,17'd30978,17'd55942,17'd59701,17'd59701,17'd59701,17'd32129,17'd58312,17'd59702,17'd59703,17'd29648,17'd29647,17'd30371,17'd37985,17'd36214,17'd37985,17'd37985,17'd30372,17'd29785,17'd29067,17'd28461,17'd28571,17'd28572,17'd27235,17'd27234,17'd16557,17'd18200,17'd12108,17'd19408,17'd11959,17'd19920,17'd13646,17'd13253,17'd13762,17'd23337,17'd17236,17'd12863,17'd10479,17'd51790,17'd24037,17'd9345,17'd9348,17'd8578,17'd13653,17'd14533,17'd59704,17'd59705,17'd59706,17'd21989,17'd59707,17'd13376,17'd17483,17'd9196,17'd15429,17'd8886,17'd9040,17'd29637,17'd12424,17'd32923,17'd59708,17'd20049,17'd12730,17'd15065,17'd59709,17'd59710,17'd59711,17'd59712,17'd59713,17'd59714,17'd59715,17'd59716,17'd59577,17'd59717,17'd59718,17'd48152,17'd47638,17'd46661,17'd48526,17'd47927,17'd42147,17'd49273,17'd42299,17'd50264,17'd50562,17'd43553,17'd31034,17'd35159,17'd29242,17'd32351,17'd22679,17'd22678,17'd32827,17'd32351,17'd29530,17'd23732,17'd30879,17'd23731,17'd24249,17'd32186,17'd23733,17'd23565,17'd29376,17'd29530,17'd29829,17'd29974,17'd37116,17'd36986,17'd22680,17'd34458,17'd22857,17'd22857,17'd22506,17'd22860,17'd33311,17'd32827,17'd36543,17'd31828,17'd37511,17'd31828,17'd59719,17'd52074,17'd57077,17'd39440,17'd59720,17'd59721,17'd58825,17'd58583,17'd59722,17'd50465,17'd53331,17'd53557,17'd29976,17'd24897,17'd28254,17'd25178,17'd27511,17'd25317,17'd25567,17'd27765,17'd28598,17'd28598,17'd28594,17'd28723,17'd25566,17'd28720,17'd28594,17'd25176,17'd23912,17'd25709,17'd28484,17'd33345,17'd29256,17'd32690,17'd59723,17'd59724,17'd59725,17'd37406,17'd33343,17'd32690,17'd59213,17'd36287,17'd39293,17'd36985,17'd59726,17'd59727,17'd59728,17'd22866,17'd46864,17'd59729,17'd59730,17'd59731,17'd59732,17'd59733,17'd59734,17'd59735,17'd59736,17'd59737,17'd59738,17'd29138,17'd59475,17'd59739,17'd59740,17'd59741,17'd59742,17'd59742,17'd20974,17'd59743,17'd22218,17'd23791,17'd55553,17'd23796,17'd23105,17'd23451,17'd55553,17'd7659,17'd5322,17'd5912,17'd5756,17'd33991,17'd42180,17'd4189,17'd33841,17'd34657,17'd28778,17'd28418,17'd5002,17'd25627,17'd5762,17'd5337,17'd5165,17'd5009,17'd5004,17'd5005,17'd4841,17'd4526,17'd54862,17'd59744,17'd59745,17'd4203,17'd59746,17'd59747,17'd59748,17'd36037,17'd58733,17'd58850,17'd36590,17'd49004,17'd3543,17'd58612,17'd58731,17'd59749,17'd59750,17'd59751,17'd49106,17'd59752,17'd59753,17'd47084,17'd47084,17'd59754,17'd59755,17'd59756,17'd59757,17'd59758,17'd59759,17'd57740,17'd59760,17'd57357,17'd59761,17'd59762,17'd59762,17'd53667,17'd59761,17'd53739,17'd56211,17'd59763,17'd58251,17'd56670,17'd59764,17'd59765,17'd59766,17'd1088,17'd1092,17'd3100,17'd209,17'd954,17'd1396,17'd1394,17'd1272,17'd1409,17'd1111,17'd425,17'd643,17'd3746,17'd606,17'd204,17'd598,17'd12644,17'd28916,17'd28066,17'd31729,17'd31101,17'd37168,17'd36903,17'd11882,17'd5958,17'd3897,17'd5939,17'd51671,17'd5937,17'd5937,17'd38202,17'd11048,17'd39179,17'd6404,17'd3220,17'd59767,17'd23299,17'd56883,17'd59768,17'd57100,17'd59769,17'd57482,17'd56544,17'd59770,17'd59771,17'd59772
},
'{
17'd291,17'd59625,17'd2258,17'd2597,17'd2257,17'd1414,17'd16,17'd17,17'd19,17'd10,17'd808,17'd10,17'd11,17'd11,17'd19,17'd18,17'd17,17'd1414,17'd2257,17'd2257,17'd1831,17'd2422,17'd2935,17'd3101,17'd3427,17'd35619,17'd3593,17'd52621,17'd31,17'd30,17'd289,17'd1692,17'd3752,17'd10924,17'd16011,17'd15878,17'd57896,17'd58016,17'd59773,17'd59774,17'd59775,17'd59251,17'd59627,17'd59001,17'd57110,17'd56892,17'd57113,17'd57251,17'd1293,17'd57252,17'd59776,17'd59628,17'd1432,17'd57253,17'd311,17'd59777,17'd2272,17'd34009,17'd59778,17'd58635,17'd57117,17'd59505,17'd59779,17'd59387,17'd59780,17'd59781,17'd59782,17'd59783,17'd18887,17'd6134,17'd4464,17'd3785,17'd3633,17'd3957,17'd59784,17'd59785,17'd59786,17'd3137,17'd59643,17'd4288,17'd3781,17'd59787,17'd4467,17'd2987,17'd59788,17'd59644,17'd59267,17'd53608,17'd54350,17'd53756,17'd54253,17'd54347,17'd59646,17'd54347,17'd59646,17'd59789,17'd56580,17'd56909,17'd59393,17'd59790,17'd59791,17'd59648,17'd59019,17'd58036,17'd59792,17'd58660,17'd59793,17'd59794,17'd59795,17'd59796,17'd59650,17'd59655,17'd56914,17'd59797,17'd55494,17'd59798,17'd59799,17'd59800,17'd56916,17'd2501,17'd59801,17'd59802,17'd59803,17'd59804,17'd59805,17'd59806,17'd59807,17'd59808,17'd58422,17'd59809,17'd59810,17'd59811,17'd57036,17'd58179,17'd58177,17'd59812,17'd59813,17'd59814,17'd59539,17'd59815,17'd59674,17'd59816,17'd59817,17'd59677,17'd59818,17'd59819,17'd59820,17'd59302,17'd59821,17'd59822,17'd59685,17'd59823,17'd59824,17'd59825,17'd59826,17'd59827,17'd59828,17'd59829,17'd59429,17'd59830,17'd59831,17'd59832,17'd59833,17'd59834,17'd59834,17'd59835,17'd12977,17'd57546,17'd13750,17'd59836,17'd59837,17'd55416,17'd56616,17'd38365,17'd39661,17'd39661,17'd57688,17'd31949,17'd31949,17'd59838,17'd59839,17'd58077,17'd38237,17'd58693,17'd29647,17'd30372,17'd37985,17'd37985,17'd32597,17'd37985,17'd30371,17'd36937,17'd31587,17'd28686,17'd28571,17'd28818,17'd28348,17'd27348,17'd27486,17'd16913,17'd18564,17'd14807,17'd11959,17'd11960,17'd13520,17'd11667,17'd11807,17'd11397,17'd37196,17'd12584,17'd10479,17'd18196,17'd23857,17'd15180,17'd10174,17'd8724,17'd19780,17'd59840,17'd14142,17'd55217,17'd59841,17'd59842,17'd59843,17'd59844,17'd16919,17'd17352,17'd59845,17'd8413,17'd8724,17'd9040,17'd48326,17'd23517,17'd32923,17'd59321,17'd59846,17'd55030,17'd59847,17'd59848,17'd59849,17'd59850,17'd59851,17'd59852,17'd59853,17'd59854,17'd59855,17'd59856,17'd59857,17'd59718,17'd48451,17'd47443,17'd46433,17'd44477,17'd43020,17'd42147,17'd45036,17'd48784,17'd54938,17'd53841,17'd39443,17'd29103,17'd32659,17'd29827,17'd23218,17'd22678,17'd22859,17'd39131,17'd23218,17'd29829,17'd23565,17'd28722,17'd30879,17'd24087,17'd29527,17'd29241,17'd31502,17'd29530,17'd32191,17'd23389,17'd32827,17'd22330,17'd30276,17'd22332,17'd32344,17'd30426,17'd30426,17'd22506,17'd22681,17'd30276,17'd22329,17'd36543,17'd37511,17'd37511,17'd39133,17'd59719,17'd59858,17'd46096,17'd59720,17'd59859,17'd59860,17'd59861,17'd57196,17'd57840,17'd59862,17'd59863,17'd38667,17'd24895,17'd24897,17'd28254,17'd25177,17'd28369,17'd27765,17'd25567,17'd27638,17'd28598,17'd27638,17'd28720,17'd28723,17'd28723,17'd28720,17'd27765,17'd24079,17'd27882,17'd28369,17'd33814,17'd26403,17'd26176,17'd29701,17'd59864,17'd59865,17'd59866,17'd37406,17'd59867,17'd59868,17'd59869,17'd59870,17'd59871,17'd59872,17'd59873,17'd59874,17'd59875,17'd47751,17'd59876,17'd59877,17'd59878,17'd59879,17'd59880,17'd22700,17'd59881,17'd59882,17'd59883,17'd59884,17'd59885,17'd59886,17'd33521,17'd59887,17'd59888,17'd59889,17'd59742,17'd59890,17'd21117,17'd22226,17'd22392,17'd24142,17'd23454,17'd23277,17'd55348,17'd57589,17'd22933,17'd10196,17'd26217,17'd5912,17'd4681,17'd4358,17'd4358,17'd4189,17'd33841,17'd34657,17'd37432,17'd30180,17'd25627,17'd5160,17'd5762,17'd5168,17'd5163,17'd5008,17'd30637,17'd4842,17'd4841,17'd4526,17'd54227,17'd59230,17'd59482,17'd57734,17'd59365,17'd36037,17'd35900,17'd59891,17'd59892,17'd58977,17'd58977,17'd49004,17'd59232,17'd58612,17'd58731,17'd59750,17'd59234,17'd58977,17'd59893,17'd59484,17'd59894,17'd59895,17'd59753,17'd59896,17'd59897,17'd59898,17'd59899,17'd59758,17'd41309,17'd57602,17'd53738,17'd57357,17'd59761,17'd59900,17'd59900,17'd59901,17'd59902,17'd53739,17'd53740,17'd59903,17'd59904,17'd59905,17'd59906,17'd59907,17'd930,17'd784,17'd622,17'd428,17'd7512,17'd1666,17'd781,17'd1525,17'd423,17'd1099,17'd952,17'd1111,17'd425,17'd206,17'd605,17'd1272,17'd1669,17'd2394,17'd32082,17'd31562,17'd31101,17'd36905,17'd36905,17'd35487,17'd2906,17'd6581,17'd4575,17'd5939,17'd51671,17'd59908,17'd58745,17'd39327,17'd11048,17'd3872,17'd8787,17'd59909,17'd19237,17'd51333,17'd58747,17'd59622,17'd59130,17'd59769,17'd57482,17'd56544,17'd59770,17'd59771,17'd59910
},
'{
17'd982,17'd2259,17'd2258,17'd2597,17'd2425,17'd1414,17'd17,17'd3905,17'd11,17'd10,17'd808,17'd808,17'd11,17'd11,17'd18,17'd18,17'd17,17'd17,17'd1414,17'd2257,17'd1688,17'd2422,17'd2935,17'd3101,17'd3428,17'd35619,17'd10669,17'd52621,17'd1129,17'd468,17'd2938,17'd468,17'd2596,17'd10802,17'd57896,17'd15118,17'd58016,17'd58016,17'd1279,17'd59911,17'd59912,17'd59913,17'd59627,17'd56672,17'd57002,17'd56892,17'd57113,17'd57113,17'd57006,17'd1293,17'd59914,17'd58382,17'd59915,17'd57253,17'd312,17'd59916,17'd2271,17'd32887,17'd59917,17'd59004,17'd2803,17'd59918,17'd59919,17'd59920,17'd59921,17'd59922,17'd59923,17'd59924,17'd59925,17'd6134,17'd4766,17'd4924,17'd59926,17'd3464,17'd3958,17'd4929,17'd59927,17'd3135,17'd3780,17'd3946,17'd3946,17'd4466,17'd2983,17'd2982,17'd59928,17'd59929,17'd59267,17'd53523,17'd59143,17'd53880,17'd57773,17'd59646,17'd54705,17'd54895,17'd57126,17'd59930,17'd56351,17'd59931,17'd57783,17'd59024,17'd59932,17'd58527,17'd57778,17'd59933,17'd59934,17'd57922,17'd59282,17'd59935,17'd59936,17'd59937,17'd59938,17'd57518,17'd59939,17'd59937,17'd59940,17'd59941,17'd57281,17'd59942,17'd58164,17'd2501,17'd59943,17'd59944,17'd59945,17'd59946,17'd59947,17'd59948,17'd58670,17'd59949,17'd59950,17'd59951,17'd59952,17'd59953,17'd56711,17'd57668,17'd58177,17'd59041,17'd59164,17'd59954,17'd59954,17'd59673,17'd59815,17'd59955,17'd59956,17'd59957,17'd59818,17'd59958,17'd59959,17'd59960,17'd59961,17'd59962,17'd59686,17'd59824,17'd59963,17'd59964,17'd59826,17'd59965,17'd59828,17'd59966,17'd59967,17'd59968,17'd59969,17'd59970,17'd59971,17'd59972,17'd59833,17'd59973,17'd13232,17'd11930,17'd59974,17'd59975,17'd59976,17'd55609,17'd57953,17'd56616,17'd56616,17'd55699,17'd57688,17'd31949,17'd57688,17'd57688,17'd30977,17'd58077,17'd58693,17'd30531,17'd30372,17'd30678,17'd37985,17'd37985,17'd37985,17'd37985,17'd30371,17'd29647,17'd30373,17'd29645,17'd50213,17'd28572,17'd28348,17'd27348,17'd25528,17'd23855,17'd12254,17'd14807,17'd14130,17'd11960,17'd13646,17'd11807,17'd16068,17'd10990,17'd21206,17'd14134,17'd10479,17'd18196,17'd25281,17'd16318,17'd9041,17'd8572,17'd8251,17'd52875,17'd15444,17'd59977,17'd12269,17'd59978,17'd23869,17'd20613,17'd15693,17'd8252,17'd25679,17'd17481,17'd8724,17'd9348,17'd48326,17'd23517,17'd32923,17'd59979,17'd25534,17'd55030,17'd59570,17'd59848,17'd59980,17'd59981,17'd59982,17'd59983,17'd59984,17'd59985,17'd47528,17'd59986,17'd59987,17'd59988,17'd48142,17'd49580,17'd49378,17'd41864,17'd33155,17'd32995,17'd43156,17'd59989,17'd51828,17'd53841,17'd39443,17'd29244,17'd30431,17'd29686,17'd32827,17'd22677,17'd39911,17'd31656,17'd32827,17'd30128,17'd29242,17'd23384,17'd30275,17'd24086,17'd29241,17'd23733,17'd29376,17'd32191,17'd39278,17'd23740,17'd36288,17'd34458,17'd22677,17'd32344,17'd30426,17'd30426,17'd30426,17'd22506,17'd22332,17'd30276,17'd22503,17'd37116,17'd29974,17'd41587,17'd58950,17'd59719,17'd39280,17'd50732,17'd59720,17'd59990,17'd59860,17'd59206,17'd50819,17'd59991,17'd49680,17'd34113,17'd30126,17'd24744,17'd24897,17'd27637,17'd25438,17'd29101,17'd25317,17'd25567,17'd27638,17'd27638,17'd28594,17'd28723,17'd25566,17'd28723,17'd27765,17'd28597,17'd28717,17'd29101,17'd29101,17'd30903,17'd59992,17'd59993,17'd59994,17'd59995,17'd59996,17'd59997,17'd59998,17'd26783,17'd59999,17'd34636,17'd60000,17'd52327,17'd47160,17'd60001,17'd60002,17'd47549,17'd60003,17'd60004,17'd60005,17'd60006,17'd60007,17'd60008,17'd60009,17'd60010,17'd60011,17'd60012,17'd60013,17'd60014,17'd60015,17'd60016,17'd60017,17'd60018,17'd60019,17'd59890,17'd20673,17'd40541,17'd22922,17'd23620,17'd22933,17'd24306,17'd23108,17'd55348,17'd23276,17'd26111,17'd10196,17'd24649,17'd5756,17'd4681,17'd4358,17'd4358,17'd4189,17'd41891,17'd5154,17'd4684,17'd5005,17'd25627,17'd5336,17'd5762,17'd5166,17'd5009,17'd30637,17'd30180,17'd28418,17'd4684,17'd50176,17'd58608,17'd36445,17'd59482,17'd59483,17'd59483,17'd59748,17'd60020,17'd60021,17'd60022,17'd58977,17'd58977,17'd49004,17'd60023,17'd58483,17'd59609,17'd59234,17'd59234,17'd59609,17'd58732,17'd36317,17'd50179,17'd60024,17'd21319,17'd20705,17'd52452,17'd60025,17'd50590,17'd59370,17'd41900,17'd57355,17'd53738,17'd57232,17'd59761,17'd60026,17'd59900,17'd53667,17'd58986,17'd58241,17'd60027,17'd58874,17'd60028,17'd56998,17'd60029,17'd18758,17'd24496,17'd1379,17'd1257,17'd627,17'd954,17'd1396,17'd604,17'd1408,17'd598,17'd951,17'd603,17'd191,17'd1111,17'd643,17'd971,17'd422,17'd415,17'd26965,17'd29037,17'd27949,17'd31101,17'd60030,17'd36904,17'd11882,17'd2906,17'd6581,17'd4713,17'd3423,17'd51671,17'd58745,17'd39948,17'd38334,17'd5355,17'd4864,17'd60031,17'd60032,17'd22778,17'd40560,17'd52532,17'd60033,17'd60034,17'd57605,17'd57482,17'd57482,17'd2072,17'd54510,17'd60035
},
'{
17'd982,17'd2259,17'd2258,17'd2597,17'd2258,17'd2257,17'd17,17'd17,17'd19,17'd10,17'd808,17'd808,17'd11,17'd1128,17'd18,17'd18,17'd16,17'd17,17'd1414,17'd2257,17'd1688,17'd2422,17'd2935,17'd3101,17'd3428,17'd35619,17'd10670,17'd10547,17'd291,17'd30,17'd468,17'd468,17'd2596,17'd10669,17'd16392,17'd15118,17'd15118,17'd58504,17'd1279,17'd15497,17'd60036,17'd60037,17'd60038,17'd60039,17'd56891,17'd60040,17'd57006,17'd57113,17'd57006,17'd1292,17'd57899,17'd60041,17'd58382,17'd57253,17'd312,17'd56797,17'd56562,17'd32733,17'd34803,17'd58753,17'd21172,17'd16148,17'd59505,17'd60042,17'd60043,17'd60044,17'd58880,17'd60045,17'd60046,17'd21966,17'd4928,17'd5250,17'd4293,17'd3299,17'd2976,17'd4297,17'd60047,17'd60048,17'd3295,17'd3471,17'd3300,17'd59642,17'd2982,17'd2825,17'd4931,17'd4297,17'd59514,17'd53523,17'd59143,17'd58028,17'd54532,17'd54530,17'd59930,17'd59930,17'd57506,17'd58273,17'd60049,17'd58152,17'd60050,17'd58160,17'd59019,17'd60051,17'd60052,17'd56914,17'd57784,17'd59792,17'd60053,17'd58156,17'd60054,17'd60055,17'd60056,17'd60057,17'd60058,17'd60059,17'd60060,17'd55681,17'd60061,17'd60062,17'd58164,17'd60063,17'd60064,17'd1606,17'd59028,17'd59289,17'd60065,17'd60066,17'd57145,17'd60067,17'd60068,17'd60069,17'd60070,17'd60071,17'd56472,17'd57932,17'd58177,17'd59041,17'd60072,17'd60073,17'd60074,17'd59296,17'd59297,17'd60075,17'd59676,17'd60076,17'd59957,17'd60077,17'd59959,17'd60078,17'd60079,17'd60080,17'd60081,17'd59963,17'd60082,17'd60083,17'd60084,17'd60085,17'd60086,17'd60087,17'd60088,17'd60089,17'd60090,17'd60091,17'd59557,17'd60092,17'd60093,17'd59560,17'd60094,17'd60095,17'd60096,17'd15801,17'd60097,17'd58931,17'd58076,17'd60098,17'd56616,17'd18685,17'd56947,17'd57688,17'd57688,17'd59838,17'd58077,17'd58077,17'd30531,17'd30680,17'd30678,17'd30678,17'd37985,17'd37985,17'd37985,17'd30371,17'd57554,17'd29646,17'd30373,17'd29645,17'd50213,17'd28350,17'd27349,17'd26373,17'd18200,17'd12254,17'd12579,17'd14130,17'd11960,17'd13366,17'd11667,17'd16068,17'd14931,17'd11132,17'd15176,17'd11527,17'd9883,17'd17011,17'd13887,17'd8721,17'd8724,17'd24213,17'd9622,17'd15059,17'd15307,17'd60099,17'd23875,17'd60100,17'd60101,17'd14530,17'd16802,17'd16691,17'd8733,17'd17481,17'd8725,17'd9348,17'd48326,17'd22473,17'd32923,17'd59979,17'd25534,17'd55030,17'd59570,17'd60102,17'd60103,17'd60104,17'd60105,17'd60106,17'd60107,17'd60108,17'd48032,17'd47528,17'd60109,17'd60110,17'd49270,17'd60111,17'd51561,17'd43548,17'd44231,17'd32995,17'd42884,17'd52260,17'd52426,17'd48895,17'd39443,17'd29244,17'd24249,17'd29374,17'd39131,17'd22857,17'd52752,17'd39911,17'd39131,17'd32351,17'd23386,17'd29689,17'd23564,17'd23733,17'd23733,17'd29376,17'd29686,17'd37117,17'd32830,17'd36288,17'd22859,17'd22677,17'd30426,17'd30426,17'd30427,17'd30427,17'd30426,17'd22677,17'd22856,17'd22331,17'd22503,17'd37116,17'd29974,17'd31828,17'd59719,17'd56397,17'd37116,17'd36543,17'd60112,17'd60113,17'd52502,17'd59083,17'd51307,17'd51735,17'd49680,17'd28977,17'd23561,17'd28595,17'd28596,17'd25320,17'd28850,17'd25317,17'd27765,17'd25567,17'd27638,17'd28594,17'd28723,17'd25566,17'd25566,17'd28720,17'd25567,17'd25709,17'd25177,17'd32689,17'd59457,17'd59999,17'd60114,17'd27261,17'd60115,17'd60116,17'd42156,17'd38825,17'd26783,17'd60117,17'd32373,17'd60118,17'd57847,17'd31660,17'd60119,17'd60120,17'd60121,17'd49796,17'd60122,17'd60123,17'd60124,17'd30458,17'd60125,17'd60126,17'd60127,17'd60128,17'd60129,17'd60130,17'd60131,17'd60132,17'd54952,17'd60133,17'd60134,17'd56984,17'd60135,17'd20673,17'd20974,17'd60136,17'd58231,17'd30028,17'd24792,17'd24306,17'd23277,17'd55986,17'd60137,17'd22587,17'd7007,17'd60138,17'd4992,17'd4837,17'd34157,17'd33991,17'd4189,17'd41891,17'd28778,17'd29024,17'd25627,17'd5160,17'd5762,17'd5336,17'd5163,17'd5009,17'd30180,17'd28418,17'd4684,17'd39015,17'd50588,17'd60139,17'd36313,17'd60140,17'd59747,17'd59606,17'd59748,17'd60020,17'd60141,17'd60141,17'd58732,17'd58732,17'd3543,17'd60142,17'd58483,17'd59609,17'd59234,17'd59234,17'd50178,17'd50285,17'd3543,17'd59484,17'd48728,17'd48728,17'd59896,17'd48382,17'd50590,17'd46879,17'd45182,17'd42192,17'd57884,17'd57097,17'd60143,17'd57357,17'd60144,17'd60026,17'd60145,17'd53739,17'd56663,17'd55072,17'd53937,17'd58375,17'd55887,17'd60146,17'd34510,17'd52104,17'd798,17'd226,17'd626,17'd1256,17'd3743,17'd192,17'd598,17'd193,17'd951,17'd193,17'd1668,17'd411,17'd425,17'd411,17'd951,17'd1672,17'd29037,17'd29610,17'd31729,17'd31101,17'd60030,17'd60030,17'd34002,17'd11061,17'd6416,17'd4883,17'd5182,17'd5938,17'd38202,17'd38334,17'd38334,17'd18383,17'd6404,17'd58008,17'd60147,17'd39324,17'd40714,17'd60148,17'd60149,17'd57605,17'd59769,17'd57482,17'd57482,17'd2072,17'd54510,17'd54082
},
'{
17'd982,17'd2259,17'd3752,17'd2597,17'd2258,17'd2257,17'd17,17'd3905,17'd11,17'd10,17'd808,17'd808,17'd10,17'd1128,17'd18,17'd18,17'd16,17'd17,17'd1416,17'd2257,17'd1688,17'd1831,17'd3252,17'd2935,17'd3427,17'd60150,17'd54978,17'd10547,17'd2426,17'd1414,17'd1692,17'd468,17'd1414,17'd52621,17'd16501,17'd15118,17'd14989,17'd14989,17'd986,17'd15362,17'd58505,17'd47,17'd59626,17'd56891,17'd60151,17'd60152,17'd1292,17'd57006,17'd1430,17'd57006,17'd57113,17'd57899,17'd59914,17'd57253,17'd492,17'd60153,17'd60154,17'd23491,17'd32887,17'd2131,17'd2278,17'd2803,17'd18045,17'd60155,17'd60156,17'd60157,17'd60158,17'd60159,17'd60160,17'd5995,17'd5256,17'd5688,17'd3950,17'd3299,17'd3133,17'd2648,17'd4616,17'd60161,17'd2824,17'd3468,17'd3139,17'd53303,17'd60162,17'd60163,17'd60164,17'd2649,17'd60165,17'd59269,17'd60166,17'd53522,17'd60167,17'd60168,17'd60169,17'd60170,17'd60171,17'd60172,17'd60173,17'd56351,17'd60174,17'd60175,17'd60176,17'd57778,17'd59793,17'd59276,17'd57784,17'd59655,17'd58654,17'd60177,17'd60178,17'd60179,17'd60180,17'd60181,17'd60182,17'd60183,17'd59394,17'd60184,17'd59940,17'd56246,17'd60185,17'd60186,17'd60187,17'd59405,17'd709,17'd60188,17'd60189,17'd60190,17'd60191,17'd60192,17'd60193,17'd53959,17'd60194,17'd60195,17'd60196,17'd60197,17'd60198,17'd60199,17'd60200,17'd58912,17'd60201,17'd60202,17'd59814,17'd60203,17'd60204,17'd60076,17'd60205,17'd60077,17'd60206,17'd60207,17'd60208,17'd60209,17'd60210,17'd60211,17'd60212,17'd60213,17'd60084,17'd60214,17'd60215,17'd60086,17'd59688,17'd59829,17'd60216,17'd60217,17'd60218,17'd60219,17'd58924,17'd60220,17'd58800,17'd60221,17'd60222,17'd60223,17'd60224,17'd60225,17'd55316,17'd60226,17'd60227,17'd19031,17'd56272,17'd55942,17'd57688,17'd59701,17'd59839,17'd32129,17'd30681,17'd59189,17'd30678,17'd37985,17'd37985,17'd37985,17'd29785,17'd30220,17'd29646,17'd36211,17'd30373,17'd36347,17'd28572,17'd28348,17'd27348,17'd27486,17'd23855,17'd12108,17'd20314,17'd18198,17'd13135,17'd11807,17'd16069,17'd17236,17'd11132,17'd10326,17'd11670,17'd9883,17'd11136,17'd9346,17'd9038,17'd8569,17'd15429,17'd8419,17'd35371,17'd39823,17'd15062,17'd21992,17'd8431,17'd59706,17'd59071,17'd7294,17'd16802,17'd7947,17'd8418,17'd9349,17'd8725,17'd8878,17'd60228,17'd22473,17'd60229,17'd59979,17'd60230,17'd60231,17'd60232,17'd60233,17'd60234,17'd60235,17'd60236,17'd60237,17'd60238,17'd60239,17'd48032,17'd59855,17'd49972,17'd60240,17'd57073,17'd51556,17'd46203,17'd47334,17'd32995,17'd49273,17'd48258,17'd50152,17'd52426,17'd53841,17'd39443,17'd30432,17'd24087,17'd37386,17'd22678,17'd22161,17'd31657,17'd35711,17'd34458,17'd30277,17'd29686,17'd29827,17'd29099,17'd31502,17'd29099,17'd23387,17'd32191,17'd23216,17'd32827,17'd22331,17'd22856,17'd22333,17'd30426,17'd22161,17'd22158,17'd30427,17'd30426,17'd22677,17'd30276,17'd22500,17'd22503,17'd37116,17'd37511,17'd31655,17'd57077,17'd39440,17'd22503,17'd39588,17'd60241,17'd59721,17'd60242,17'd59454,17'd50819,17'd57205,17'd50364,17'd28601,17'd29240,17'd34283,17'd28254,17'd29244,17'd29101,17'd25317,17'd25567,17'd28597,17'd27638,17'd28720,17'd25566,17'd25566,17'd25435,17'd28130,17'd28597,17'd25709,17'd34127,17'd38812,17'd33345,17'd29256,17'd32524,17'd60243,17'd59995,17'd31846,17'd31364,17'd29992,17'd32524,17'd60244,17'd59869,17'd55960,17'd50165,17'd41112,17'd52439,17'd51068,17'd60245,17'd60246,17'd60247,17'd60248,17'd60249,17'd60250,17'd23233,17'd22879,17'd60251,17'd60252,17'd60253,17'd60254,17'd33189,17'd60255,17'd60256,17'd60257,17'd60258,17'd60259,17'd21277,17'd60260,17'd60261,17'd60262,17'd22565,17'd55740,17'd24305,17'd24306,17'd23277,17'd56655,17'd24793,17'd8608,17'd6545,17'd5325,17'd4682,17'd4838,17'd34157,17'd33991,17'd4189,17'd41891,17'd5327,17'd5002,17'd5160,17'd28185,17'd5762,17'd5335,17'd5008,17'd5008,17'd4842,17'd4685,17'd49995,17'd50176,17'd60263,17'd60264,17'd6566,17'd6566,17'd60265,17'd35899,17'd35900,17'd60020,17'd60141,17'd60141,17'd60266,17'd60267,17'd59484,17'd59113,17'd58483,17'd59609,17'd36446,17'd36446,17'd36446,17'd50285,17'd59232,17'd20857,17'd36450,17'd60268,17'd52452,17'd48182,17'd60269,17'd59370,17'd41900,17'd60270,17'd59760,17'd57231,17'd57231,17'd57356,17'd60271,17'd60271,17'd59761,17'd53798,17'd60027,17'd54972,17'd1927,17'd60272,17'd55565,17'd60273,17'd1809,17'd451,17'd234,17'd3248,17'd626,17'd1666,17'd604,17'd6868,17'd193,17'd193,17'd951,17'd193,17'd603,17'd971,17'd606,17'd1272,17'd194,17'd777,17'd2741,17'd29610,17'd31729,17'd31101,17'd36905,17'd36905,17'd33051,17'd11061,17'd6416,17'd4729,17'd3424,17'd5182,17'd38203,17'd41481,17'd11867,17'd41160,17'd50841,17'd18981,17'd60274,17'd39324,17'd56547,17'd60148,17'd60149,17'd57605,17'd60275,17'd2070,17'd2070,17'd59903,17'd60276,17'd60277
},
'{
17'd982,17'd982,17'd3752,17'd3752,17'd2258,17'd2258,17'd1415,17'd17,17'd19,17'd10,17'd808,17'd808,17'd10,17'd1128,17'd18,17'd19,17'd16,17'd17,17'd1416,17'd1416,17'd4247,17'd1688,17'd2422,17'd2935,17'd3427,17'd60150,17'd59496,17'd10802,17'd10547,17'd2596,17'd2599,17'd468,17'd1414,17'd3429,17'd11888,17'd58016,17'd14989,17'd14989,17'd58016,17'd986,17'd59911,17'd60278,17'd60279,17'd60280,17'd60281,17'd60152,17'd1152,17'd1292,17'd57005,17'd1430,17'd57006,17'd57113,17'd1562,17'd78,17'd77,17'd60153,17'd59777,17'd2617,17'd60282,17'd60283,17'd59917,17'd21172,17'd3770,17'd60284,17'd60042,17'd60285,17'd60286,17'd60287,17'd4454,17'd60288,17'd60289,17'd4928,17'd60290,17'd3946,17'd3293,17'd60291,17'd4774,17'd53610,17'd5695,17'd60292,17'd3136,17'd3136,17'd60293,17'd60294,17'd60295,17'd4932,17'd4929,17'd60296,17'd60166,17'd53607,17'd54435,17'd60297,17'd60298,17'd60299,17'd56688,17'd54892,17'd55093,17'd58522,17'd60300,17'd60301,17'd58160,17'd60302,17'd60303,17'd59793,17'd60304,17'd57784,17'd59024,17'd60305,17'd60306,17'd60179,17'd56698,17'd60307,17'd60305,17'd60305,17'd60308,17'd60309,17'd59657,17'd60310,17'd56586,17'd60311,17'd60312,17'd60313,17'd60314,17'd60315,17'd60316,17'd60317,17'd60318,17'd60319,17'd60320,17'd60321,17'd59536,17'd60070,17'd60322,17'd60323,17'd60324,17'd60199,17'd60325,17'd58787,17'd60326,17'd60327,17'd60328,17'd60203,17'd60329,17'd60330,17'd60205,17'd60205,17'd60206,17'd60331,17'd60332,17'd60078,17'd60333,17'd60334,17'd60335,17'd60335,17'd60336,17'd60337,17'd60338,17'd60215,17'd60339,17'd60340,17'd60341,17'd60342,17'd60343,17'd59692,17'd59831,17'd58924,17'd59056,17'd60344,17'd60345,17'd60346,17'd60347,17'd54276,17'd57057,17'd57953,17'd60227,17'd19031,17'd17844,17'd56272,17'd57688,17'd31950,17'd59839,17'd30681,17'd59189,17'd30680,17'd37985,17'd37985,17'd30371,17'd30371,17'd30220,17'd29646,17'd36211,17'd29481,17'd30373,17'd36347,17'd28572,17'd27235,17'd27486,17'd23855,17'd12108,17'd21671,17'd11959,17'd14261,17'd11667,17'd16068,17'd17838,17'd13886,17'd11133,17'd10479,17'd9883,17'd9741,17'd10744,17'd8874,17'd25677,17'd8731,17'd8578,17'd18203,17'd18085,17'd19419,17'd19421,17'd60348,17'd24052,17'd59706,17'd60349,17'd24868,17'd11534,17'd17241,17'd19780,17'd9887,17'd24368,17'd8878,17'd60228,17'd10607,17'd34829,17'd59979,17'd60230,17'd60350,17'd55954,17'd60351,17'd60352,17'd60353,17'd60354,17'd60355,17'd60356,17'd60357,17'd58326,17'd59333,17'd60358,17'd49471,17'd55038,17'd51645,17'd50825,17'd46753,17'd32995,17'd49273,17'd48612,17'd46202,17'd50360,17'd59209,17'd38406,17'd29533,17'd31033,17'd23217,17'd22332,17'd22161,17'd31657,17'd31657,17'd23573,17'd22329,17'd29828,17'd23386,17'd29376,17'd35865,17'd35865,17'd30579,17'd23569,17'd22501,17'd22327,17'd22325,17'd22681,17'd22159,17'd22159,17'd22161,17'd22161,17'd30426,17'd23573,17'd22332,17'd22330,17'd22328,17'd22501,17'd37116,17'd41587,17'd31828,17'd51552,17'd33158,17'd22502,17'd60359,17'd60360,17'd50815,17'd51473,17'd58824,17'd50730,17'd60361,17'd23917,17'd23562,17'd29240,17'd28596,17'd25320,17'd27511,17'd25317,17'd27765,17'd25567,17'd25567,17'd28594,17'd28723,17'd25566,17'd25566,17'd28600,17'd25567,17'd28597,17'd25709,17'd30903,17'd29256,17'd29256,17'd60362,17'd32524,17'd32038,17'd60363,17'd42156,17'd60364,17'd60365,17'd60366,17'd60367,17'd60368,17'd60369,17'd21694,17'd57974,17'd60370,17'd60371,17'd48627,17'd60372,17'd60373,17'd60374,17'd36563,17'd60375,17'd23408,17'd60376,17'd60377,17'd60378,17'd60379,17'd60380,17'd43035,17'd60381,17'd60382,17'd60383,17'd60384,17'd60385,17'd20972,17'd29422,17'd21895,17'd29882,17'd23619,17'd53503,17'd24792,17'd24306,17'd23277,17'd23455,17'd60386,17'd26449,17'd6546,17'd5325,17'd4682,17'd5144,17'd33991,17'd33838,17'd33841,17'd41459,17'd4686,17'd5004,17'd28185,17'd27935,17'd5336,17'd25627,17'd37029,17'd37288,17'd28418,17'd4685,17'd60387,17'd56203,17'd60388,17'd60389,17'd60390,17'd60391,17'd6400,17'd4209,17'd49709,17'd35900,17'd60392,17'd3545,17'd49998,17'd60267,17'd60393,17'd60393,17'd3543,17'd58977,17'd36446,17'd36446,17'd58484,17'd58357,17'd58483,17'd3543,17'd20857,17'd59754,17'd48182,17'd59369,17'd46879,17'd58122,17'd42192,17'd60270,17'd60394,17'd57231,17'd57231,17'd57356,17'd60271,17'd60145,17'd60395,17'd56663,17'd55266,17'd59903,17'd60396,17'd60397,17'd55885,17'd19361,17'd8788,17'd448,17'd447,17'd626,17'd1263,17'd4727,17'd6868,17'd2409,17'd602,17'd602,17'd951,17'd193,17'd603,17'd424,17'd606,17'd1272,17'd778,17'd1949,17'd29610,17'd29610,17'd31101,17'd31101,17'd36905,17'd37168,17'd34002,17'd9124,17'd35769,17'd60398,17'd5182,17'd38203,17'd44019,17'd60399,17'd39032,17'd3871,17'd50002,17'd60400,17'd60401,17'd58374,17'd40258,17'd60402,17'd60403,17'd57482,17'd2071,17'd2070,17'd2071,17'd59903,17'd60276,17'd60277
},
'{
17'd3429,17'd3429,17'd3752,17'd3752,17'd2426,17'd2425,17'd1416,17'd1416,17'd19,17'd19,17'd10,17'd808,17'd10,17'd1128,17'd18,17'd19,17'd18,17'd3905,17'd1416,17'd1416,17'd4247,17'd1688,17'd2422,17'd2935,17'd2934,17'd35619,17'd54242,17'd10802,17'd12195,17'd2596,17'd2599,17'd809,17'd22965,17'd2258,17'd3751,17'd4893,17'd15117,17'd14989,17'd58016,17'd659,17'd15497,17'd60404,17'd59913,17'd60039,17'd60281,17'd60152,17'd1152,17'd57372,17'd57005,17'd1430,17'd59500,17'd57111,17'd57898,17'd77,17'd59629,17'd60405,17'd59916,17'd2440,17'd41162,17'd60406,17'd34170,17'd21640,17'd3276,17'd60407,17'd60408,17'd60409,17'd60410,17'd3614,17'd60411,17'd60412,17'd22461,17'd5256,17'd4768,17'd3949,17'd3136,17'd60291,17'd60413,17'd60414,17'd60415,17'd53815,17'd5690,17'd2984,17'd60416,17'd60294,17'd60417,17'd60164,17'd4772,17'd60418,17'd60419,17'd58765,17'd60420,17'd60421,17'd60169,17'd60422,17'd57015,17'd56351,17'd56689,17'd60049,17'd60422,17'd60423,17'd58408,17'd59523,17'd59147,17'd60303,17'd59025,17'd59150,17'd56697,17'd58157,17'd60424,17'd60425,17'd60426,17'd56355,17'd60427,17'd60428,17'd57644,17'd57778,17'd60060,17'd60429,17'd59798,17'd58285,17'd60430,17'd60431,17'd60432,17'd3020,17'd60433,17'd60434,17'd60435,17'd60436,17'd60437,17'd60438,17'd60439,17'd60440,17'd60441,17'd60442,17'd60443,17'd58547,17'd60444,17'd58787,17'd60326,17'd60445,17'd60328,17'd60446,17'd60447,17'd60448,17'd60449,17'd60205,17'd60450,17'd60451,17'd60331,17'd60452,17'd60453,17'd60454,17'd60455,17'd60456,17'd60457,17'd60458,17'd60459,17'd60338,17'd60338,17'd60339,17'd60087,17'd60460,17'd60216,17'd60461,17'd60462,17'd60463,17'd59313,17'd59315,17'd13116,17'd57545,17'd12707,17'd60464,17'd54645,17'd59436,17'd60465,17'd18685,17'd38910,17'd38910,17'd57688,17'd59701,17'd58077,17'd32129,17'd58932,17'd30680,17'd30372,17'd30372,17'd29647,17'd29647,17'd29482,17'd30373,17'd29481,17'd29481,17'd36347,17'd28572,17'd27235,17'd27234,17'd23855,17'd12254,17'd14807,17'd11959,17'd11961,17'd13764,17'd16069,17'd17236,17'd10477,17'd11528,17'd9739,17'd15048,17'd10742,17'd16554,17'd9339,17'd9038,17'd9046,17'd21987,17'd17352,17'd13006,17'd25004,17'd19647,17'd16807,17'd60466,17'd8431,17'd12431,17'd60349,17'd41932,17'd14932,17'd17241,17'd10028,17'd9349,17'd8726,17'd8879,17'd50864,17'd8572,17'd34829,17'd59979,17'd60467,17'd60468,17'd60469,17'd60470,17'd60471,17'd60472,17'd60473,17'd60474,17'd60475,17'd60357,17'd60476,17'd49675,17'd60477,17'd56970,17'd48033,17'd60478,17'd51653,17'd46753,17'd49273,17'd47438,17'd48784,17'd49274,17'd56636,17'd59209,17'd38406,17'd29533,17'd23920,17'd23389,17'd22333,17'd22008,17'd23040,17'd31829,17'd30427,17'd22331,17'd23217,17'd30128,17'd30579,17'd29829,17'd23388,17'd23569,17'd22501,17'd22328,17'd22325,17'd22505,17'd22334,17'd22683,17'd22683,17'd35292,17'd22159,17'd22159,17'd22506,17'd22856,17'd22330,17'd22503,17'd22501,17'd36543,17'd50732,17'd39440,17'd36543,17'd30277,17'd51229,17'd60479,17'd60241,17'd59859,17'd52668,17'd60480,17'd56973,17'd30424,17'd24902,17'd34884,17'd28595,17'd27637,17'd29103,17'd27511,17'd25317,17'd27765,17'd25567,17'd28594,17'd28720,17'd28723,17'd25566,17'd28723,17'd27765,17'd27882,17'd27882,17'd27882,17'd30903,17'd59999,17'd59213,17'd60114,17'd60117,17'd60481,17'd30148,17'd41119,17'd60482,17'd60483,17'd60484,17'd60485,17'd60486,17'd45162,17'd41584,17'd53494,17'd60487,17'd47163,17'd31345,17'd60488,17'd60489,17'd60490,17'd25039,17'd23058,17'd60491,17'd60492,17'd60493,17'd60494,17'd60495,17'd60496,17'd43449,17'd60497,17'd60498,17'd60499,17'd33685,17'd20513,17'd21278,17'd21894,17'd60500,17'd22395,17'd60501,17'd24792,17'd24643,17'd24306,17'd23277,17'd24644,17'd24650,17'd6546,17'd4993,17'd5325,17'd6067,17'd5145,17'd33838,17'd33838,17'd33841,17'd5155,17'd4687,17'd5002,17'd5335,17'd27935,17'd5160,17'd5004,17'd29024,17'd4685,17'd4841,17'd4684,17'd4370,17'd37808,17'd4380,17'd5488,17'd60502,17'd5925,17'd6568,17'd7844,17'd49709,17'd49709,17'd60392,17'd3545,17'd60503,17'd60504,17'd60393,17'd59484,17'd3543,17'd50285,17'd36446,17'd36446,17'd58357,17'd60505,17'd58851,17'd36449,17'd60506,17'd36742,17'd52837,17'd58982,17'd45182,17'd58489,17'd60507,17'd60508,17'd58858,17'd59485,17'd60394,17'd59760,17'd60271,17'd60145,17'd58241,17'd53740,17'd60509,17'd58748,17'd60510,17'd60511,17'd56550,17'd60512,17'd52363,17'd2587,17'd623,17'd625,17'd1680,17'd3743,17'd2409,17'd2589,17'd415,17'd421,17'd2763,17'd422,17'd603,17'd1272,17'd1537,17'd598,17'd777,17'd26228,17'd27707,17'd29610,17'd31251,17'd31251,17'd36905,17'd38719,17'd9124,17'd7538,17'd35769,17'd37445,17'd58991,17'd4867,17'd38072,17'd39033,17'd48559,17'd7191,17'd3218,17'd60513,17'd60514,17'd60515,17'd52458,17'd60402,17'd60403,17'd58621,17'd60516,17'd58874,17'd2071,17'd60517,17'd54320,17'd54082
},
'{
17'd3429,17'd3429,17'd3752,17'd3752,17'd2426,17'd2258,17'd1414,17'd1416,17'd19,17'd19,17'd10,17'd808,17'd10,17'd1128,17'd18,17'd19,17'd18,17'd3905,17'd1416,17'd1416,17'd4247,17'd1688,17'd2422,17'd2935,17'd2934,17'd35619,17'd60518,17'd10924,17'd10670,17'd10268,17'd291,17'd809,17'd22965,17'd2258,17'd3751,17'd4893,17'd15117,17'd15117,17'd58016,17'd14320,17'd15362,17'd60519,17'd60037,17'd59001,17'd60520,17'd844,17'd60040,17'd57372,17'd1430,17'd1430,17'd59500,17'd59500,17'd57006,17'd1562,17'd77,17'd60521,17'd73,17'd308,17'd670,17'd60522,17'd60523,17'd60524,17'd60525,17'd18396,17'd59006,17'd60409,17'd60526,17'd60527,17'd60528,17'd3938,17'd59510,17'd5996,17'd60529,17'd4463,17'd3139,17'd2825,17'd53611,17'd54901,17'd60530,17'd60531,17'd53689,17'd60532,17'd60416,17'd60294,17'd60533,17'd60294,17'd2654,17'd60534,17'd60535,17'd60296,17'd60420,17'd60536,17'd60537,17'd60538,17'd54802,17'd56580,17'd60539,17'd55092,17'd60540,17'd56582,17'd55378,17'd58885,17'd56583,17'd60303,17'd56811,17'd58661,17'd60541,17'd59522,17'd60542,17'd59647,17'd60543,17'd60544,17'd59144,17'd59024,17'd58157,17'd60545,17'd60309,17'd55681,17'd59941,17'd60546,17'd60547,17'd60313,17'd60548,17'd3507,17'd60549,17'd60550,17'd60551,17'd60552,17'd60553,17'd60554,17'd60555,17'd53528,17'd40875,17'd60556,17'd60557,17'd60558,17'd60559,17'd59039,17'd60560,17'd59954,17'd60446,17'd60328,17'd60561,17'd60562,17'd60563,17'd60449,17'd60564,17'd60450,17'd60565,17'd60566,17'd60452,17'd60332,17'd60567,17'd60568,17'd60456,17'd60569,17'd60570,17'd60571,17'd60572,17'd60573,17'd60339,17'd60574,17'd60341,17'd60216,17'd60343,17'd60575,17'd60576,17'd58685,17'd13346,17'd57808,17'd15041,17'd60577,17'd54730,17'd57314,17'd38238,17'd28233,17'd18448,17'd38910,17'd55942,17'd60578,17'd31135,17'd59839,17'd30681,17'd30680,17'd29647,17'd29647,17'd29647,17'd29482,17'd30373,17'd30373,17'd29481,17'd36347,17'd28572,17'd28348,17'd27234,17'd24991,17'd12254,17'd16203,17'd14130,17'd14261,17'd11807,17'd16069,17'd17236,17'd11400,17'd10479,17'd12116,17'd9620,17'd9344,17'd9342,17'd13887,17'd8873,17'd9195,17'd8576,17'd8419,17'd9889,17'd16689,17'd8258,17'd19924,17'd17856,17'd59842,17'd55829,17'd59706,17'd60349,17'd11969,17'd14681,17'd17241,17'd8580,17'd24213,17'd8412,17'd10027,17'd50864,17'd15429,17'd34829,17'd60579,17'd60580,17'd60581,17'd60582,17'd60583,17'd60584,17'd60585,17'd60586,17'd60587,17'd60588,17'd60357,17'd60589,17'd50064,17'd60590,17'd57073,17'd49472,17'd60478,17'd51653,17'd46753,17'd49273,17'd43286,17'd50264,17'd50157,17'd55847,17'd60591,17'd53720,17'd34276,17'd30127,17'd41273,17'd22334,17'd22008,17'd23040,17'd37385,17'd37510,17'd22856,17'd23389,17'd32191,17'd29829,17'd32008,17'd23217,17'd23218,17'd36986,17'd22678,17'd22332,17'd22333,17'd22160,17'd35292,17'd22507,17'd22683,17'd22160,17'd22506,17'd22332,17'd22680,17'd36986,17'd22328,17'd33158,17'd33158,17'd37116,17'd37116,17'd30277,17'd30277,17'd45746,17'd60592,17'd52965,17'd59337,17'd52815,17'd57455,17'd30578,17'd24086,17'd28852,17'd24252,17'd34283,17'd25177,17'd28850,17'd28369,17'd25567,17'd25567,17'd27638,17'd28720,17'd28723,17'd25566,17'd25566,17'd28600,17'd28369,17'd25709,17'd27882,17'd30903,17'd29256,17'd30292,17'd60593,17'd36267,17'd31361,17'd60594,17'd60595,17'd60595,17'd36135,17'd39751,17'd60596,17'd60597,17'd60598,17'd23221,17'd60599,17'd47250,17'd60600,17'd48164,17'd23926,17'd60601,17'd60602,17'd60603,17'd22699,17'd60604,17'd60376,17'd60605,17'd60606,17'd60607,17'd60608,17'd60609,17'd60610,17'd60611,17'd60612,17'd60613,17'd58842,17'd59107,17'd20977,17'd60614,17'd60615,17'd22567,17'd54496,17'd24792,17'd22934,17'd24306,17'd23108,17'd23110,17'd5147,17'd5148,17'd4993,17'd5325,17'd6067,17'd5145,17'd4189,17'd41891,17'd5154,17'd40397,17'd5002,17'd5004,17'd28185,17'd5614,17'd25627,17'd30637,17'd29024,17'd37433,17'd5328,17'd49995,17'd55869,17'd60616,17'd5622,17'd60617,17'd60618,17'd5925,17'd6862,17'd7844,17'd49709,17'd49709,17'd60392,17'd3545,17'd60503,17'd60619,17'd59484,17'd36317,17'd3543,17'd49004,17'd58733,17'd58484,17'd60505,17'd60505,17'd50285,17'd3542,17'd52187,17'd36742,17'd52837,17'd44738,17'd57996,17'd42192,17'd60507,17'd53431,17'd58619,17'd59485,17'd59760,17'd59760,17'd60271,17'd53667,17'd57233,17'd60620,17'd60621,17'd59904,17'd60622,17'd60623,17'd60624,17'd58129,17'd629,17'd1402,17'd446,17'd1261,17'd5050,17'd11337,17'd413,17'd1383,17'd415,17'd1529,17'd2763,17'd422,17'd598,17'd1272,17'd424,17'd2589,17'd1949,17'd26228,17'd27707,17'd29610,17'd60625,17'd60625,17'd36905,17'd60626,17'd7538,17'd7538,17'd6417,17'd60627,17'd38459,17'd13420,17'd44019,17'd38859,17'd39179,17'd5932,17'd60628,17'd20861,17'd60629,17'd60630,17'd60631,17'd37041,17'd60632,17'd58621,17'd60516,17'd58874,17'd2071,17'd60517,17'd54320,17'd54082
},
'{
17'd52621,17'd3429,17'd3752,17'd3752,17'd2258,17'd2258,17'd2257,17'd1416,17'd13,17'd12,17'd10,17'd808,17'd10,17'd1128,17'd19,17'd979,17'd18,17'd18,17'd3905,17'd17,17'd1414,17'd2597,17'd2422,17'd2784,17'd2934,17'd3428,17'd35619,17'd15358,17'd10670,17'd3429,17'd2597,17'd2257,17'd22965,17'd2258,17'd2593,17'd4086,17'd15117,17'd14744,17'd5203,17'd14320,17'd1279,17'd815,17'd47,17'd60633,17'd60634,17'd60635,17'd57002,17'd57002,17'd60636,17'd56795,17'd56793,17'd60637,17'd20406,17'd674,17'd77,17'd492,17'd311,17'd1000,17'd485,17'd837,17'd60406,17'd60638,17'd21640,17'd2803,17'd60639,17'd60640,17'd60285,17'd60641,17'd60642,17'd60643,17'd60644,17'd5995,17'd6302,17'd4768,17'd3627,17'd5690,17'd53815,17'd60645,17'd60646,17'd60647,17'd60648,17'd5697,17'd60649,17'd60650,17'd60649,17'd60649,17'd60651,17'd2655,17'd4296,17'd59784,17'd3304,17'd60652,17'd60653,17'd60654,17'd60300,17'd60655,17'd60656,17'd55282,17'd55674,17'd56236,17'd60657,17'd57647,17'd59523,17'd57917,17'd60658,17'd60659,17'd56811,17'd58769,17'd60660,17'd58769,17'd60658,17'd60661,17'd60662,17'd60427,17'd60663,17'd60664,17'd60665,17'd55587,17'd60666,17'd60667,17'd58665,17'd59404,17'd60668,17'd60669,17'd60670,17'd60671,17'd60672,17'd60673,17'd60674,17'd60675,17'd60676,17'd60677,17'd60678,17'd38350,17'd60679,17'd60680,17'd57933,17'd58424,17'd59298,17'd60681,17'd60682,17'd60683,17'd60684,17'd60685,17'd60686,17'd59956,17'd60687,17'd60450,17'd60451,17'd60688,17'd60689,17'd60690,17'd60567,17'd60691,17'd60692,17'd60693,17'd60694,17'd60695,17'd60696,17'd60697,17'd60698,17'd60086,17'd60699,17'd60700,17'd60701,17'd60702,17'd59430,17'd60703,17'd59316,17'd58443,17'd60704,17'd15671,17'd54822,17'd54374,17'd38238,17'd37738,17'd18448,17'd18448,17'd39825,17'd57817,17'd30977,17'd58077,17'd58312,17'd58312,17'd29786,17'd29648,17'd29481,17'd29481,17'd36347,17'd28345,17'd28818,17'd28460,17'd27858,17'd26758,17'd18200,17'd12254,17'd12579,17'd11959,17'd13135,17'd11807,17'd16069,17'd17236,17'd12863,17'd9884,17'd9620,17'd9339,17'd9189,17'd9038,17'd9193,17'd29063,17'd8877,17'd8731,17'd60705,17'd15056,17'd56166,17'd15813,17'd21059,17'd15575,17'd19650,17'd60706,17'd60707,17'd60100,17'd60708,17'd60709,17'd7789,17'd7949,17'd10028,17'd25147,17'd11966,17'd8878,17'd8725,17'd8413,17'd60710,17'd57692,17'd60580,17'd53111,17'd60711,17'd60712,17'd60713,17'd60714,17'd60715,17'd60716,17'd60717,17'd60718,17'd49373,17'd60477,17'd60590,17'd47923,17'd49473,17'd46662,17'd51746,17'd43979,17'd49273,17'd45036,17'd54205,17'd60719,17'd53986,17'd60591,17'd53557,17'd38808,17'd29099,17'd36426,17'd22159,17'd22861,17'd23040,17'd32345,17'd37659,17'd36009,17'd39131,17'd23218,17'd22501,17'd33158,17'd37533,17'd30729,17'd35017,17'd35736,17'd40052,17'd22158,17'd22507,17'd22683,17'd35292,17'd35292,17'd22160,17'd22333,17'd22856,17'd22330,17'd22329,17'd22501,17'd22501,17'd36543,17'd51229,17'd22328,17'd32827,17'd45616,17'd60720,17'd52965,17'd52965,17'd57077,17'd56751,17'd40680,17'd23733,17'd24902,17'd29100,17'd28718,17'd25320,17'd25438,17'd27511,17'd28369,17'd25567,17'd25567,17'd28594,17'd28723,17'd28723,17'd25566,17'd28721,17'd28600,17'd27882,17'd25438,17'd27511,17'd33345,17'd32040,17'd25952,17'd59993,17'd60721,17'd60722,17'd60723,17'd60724,17'd60725,17'd60726,17'd60727,17'd32851,17'd60728,17'd60729,17'd50478,17'd60730,17'd60731,17'd60732,17'd60733,17'd31663,17'd60734,17'd60735,17'd36863,17'd60736,17'd60737,17'd25974,17'd60738,17'd60739,17'd60740,17'd60741,17'd60742,17'd60743,17'd60744,17'd60745,17'd60746,17'd60747,17'd21278,17'd60748,17'd60749,17'd23100,17'd23620,17'd54593,17'd24792,17'd30793,17'd22933,17'd23278,17'd23110,17'd6546,17'd5150,17'd5325,17'd5324,17'd4682,17'd5145,17'd41891,17'd4998,17'd5154,17'd4847,17'd5005,17'd5335,17'd5614,17'd28185,17'd30637,17'd53578,17'd37433,17'd40397,17'd4847,17'd38568,17'd56203,17'd6072,17'd60750,17'd60751,17'd5925,17'd60752,17'd7188,17'd19858,17'd49403,17'd49403,17'd3545,17'd60753,17'd21010,17'd60754,17'd60754,17'd60619,17'd3543,17'd3543,17'd60755,17'd60756,17'd58357,17'd60505,17'd50285,17'd59233,17'd59614,17'd52767,17'd60757,17'd41309,17'd42040,17'd42040,17'd60758,17'd60759,17'd60508,17'd60760,17'd60761,17'd59760,17'd60144,17'd57742,17'd60027,17'd60509,17'd60762,17'd60763,17'd60764,17'd60765,17'd60766,17'd60767,17'd2587,17'd231,17'd1263,17'd1261,17'd5957,17'd6868,17'd2589,17'd1383,17'd194,17'd1529,17'd1529,17'd1529,17'd1669,17'd202,17'd598,17'd413,17'd1949,17'd28429,17'd27708,17'd29170,17'd31251,17'd36905,17'd35487,17'd33051,17'd7538,17'd7538,17'd60768,17'd37445,17'd48187,17'd14177,17'd38334,17'd5355,17'd3871,17'd40715,17'd60513,17'd60769,17'd60770,17'd60630,17'd51493,17'd36900,17'd60771,17'd58621,17'd60772,17'd54159,17'd2071,17'd24320,17'd54320,17'd60035
},
'{
17'd52621,17'd3429,17'd3752,17'd3752,17'd2258,17'd2258,17'd2257,17'd1414,17'd2,17'd12,17'd10,17'd808,17'd10,17'd1128,17'd18,17'd979,17'd18,17'd18,17'd18,17'd17,17'd1414,17'd2597,17'd2422,17'd2784,17'd2934,17'd3428,17'd35619,17'd35619,17'd10670,17'd10669,17'd3752,17'd2597,17'd2257,17'd2258,17'd2935,17'd3592,17'd5203,17'd5203,17'd5511,17'd5204,17'd58016,17'd15497,17'd60773,17'd60774,17'd60039,17'd60281,17'd56672,17'd56892,17'd56438,17'd56795,17'd56793,17'd60775,17'd60776,17'd20406,17'd312,17'd492,17'd20406,17'd1000,17'd305,17'd18151,17'd2794,17'd60523,17'd60524,17'd2451,17'd60777,17'd60778,17'd60779,17'd60157,17'd60780,17'd60781,17'd60782,17'd5684,17'd31269,17'd5835,17'd60783,17'd3470,17'd60784,17'd60531,17'd60785,17'd60785,17'd60786,17'd60787,17'd60788,17'd60650,17'd53759,17'd60649,17'd53759,17'd60650,17'd2655,17'd4296,17'd59514,17'd60420,17'd60536,17'd60789,17'd60790,17'd56910,17'd57019,17'd58652,17'd57277,17'd55671,17'd56128,17'd58159,17'd58885,17'd59933,17'd60791,17'd60792,17'd60793,17'd60794,17'd60795,17'd60795,17'd59147,17'd60661,17'd60796,17'd60308,17'd60183,17'd60183,17'd60797,17'd60798,17'd59940,17'd57023,17'd60799,17'd60800,17'd60668,17'd1189,17'd3808,17'd60801,17'd60802,17'd60803,17'd60804,17'd60805,17'd60806,17'd60807,17'd60808,17'd60809,17'd60810,17'd60811,17'd60812,17'd60813,17'd59298,17'd60681,17'd60814,17'd60561,17'd60815,17'd60816,17'd60817,17'd59956,17'd60818,17'd60687,17'd60450,17'd60451,17'd60688,17'd60689,17'd60207,17'd60691,17'd60819,17'd60820,17'd60821,17'd60822,17'd60823,17'd60824,17'd60825,17'd60215,17'd59828,17'd60699,17'd59689,17'd59690,17'd60343,17'd60826,17'd59833,17'd60827,17'd57680,17'd13875,17'd60828,17'd56495,17'd54825,17'd37738,17'd18685,17'd17724,17'd18448,17'd30978,17'd31135,17'd31135,17'd58806,17'd58693,17'd29648,17'd31134,17'd29481,17'd50213,17'd28818,17'd28229,17'd27857,17'd28104,17'd26758,17'd18084,17'd18564,17'd16203,17'd11959,17'd13520,17'd11807,17'd16068,17'd11524,17'd11526,17'd10169,17'd10025,17'd10173,17'd17480,17'd9194,17'd9040,17'd8721,17'd8876,17'd23517,17'd50524,17'd8888,17'd25152,17'd60829,17'd12727,17'd21366,17'd15950,17'd56276,17'd22828,17'd60830,17'd60100,17'd54649,17'd9624,17'd10180,17'd17354,17'd17240,17'd25147,17'd11966,17'd8724,17'd10607,17'd21987,17'd25680,17'd60831,17'd51882,17'd24717,17'd60832,17'd60833,17'd60834,17'd60835,17'd60836,17'd60837,17'd60475,17'd60718,17'd60838,17'd60590,17'd60839,17'd55840,17'd54939,17'd50158,17'd51746,17'd43979,17'd47727,17'd43285,17'd60840,17'd60841,17'd51554,17'd60842,17'd53193,17'd34276,17'd29099,17'd36426,17'd22160,17'd35153,17'd23040,17'd32345,17'd31496,17'd30427,17'd39131,17'd23389,17'd30277,17'd22328,17'd32015,17'd35017,17'd35158,17'd44360,17'd35296,17'd30426,17'd22158,17'd22161,17'd22159,17'd22159,17'd22506,17'd22332,17'd22680,17'd36986,17'd30277,17'd22501,17'd22501,17'd33158,17'd22503,17'd36986,17'd36986,17'd51229,17'd60843,17'd59720,17'd39280,17'd46427,17'd40680,17'd23734,17'd23384,17'd29102,17'd28601,17'd24745,17'd29244,17'd27511,17'd28369,17'd28369,17'd25567,17'd27765,17'd28720,17'd28723,17'd25566,17'd28723,17'd28600,17'd25317,17'd27511,17'd25438,17'd29103,17'd33345,17'd25952,17'd30445,17'd33019,17'd60844,17'd33181,17'd60845,17'd30291,17'd35433,17'd60846,17'd60847,17'd60848,17'd60849,17'd60850,17'd60851,17'd60852,17'd60853,17'd60854,17'd48712,17'd60855,17'd60856,17'd60857,17'd60858,17'd60859,17'd60860,17'd60861,17'd60862,17'd60863,17'd20197,17'd60864,17'd60865,17'd60866,17'd60867,17'd60868,17'd20820,17'd60869,17'd20977,17'd60870,17'd60871,17'd60872,17'd56875,17'd54593,17'd24643,17'd24305,17'd22933,17'd23109,17'd6543,17'd5325,17'd5480,17'd5325,17'd5324,17'd6067,17'd5144,17'd33992,17'd34657,17'd34791,17'd29024,17'd5004,17'd5335,17'd27935,17'd30638,17'd30180,17'd28536,17'd40397,17'd40397,17'd4527,17'd60873,17'd60874,17'd7334,17'd60875,17'd60751,17'd5925,17'd60752,17'd6717,17'd21619,17'd6568,17'd7508,17'd3545,17'd60753,17'd60267,17'd60754,17'd60754,17'd60619,17'd3543,17'd3543,17'd60756,17'd60756,17'd60756,17'd58851,17'd36893,17'd60876,17'd59896,17'd48182,17'd45652,17'd60877,17'd60878,17'd60507,17'd22602,17'd60758,17'd42328,17'd42328,17'd60760,17'd60879,17'd60880,17'd60881,17'd60882,17'd60509,17'd60883,17'd56554,17'd60884,17'd60885,17'd52534,17'd30342,17'd623,17'd1399,17'd1401,17'd5050,17'd6868,17'd2409,17'd2589,17'd1383,17'd194,17'd1529,17'd1529,17'd415,17'd421,17'd1526,17'd414,17'd15233,17'd26228,17'd28429,17'd27708,17'd31251,17'd60030,17'd36905,17'd33051,17'd9124,17'd7538,17'd60886,17'd36045,17'd60887,17'd16855,17'd13572,17'd38202,17'd47767,17'd3871,17'd40562,17'd60513,17'd60888,17'd60889,17'd60890,17'd56214,17'd37165,17'd2360,17'd58621,17'd60772,17'd58874,17'd58999,17'd24320,17'd54320,17'd54082
},
'{
17'd52621,17'd3429,17'd3752,17'd3752,17'd3429,17'd2426,17'd4247,17'd466,17'd12,17'd12,17'd10,17'd808,17'd10,17'd11,17'd18,17'd19,17'd652,17'd652,17'd18,17'd3905,17'd1416,17'd2257,17'd1831,17'd2422,17'd3101,17'd3428,17'd35619,17'd35619,17'd54978,17'd10669,17'd3752,17'd2597,17'd2257,17'd2597,17'd10669,17'd10925,17'd5204,17'd5203,17'd5511,17'd5204,17'd12504,17'd14599,17'd60891,17'd58255,17'd59499,17'd60634,17'd56891,17'd56438,17'd57003,17'd57003,17'd20272,17'd60775,17'd60892,17'd60893,17'd311,17'd491,17'd840,17'd56794,17'd68,17'd60894,17'd60895,17'd60896,17'd60897,17'd3274,17'd60898,17'd58389,17'd60899,17'd60900,17'd60901,17'd59922,17'd60902,17'd60412,17'd5833,17'd60289,17'd60903,17'd6477,17'd60904,17'd60905,17'd60906,17'd60785,17'd60907,17'd60908,17'd60909,17'd60784,17'd60784,17'd6008,17'd53526,17'd60910,17'd60651,17'd2826,17'd59929,17'd3636,17'd60911,17'd60912,17'd60913,17'd60914,17'd60915,17'd58408,17'd60916,17'd60917,17'd60918,17'd60919,17'd58772,17'd59523,17'd58279,17'd60920,17'd60792,17'd59399,17'd59282,17'd1320,17'd59282,17'd60921,17'd59277,17'd60922,17'd60545,17'd60923,17'd57022,17'd60924,17'd59657,17'd60925,17'd60926,17'd60927,17'd1038,17'd60928,17'd60929,17'd60930,17'd60931,17'd60932,17'd60933,17'd60934,17'd60935,17'd60936,17'd60937,17'd60938,17'd60939,17'd60940,17'd60941,17'd60942,17'd60943,17'd60944,17'd60945,17'd60446,17'd60815,17'd60946,17'd60817,17'd60947,17'd60563,17'd60449,17'd60564,17'd60450,17'd60948,17'd60949,17'd60950,17'd60951,17'd60952,17'd60691,17'd60953,17'd60954,17'd60955,17'd60956,17'd60957,17'd60958,17'd60959,17'd60960,17'd60961,17'd59966,17'd60962,17'd59430,17'd60963,17'd59318,17'd60964,17'd60965,17'd54557,17'd60966,17'd53900,17'd17725,17'd17724,17'd17724,17'd18448,17'd31772,17'd30978,17'd59064,17'd30976,17'd31771,17'd31771,17'd30976,17'd50213,17'd29336,17'd27857,17'd27858,17'd26872,17'd25927,17'd24207,17'd28950,17'd15184,17'd19920,17'd15185,17'd11395,17'd14810,17'd13001,17'd10330,17'd10169,17'd9340,17'd10335,17'd17123,17'd29920,17'd9046,17'd8724,17'd8567,17'd8568,17'd8575,17'd60967,17'd16333,17'd24216,17'd60968,17'd10747,17'd18809,17'd15061,17'd60969,17'd60970,17'd60971,17'd60972,17'd10182,17'd18205,17'd14680,17'd9622,17'd8250,17'd8578,17'd8572,17'd12425,17'd8571,17'd9196,17'd17352,17'd60973,17'd59846,17'd60974,17'd60832,17'd60975,17'd60976,17'd60977,17'd60978,17'd60979,17'd60980,17'd60981,17'd60982,17'd60983,17'd60984,17'd55840,17'd47530,17'd57713,17'd51746,17'd43979,17'd47629,17'd54480,17'd60985,17'd60986,17'd60987,17'd57325,17'd53193,17'd34276,17'd29099,17'd30425,17'd22506,17'd22507,17'd32497,17'd30580,17'd32660,17'd32344,17'd22678,17'd36986,17'd36986,17'd22330,17'd44702,17'd34278,17'd40523,17'd33645,17'd46958,17'd33944,17'd32344,17'd22159,17'd22159,17'd22506,17'd22333,17'd30276,17'd22331,17'd22329,17'd30277,17'd22501,17'd22503,17'd22328,17'd22330,17'd22331,17'd22327,17'd39912,17'd39744,17'd45746,17'd51552,17'd38980,17'd23734,17'd23565,17'd29378,17'd28852,17'd24744,17'd29976,17'd29103,17'd27511,17'd28369,17'd28369,17'd27765,17'd28130,17'd28723,17'd25566,17'd25566,17'd28720,17'd27765,17'd27882,17'd34127,17'd60988,17'd60989,17'd60990,17'd60362,17'd36549,17'd60721,17'd60482,17'd60845,17'd37405,17'd60991,17'd38038,17'd34888,17'd60992,17'd60993,17'd43438,17'd60994,17'd60995,17'd60996,17'd60997,17'd60998,17'd60999,17'd61000,17'd61001,17'd61002,17'd61003,17'd31686,17'd61004,17'd61005,17'd61006,17'd61007,17'd61008,17'd61009,17'd39763,17'd26208,17'd20363,17'd61010,17'd21118,17'd61011,17'd61012,17'd61013,17'd22225,17'd22394,17'd23792,17'd24305,17'd24643,17'd24305,17'd22933,17'd25222,17'd7658,17'd5325,17'd4841,17'd4683,17'd4683,17'd6067,17'd38442,17'd33992,17'd33841,17'd5156,17'd5157,17'd5329,17'd5335,17'd28185,17'd31553,17'd37288,17'd37433,17'd49995,17'd58971,17'd50587,17'd52997,17'd61014,17'd9096,17'd10785,17'd5174,17'd8945,17'd61015,17'd4212,17'd61016,17'd7188,17'd7845,17'd61017,17'd3691,17'd60504,17'd59233,17'd59232,17'd3543,17'd49004,17'd49004,17'd49004,17'd58732,17'd58732,17'd61018,17'd59233,17'd60876,17'd36742,17'd3365,17'd61019,17'd61020,17'd60507,17'd53431,17'd61021,17'd58737,17'd60270,17'd58858,17'd60394,17'd61022,17'd61023,17'd56000,17'd54972,17'd61024,17'd61025,17'd55888,17'd53595,17'd61026,17'd1378,17'd20270,17'd626,17'd230,17'd3743,17'd5371,17'd6868,17'd2409,17'd413,17'd779,17'd1671,17'd776,17'd776,17'd776,17'd941,17'd940,17'd15233,17'd28916,17'd28429,17'd61027,17'd27708,17'd31251,17'd36903,17'd35487,17'd9124,17'd7538,17'd7538,17'd60886,17'd6417,17'd16492,17'd14177,17'd44019,17'd61028,17'd47767,17'd40099,17'd40861,17'd61029,17'd61030,17'd61031,17'd50753,17'd56427,17'd61032,17'd32556,17'd2069,17'd60516,17'd60516,17'd58999,17'd61033,17'd61034,17'd54082
},
'{
17'd52621,17'd3429,17'd3752,17'd3429,17'd52621,17'd52621,17'd1831,17'd4247,17'd0,17'd12,17'd10,17'd808,17'd808,17'd11,17'd18,17'd19,17'd652,17'd652,17'd18,17'd17,17'd1414,17'd2596,17'd3250,17'd2784,17'd2934,17'd3428,17'd35619,17'd35619,17'd59496,17'd10802,17'd3429,17'd3752,17'd2597,17'd2597,17'd3429,17'd10924,17'd5204,17'd5511,17'd5511,17'd5511,17'd12653,17'd14989,17'd59497,17'd59775,17'd61035,17'd59499,17'd56891,17'd56792,17'd56892,17'd56892,17'd56795,17'd20272,17'd61036,17'd60892,17'd56796,17'd841,17'd1150,17'd56795,17'd55892,17'd61037,17'd60895,17'd61038,17'd61039,17'd61040,17'd20013,17'd61041,17'd61042,17'd61043,17'd61044,17'd59780,17'd61045,17'd60782,17'd59510,17'd5834,17'd61046,17'd61047,17'd6317,17'd6008,17'd61048,17'd61049,17'd60906,17'd61050,17'd61051,17'd61052,17'd61053,17'd6008,17'd61054,17'd60910,17'd61055,17'd2657,17'd4929,17'd3143,17'd2644,17'd2296,17'd61056,17'd61057,17'd60915,17'd61058,17'd59517,17'd61059,17'd61060,17'd56030,17'd57278,17'd58160,17'd58888,17'd60055,17'd60920,17'd60793,17'd57649,17'd60795,17'd57644,17'd59147,17'd61061,17'd61062,17'd61063,17'd59938,17'd59792,17'd61064,17'd59797,17'd61065,17'd57023,17'd61066,17'd61067,17'd60668,17'd61068,17'd2328,17'd61069,17'd61070,17'd61071,17'd61072,17'd60553,17'd61073,17'd61074,17'd61075,17'd61076,17'd61077,17'd61078,17'd61079,17'd61080,17'd61081,17'd60944,17'd60814,17'd61082,17'd61083,17'd60817,17'd61084,17'd60563,17'd61085,17'd61086,17'd60564,17'd61087,17'd60948,17'd61088,17'd61089,17'd61090,17'd60951,17'd61091,17'd61092,17'd60955,17'd60956,17'd61093,17'd60825,17'd61094,17'd61095,17'd60959,17'd59828,17'd60341,17'd60702,17'd61096,17'd59314,17'd60221,17'd61097,17'd61098,17'd54559,17'd53706,17'd54825,17'd17013,17'd17013,17'd17724,17'd18448,17'd39661,17'd39661,17'd31136,17'd30976,17'd30976,17'd28572,17'd28572,17'd27857,17'd27737,17'd27123,17'd25927,17'd24707,17'd16324,17'd15055,17'd19920,17'd15185,17'd11395,17'd14810,17'd13886,17'd11527,17'd10169,17'd17965,17'd14674,17'd16795,17'd29920,17'd12425,17'd8571,17'd8571,17'd8569,17'd10607,17'd61099,17'd52404,17'd15440,17'd60968,17'd22995,17'd24869,17'd14387,17'd24370,17'd8430,17'd22303,17'd61100,17'd61101,17'd21367,17'd18205,17'd7790,17'd9622,17'd8250,17'd37734,17'd24711,17'd8731,17'd8573,17'd8578,17'd25411,17'd61102,17'd61103,17'd61104,17'd61105,17'd61106,17'd61107,17'd61108,17'd61109,17'd61110,17'd61111,17'd60981,17'd49781,17'd61112,17'd61113,17'd48033,17'd50994,17'd50070,17'd42299,17'd44106,17'd44230,17'd61114,17'd61115,17'd61116,17'd58710,17'd50646,17'd53193,17'd28368,17'd29376,17'd30425,17'd22333,17'd22162,17'd30580,17'd32660,17'd22161,17'd22333,17'd22331,17'd36986,17'd22680,17'd22678,17'd44591,17'd34278,17'd40523,17'd40523,17'd23926,17'd39441,17'd22333,17'd22506,17'd22506,17'd22677,17'd22856,17'd22331,17'd22329,17'd22328,17'd30277,17'd22501,17'd22503,17'd22329,17'd22680,17'd22331,17'd45874,17'd53781,17'd45874,17'd39588,17'd39280,17'd38806,17'd29376,17'd29972,17'd23563,17'd24742,17'd29976,17'd29103,17'd27511,17'd28850,17'd28369,17'd28369,17'd27765,17'd28600,17'd25566,17'd25566,17'd25566,17'd28130,17'd28369,17'd34127,17'd60988,17'd33345,17'd60989,17'd59213,17'd36549,17'd36135,17'd35859,17'd61117,17'd35714,17'd61118,17'd33808,17'd29264,17'd33957,17'd34889,17'd61119,17'd61120,17'd46335,17'd61121,17'd61122,17'd61123,17'd61124,17'd41121,17'd61125,17'd61126,17'd61127,17'd61128,17'd61129,17'd61130,17'd61131,17'd61132,17'd30911,17'd61133,17'd61134,17'd61135,17'd26102,17'd27925,17'd17742,17'd61136,17'd61137,17'd61138,17'd61139,17'd22927,17'd23445,17'd24305,17'd25222,17'd23109,17'd24305,17'd24643,17'd24794,17'd7325,17'd4993,17'd4841,17'd4683,17'd4683,17'd5145,17'd33532,17'd4998,17'd5155,17'd4846,17'd5162,17'd5160,17'd5335,17'd30638,17'd32553,17'd61140,17'd37433,17'd49995,17'd49896,17'd61141,17'd37033,17'd8160,17'd22769,17'd61142,17'd5020,17'd8944,17'd61015,17'd4701,17'd61143,17'd4041,17'd61144,17'd49601,17'd61145,17'd60504,17'd36449,17'd59232,17'd3543,17'd49004,17'd49004,17'd49004,17'd58732,17'd61018,17'd53142,17'd53142,17'd52607,17'd61146,17'd3193,17'd60877,17'd61147,17'd61148,17'd61149,17'd61021,17'd53431,17'd58738,17'd58984,17'd57357,17'd61150,17'd61151,17'd61152,17'd59903,17'd61153,17'd57755,17'd61154,17'd61155,17'd61156,17'd1090,17'd772,17'd1262,17'd1401,17'd4880,17'd5372,17'd2409,17'd412,17'd413,17'd779,17'd1671,17'd776,17'd776,17'd776,17'd776,17'd776,17'd27094,17'd29037,17'd28429,17'd29441,17'd31251,17'd31251,17'd36903,17'd35487,17'd9124,17'd61157,17'd60886,17'd61158,17'd39791,17'd16132,17'd14584,17'd38580,17'd40101,17'd47767,17'd4225,17'd50001,17'd61159,17'd61160,17'd54974,17'd53744,17'd61161,17'd61162,17'd61163,17'd56544,17'd2071,17'd60772,17'd61164,17'd61165,17'd54320,17'd54082
},
'{
17'd52621,17'd3429,17'd10546,17'd3593,17'd52621,17'd52621,17'd1831,17'd4247,17'd0,17'd12,17'd806,17'd465,17'd808,17'd11,17'd18,17'd18,17'd652,17'd652,17'd18,17'd3905,17'd17,17'd1414,17'd1688,17'd3250,17'd2935,17'd3427,17'd35619,17'd60150,17'd59496,17'd10670,17'd52621,17'd3752,17'd1129,17'd1129,17'd2597,17'd52621,17'd3428,17'd5511,17'd5511,17'd5511,17'd12504,17'd15118,17'd61166,17'd45,17'd59251,17'd59499,17'd56790,17'd56672,17'd57002,17'd56892,17'd1430,17'd20406,17'd310,17'd60892,17'd56796,17'd56795,17'd1150,17'd57005,17'd60892,17'd61167,17'd61168,17'd61169,17'd55086,17'd34349,17'd61170,17'd2452,17'd61171,17'd60156,17'd61172,17'd60780,17'd60781,17'd61173,17'd5405,17'd5543,17'd5685,17'd61174,17'd61175,17'd6000,17'd61176,17'd61177,17'd61178,17'd61179,17'd5707,17'd61180,17'd60784,17'd6008,17'd61054,17'd60533,17'd61181,17'd5546,17'd61182,17'd2990,17'd2465,17'd61183,17'd61184,17'd60913,17'd61185,17'd61186,17'd57275,17'd57275,17'd57642,17'd61187,17'd61188,17'd61189,17'd61190,17'd61191,17'd61192,17'd61193,17'd58661,17'd58769,17'd60427,17'd59401,17'd61194,17'd61195,17'd60658,17'd59279,17'd59024,17'd57022,17'd59276,17'd59151,17'd59026,17'd60667,17'd61196,17'd59800,17'd59527,17'd60928,17'd61197,17'd61198,17'd61199,17'd61200,17'd61201,17'd60437,17'd54811,17'd61202,17'd61203,17'd60322,17'd61204,17'd61205,17'd61206,17'd61207,17'd60944,17'd61208,17'd60685,17'd60685,17'd61209,17'd61210,17'd61211,17'd61212,17'd61085,17'd61086,17'd61213,17'd61214,17'd61215,17'd61216,17'd61217,17'd61089,17'd61218,17'd61219,17'd60955,17'd61220,17'd61221,17'd61222,17'd61223,17'd61224,17'd61225,17'd61226,17'd59966,17'd59555,17'd61227,17'd59431,17'd59182,17'd57808,17'd13497,17'd54729,17'd53468,17'd45209,17'd61228,17'd17235,17'd17726,17'd17726,17'd28233,17'd28349,17'd31136,17'd31136,17'd28945,17'd28350,17'd28348,17'd27737,17'd18083,17'd24207,17'd25671,17'd30229,17'd14261,17'd14379,17'd11522,17'd16068,17'd12720,17'd10605,17'd17720,17'd9740,17'd10743,17'd15187,17'd37605,17'd39660,17'd8724,17'd15429,17'd21987,17'd24710,17'd8730,17'd8575,17'd61229,17'd13765,17'd25004,17'd15572,17'd10747,17'd15691,17'd14387,17'd14817,17'd61230,17'd61231,17'd61232,17'd61233,17'd10483,17'd13528,17'd7618,17'd12120,17'd8250,17'd19923,17'd8571,17'd8571,17'd21987,17'd8733,17'd15056,17'd53979,17'd61234,17'd25296,17'd61235,17'd61236,17'd61237,17'd61238,17'd61239,17'd59714,17'd61240,17'd60981,17'd50064,17'd61241,17'd61113,17'd48033,17'd50994,17'd49978,17'd42597,17'd44230,17'd43285,17'd58953,17'd54837,17'd61242,17'd61243,17'd51233,17'd49080,17'd34106,17'd23565,17'd29973,17'd22332,17'd37510,17'd32660,17'd22158,17'd22334,17'd22504,17'd22500,17'd36986,17'd22680,17'd22677,17'd40523,17'd48913,17'd48913,17'd23391,17'd23391,17'd48913,17'd40523,17'd34107,17'd22332,17'd22678,17'd22331,17'd36986,17'd22328,17'd30277,17'd30277,17'd30277,17'd22328,17'd36986,17'd22680,17'd22331,17'd47457,17'd47457,17'd22327,17'd51229,17'd41587,17'd23923,17'd29529,17'd29532,17'd28601,17'd25031,17'd31034,17'd27511,17'd25438,17'd27511,17'd28369,17'd28369,17'd28130,17'd28721,17'd32658,17'd25566,17'd25435,17'd27765,17'd25835,17'd30903,17'd33345,17'd59213,17'd61244,17'd61245,17'd42006,17'd35859,17'd38161,17'd61246,17'd33326,17'd38166,17'd61247,17'd61248,17'd24102,17'd61249,17'd61250,17'd47166,17'd51005,17'd61251,17'd61252,17'd61253,17'd43162,17'd61254,17'd61255,17'd61256,17'd61257,17'd61258,17'd61259,17'd21719,17'd61260,17'd61261,17'd61262,17'd19303,17'd50280,17'd61263,17'd61264,17'd61265,17'd21743,17'd21584,17'd21284,17'd61266,17'd61267,17'd22928,17'd23106,17'd61268,17'd10881,17'd10881,17'd23109,17'd23109,17'd22759,17'd7163,17'd4993,17'd5328,17'd4683,17'd4682,17'd41891,17'd46979,17'd39470,17'd5155,17'd4846,17'd5162,17'd5166,17'd37030,17'd5165,17'd37288,17'd37433,17'd40397,17'd4690,17'd55457,17'd61269,17'd4540,17'd20700,17'd21936,17'd61270,17'd61271,17'd19857,17'd8944,17'd4701,17'd4213,17'd61272,17'd33045,17'd61017,17'd61273,17'd36449,17'd36448,17'd58483,17'd60756,17'd49004,17'd49004,17'd36317,17'd36317,17'd61274,17'd60506,17'd59755,17'd59369,17'd59759,17'd60877,17'd61275,17'd58616,17'd53286,17'd53286,17'd61148,17'd61148,17'd61276,17'd57357,17'd57742,17'd57099,17'd24662,17'd61277,17'd58874,17'd61278,17'd61279,17'd61280,17'd58862,17'd59766,17'd1959,17'd259,17'd1823,17'd3743,17'd5371,17'd6415,17'd412,17'd602,17'd1529,17'd415,17'd1671,17'd776,17'd29440,17'd29440,17'd33847,17'd33847,17'd29169,17'd29610,17'd27708,17'd29039,17'd31251,17'd29611,17'd58990,17'd11882,17'd7537,17'd8507,17'd6418,17'd36045,17'd60887,17'd16623,17'd13420,17'd38860,17'd40101,17'd10790,17'd53591,17'd50183,17'd61159,17'd41477,17'd61281,17'd41477,17'd51408,17'd61282,17'd61283,17'd2069,17'd60516,17'd61284,17'd61164,17'd60517,17'd54320,17'd60035
},
'{
17'd52621,17'd3429,17'd10546,17'd3593,17'd52621,17'd52621,17'd1831,17'd1688,17'd14,17'd0,17'd3,17'd465,17'd808,17'd10,17'd18,17'd18,17'd652,17'd652,17'd18,17'd16,17'd1415,17'd2596,17'd3250,17'd2592,17'd2782,17'd2934,17'd15358,17'd60150,17'd61285,17'd54978,17'd52621,17'd3429,17'd1129,17'd1129,17'd2597,17'd52621,17'd3427,17'd15496,17'd5511,17'd5203,17'd16392,17'd57896,17'd59381,17'd61286,17'd61287,17'd61035,17'd60280,17'd56891,17'd57002,17'd57372,17'd61288,17'd20406,17'd73,17'd60892,17'd55892,17'd56794,17'd56795,17'd20406,17'd75,17'd18039,17'd61168,17'd61289,17'd1709,17'd2620,17'd61290,17'd61291,17'd61292,17'd61293,17'd61294,17'd60044,17'd3456,17'd61295,17'd61296,17'd61297,17'd61298,17'd61299,17'd61300,17'd61301,17'd6144,17'd61302,17'd61049,17'd61303,17'd61304,17'd61051,17'd61052,17'd6008,17'd5697,17'd5698,17'd61055,17'd5546,17'd2651,17'd4130,17'd2990,17'd61183,17'd61305,17'd61306,17'd61307,17'd61308,17'd61309,17'd59523,17'd58885,17'd55783,17'd61310,17'd55091,17'd58525,17'd61311,17'd61312,17'd59795,17'd58894,17'd59276,17'd59273,17'd60660,17'd59520,17'd56584,17'd59653,17'd59648,17'd61313,17'd60428,17'd58769,17'd59797,17'd59657,17'd59026,17'd61314,17'd61315,17'd61316,17'd61317,17'd61318,17'd61319,17'd61320,17'd61321,17'd61322,17'd61323,17'd61324,17'd61325,17'd60937,17'd61326,17'd61327,17'd61328,17'd61329,17'd61330,17'd61331,17'd61332,17'd61333,17'd61333,17'd61209,17'd61334,17'd61335,17'd61336,17'd61337,17'd61086,17'd61213,17'd61338,17'd61339,17'd61340,17'd61341,17'd61217,17'd61342,17'd61343,17'd61344,17'd61220,17'd61221,17'd61221,17'd61345,17'd61223,17'd61346,17'd61226,17'd60087,17'd59689,17'd61347,17'd61348,17'd59559,17'd61349,17'd12698,17'd23676,17'd53774,17'd61350,17'd45209,17'd16915,17'd17235,17'd16327,17'd28232,17'd28233,17'd38365,17'd38502,17'd28350,17'd27349,17'd27737,17'd25528,17'd25670,17'd16203,17'd21505,17'd22992,17'd14264,17'd11396,17'd11274,17'd17236,17'd10605,17'd11527,17'd9739,17'd10743,17'd15187,17'd15944,17'd9194,17'd8878,17'd8412,17'd9887,17'd25148,17'd61351,17'd24546,17'd24710,17'd52404,17'd15440,17'd8108,17'd8259,17'd24869,17'd15691,17'd22138,17'd14533,17'd18454,17'd61352,17'd55833,17'd18335,17'd10483,17'd14266,17'd23518,17'd12120,17'd8250,17'd23343,17'd24711,17'd8571,17'd25147,17'd8733,17'd15435,17'd61353,17'd18569,17'd61354,17'd61355,17'd61356,17'd61357,17'd61358,17'd61359,17'd61360,17'd59715,17'd60981,17'd49879,17'd61361,17'd61113,17'd56638,17'd49785,17'd49882,17'd42597,17'd45036,17'd43285,17'd50461,17'd61362,17'd57844,17'd61243,17'd61363,17'd55722,17'd34459,17'd23733,17'd23217,17'd22680,17'd30427,17'd31343,17'd32344,17'd22860,17'd22325,17'd22327,17'd22329,17'd22680,17'd22677,17'd32190,17'd34882,17'd34882,17'd34759,17'd34759,17'd32190,17'd40523,17'd34278,17'd22680,17'd32827,17'd36986,17'd22329,17'd30277,17'd30277,17'd30277,17'd30277,17'd36986,17'd32827,17'd22680,17'd22330,17'd22325,17'd22504,17'd22500,17'd45616,17'd23569,17'd29975,17'd29526,17'd29243,17'd28851,17'd32353,17'd28850,17'd25438,17'd25438,17'd27511,17'd28369,17'd25317,17'd28600,17'd33643,17'd32658,17'd28723,17'd28130,17'd25567,17'd25835,17'd30903,17'd26403,17'd59213,17'd61364,17'd27148,17'd61365,17'd61366,17'd61246,17'd32037,17'd61367,17'd61368,17'd37919,17'd61369,17'd61370,17'd61371,17'd61372,17'd61373,17'd61374,17'd51751,17'd61375,17'd61376,17'd61377,17'd61378,17'd61379,17'd61380,17'd35312,17'd61381,17'd61382,17'd61383,17'd30460,17'd61384,17'd61385,17'd61386,17'd61387,17'd19833,17'd22727,17'd21439,17'd21744,17'd21434,17'd61388,17'd61389,17'd61390,17'd60501,17'd22933,17'd61391,17'd10881,17'd10881,17'd23109,17'd23279,17'd26216,17'd7008,17'd4994,17'd4841,17'd4683,17'd6067,17'd33992,17'd4998,17'd34657,17'd5156,17'd5157,17'd5162,17'd5166,17'd37030,17'd5164,17'd61140,17'd37433,17'd40397,17'd4690,17'd52011,17'd37033,17'd11435,17'd12011,17'd11715,17'd61392,17'd61393,17'd4383,17'd19857,17'd5489,17'd4384,17'd61394,17'd61395,17'd4039,17'd61396,17'd59232,17'd58483,17'd60755,17'd60756,17'd58852,17'd58732,17'd36317,17'd20857,17'd60506,17'd36742,17'd47267,17'd3193,17'd60877,17'd58617,17'd58616,17'd61397,17'd61398,17'd60759,17'd53431,17'd61399,17'd61400,17'd56208,17'd56423,17'd55878,17'd55072,17'd58874,17'd54013,17'd61401,17'd61402,17'd61403,17'd56431,17'd1942,17'd794,17'd1666,17'd5050,17'd5050,17'd5372,17'd1946,17'd412,17'd602,17'd1529,17'd415,17'd1671,17'd1671,17'd29440,17'd33847,17'd33847,17'd1950,17'd29037,17'd29610,17'd29170,17'd29039,17'd60625,17'd29611,17'd12923,17'd7705,17'd7537,17'd8507,17'd6418,17'd36045,17'd60887,17'd43596,17'd44019,17'd39033,17'd39790,17'd10388,17'd53591,17'd61404,17'd61405,17'd61406,17'd61407,17'd53870,17'd61408,17'd61282,17'd32722,17'd56544,17'd2071,17'd60772,17'd2070,17'd61409,17'd54320,17'd61410
},
'{
17'd10669,17'd3593,17'd10546,17'd3593,17'd52621,17'd52621,17'd1831,17'd4247,17'd2,17'd13,17'd806,17'd465,17'd16389,17'd10,17'd18,17'd18,17'd652,17'd652,17'd16,17'd16,17'd1415,17'd1414,17'd1688,17'd3250,17'd2592,17'd2934,17'd15358,17'd60150,17'd61411,17'd37047,17'd10547,17'd3429,17'd469,17'd1129,17'd2597,17'd2258,17'd3101,17'd15496,17'd5511,17'd52704,17'd3592,17'd12504,17'd986,17'd987,17'd61412,17'd61035,17'd59499,17'd56891,17'd57002,17'd1151,17'd842,17'd311,17'd673,17'd72,17'd69,17'd61413,17'd56796,17'd61414,17'd61415,17'd61416,17'd61417,17'd837,17'd2612,17'd54787,17'd61418,17'd61419,17'd61420,17'd61421,17'd61422,17'd61423,17'd61424,17'd61425,17'd61426,17'd61427,17'd47092,17'd61428,17'd61429,17'd61430,17'd6316,17'd61431,17'd61432,17'd61433,17'd61434,17'd61051,17'd6009,17'd6008,17'd53689,17'd54026,17'd54098,17'd60294,17'd61435,17'd2299,17'd4130,17'd2295,17'd61436,17'd3483,17'd61437,17'd61438,17'd61439,17'd59655,17'd58409,17'd56458,17'd56353,17'd61440,17'd58282,17'd61441,17'd61442,17'd61443,17'd61193,17'd59399,17'd56914,17'd61444,17'd61445,17'd59398,17'd61446,17'd61447,17'd61448,17'd60183,17'd61449,17'd56914,17'd55587,17'd55681,17'd59151,17'd59526,17'd57924,17'd1038,17'd60548,17'd3805,17'd61450,17'd61451,17'd61452,17'd61453,17'd59158,17'd61454,17'd61455,17'd61456,17'd61077,17'd61457,17'd61458,17'd61459,17'd61460,17'd60944,17'd61461,17'd61462,17'd61463,17'd61334,17'd61464,17'd61465,17'd61466,17'd61467,17'd61213,17'd61338,17'd61468,17'd61469,17'd61470,17'd61341,17'd60949,17'd61471,17'd61472,17'd61344,17'd61473,17'd61473,17'd61474,17'd61475,17'd61476,17'd61477,17'd60959,17'd61478,17'd59966,17'd61479,17'd59432,17'd58440,17'd61480,17'd13130,17'd52865,17'd61481,17'd61482,17'd16915,17'd17235,17'd18449,17'd16684,17'd28232,17'd28349,17'd28349,17'd27349,17'd27348,17'd25528,17'd23855,17'd22819,17'd21362,17'd14258,17'd18681,17'd11397,17'd11398,17'd11524,17'd10476,17'd10991,17'd11134,17'd9473,17'd10857,17'd9344,17'd9189,17'd9621,17'd8725,17'd15429,17'd9887,17'd23343,17'd37734,17'd24545,17'd24862,17'd17128,17'd18085,17'd8426,17'd15194,17'd15691,17'd15691,17'd15304,17'd15695,17'd61483,17'd61484,17'd8117,17'd56953,17'd61485,17'd14270,17'd10609,17'd12120,17'd8251,17'd21208,17'd8572,17'd8572,17'd21208,17'd16072,17'd13649,17'd21058,17'd61486,17'd55323,17'd61487,17'd61488,17'd61489,17'd61490,17'd61491,17'd61492,17'd61493,17'd61494,17'd61495,17'd61496,17'd61497,17'd48143,17'd51234,17'd46325,17'd42597,17'd45036,17'd50153,17'd50461,17'd61498,17'd61499,17'd57970,17'd61500,17'd52584,17'd34113,17'd29528,17'd32008,17'd22330,17'd30426,17'd30426,17'd22506,17'd22860,17'd33315,17'd22327,17'd22500,17'd30276,17'd22332,17'd39441,17'd61501,17'd34759,17'd34619,17'd47159,17'd44591,17'd45754,17'd39747,17'd36986,17'd22329,17'd22329,17'd30277,17'd30277,17'd30277,17'd30277,17'd30277,17'd32827,17'd22680,17'd30276,17'd33311,17'd22860,17'd30276,17'd22500,17'd22503,17'd23215,17'd29975,17'd29689,17'd23916,17'd32668,17'd31034,17'd27511,17'd28717,17'd27511,17'd29101,17'd28484,17'd28484,17'd25435,17'd32996,17'd32658,17'd28720,17'd25567,17'd27882,17'd34127,17'd33345,17'd59213,17'd59213,17'd61502,17'd61503,17'd60991,17'd29110,17'd30892,17'd28502,17'd29126,17'd27381,17'd61504,17'd61505,17'd61506,17'd61507,17'd61508,17'd48166,17'd61509,17'd61510,17'd61511,17'd61512,17'd61513,17'd61379,17'd61514,17'd61515,17'd61516,17'd22530,17'd61517,17'd61518,17'd61519,17'd61520,17'd61521,17'd61522,17'd22205,17'd26822,17'd22071,17'd21585,17'd61523,17'd61524,17'd61525,17'd61526,17'd61527,17'd24303,17'd22758,17'd61528,17'd8289,17'd8289,17'd23279,17'd23628,17'd25999,17'd26827,17'd5150,17'd4840,17'd4839,17'd5144,17'd4998,17'd33992,17'd49804,17'd50081,17'd34921,17'd42031,17'd5166,17'd5165,17'd51175,17'd61140,17'd61529,17'd49995,17'd55254,17'd51177,17'd5485,17'd11713,17'd12170,17'd61530,17'd61531,17'd61393,17'd61271,17'd61271,17'd9399,17'd5347,17'd4704,17'd61532,17'd3546,17'd61273,17'd59233,17'd58851,17'd58357,17'd58852,17'd61533,17'd59893,17'd36177,17'd20857,17'd60268,17'd51576,17'd61534,17'd61535,17'd60877,17'd58489,17'd41767,17'd61397,17'd61398,17'd61398,17'd61536,17'd61537,17'd56422,17'd56319,17'd56541,17'd61538,17'd61539,17'd54159,17'd61540,17'd61402,17'd61541,17'd61542,17'd37042,17'd61543,17'd1962,17'd604,17'd5957,17'd5957,17'd6415,17'd2575,17'd951,17'd951,17'd1529,17'd194,17'd1671,17'd1671,17'd33847,17'd2560,17'd29609,17'd26228,17'd27707,17'd29610,17'd29170,17'd29170,17'd29611,17'd35207,17'd11882,17'd8187,17'd6416,17'd6258,17'd6417,17'd36045,17'd16492,17'd43596,17'd44019,17'd12176,17'd39790,17'd18512,17'd61544,17'd61545,17'd61546,17'd61547,17'd19728,17'd54974,17'd61548,17'd61549,17'd32722,17'd58742,17'd53937,17'd60516,17'd56099,17'd59249,17'd61034,17'd61410
},
'{
17'd10669,17'd3593,17'd10546,17'd3429,17'd52621,17'd52621,17'd2422,17'd1688,17'd14,17'd2,17'd2423,17'd465,17'd16389,17'd10,17'd19,17'd18,17'd19,17'd652,17'd16,17'd17187,17'd1415,17'd2596,17'd1689,17'd3250,17'd2592,17'd2593,17'd15358,17'd60150,17'd60150,17'd37047,17'd10802,17'd3429,17'd3752,17'd1129,17'd2596,17'd2258,17'd3101,17'd15496,17'd5511,17'd15359,17'd5204,17'd4738,17'd58504,17'd15497,17'd45,17'd59913,17'd61550,17'd61551,17'd56672,17'd57622,17'd842,17'd840,17'd1982,17'd839,17'd1291,17'd61552,17'd61036,17'd74,17'd61553,17'd18392,17'd59777,17'd670,17'd2789,17'd61554,17'd61169,17'd61555,17'd61556,17'd61557,17'd61558,17'd61559,17'd61560,17'd61561,17'd61562,17'd61563,17'd61564,17'd60289,17'd6135,17'd61565,17'd61566,17'd61567,17'd61568,17'd61569,17'd61570,17'd61051,17'd60909,17'd6008,17'd54099,17'd61571,17'd54026,17'd54098,17'd61435,17'd61572,17'd3638,17'd2467,17'd3636,17'd61573,17'd2015,17'd61574,17'd61575,17'd59792,17'd59934,17'd58277,17'd57019,17'd61576,17'd57278,17'd57517,17'd59790,17'd60055,17'd61577,17'd61578,17'd59150,17'd55784,17'd61579,17'd56355,17'd61580,17'd61581,17'd61582,17'd60059,17'd60177,17'd56583,17'd59395,17'd60060,17'd60309,17'd61583,17'd56699,17'd58775,17'd59404,17'd61584,17'd61585,17'd61320,17'd61586,17'd61587,17'd61588,17'd61589,17'd61590,17'd61591,17'd61592,17'd61593,17'd61594,17'd61595,17'd61330,17'd61081,17'd61596,17'd61597,17'd61598,17'd61334,17'd61464,17'd61599,17'd61465,17'd61467,17'd61213,17'd61600,17'd61601,17'd61602,17'd61603,17'd61604,17'd61605,17'd61606,17'd61607,17'd61608,17'd61609,17'd61473,17'd61610,17'd61611,17'd61612,17'd61346,17'd61094,17'd60215,17'd59688,17'd61347,17'd61613,17'd58926,17'd61614,17'd19151,17'd24850,17'd18321,17'd61615,17'd16915,17'd15571,17'd15811,17'd50314,17'd16327,17'd28233,17'd37738,17'd27234,17'd25528,17'd23855,17'd23168,17'd21362,17'd18443,17'd21985,17'd24029,17'd11275,17'd11399,17'd13886,17'd11527,17'd17839,17'd10742,17'd9344,17'd9346,17'd9189,17'd9042,17'd9195,17'd8730,17'd8576,17'd23343,17'd13374,17'd13374,17'd53189,17'd23866,17'd10860,17'd61616,17'd10481,17'd15194,17'd15691,17'd15691,17'd13378,17'd23180,17'd59704,17'd61352,17'd61617,17'd56735,17'd14818,17'd14270,17'd7619,17'd12120,17'd13258,17'd8579,17'd24545,17'd8573,17'd17126,17'd8250,17'd12589,17'd61618,17'd18570,17'd61619,17'd61620,17'd61621,17'd61622,17'd61623,17'd61624,17'd61625,17'd61493,17'd61626,17'd61495,17'd61496,17'd61627,17'd49571,17'd50902,17'd49274,17'd42597,17'd45036,17'd54480,17'd50069,17'd61628,17'd61629,17'd57970,17'd58826,17'd61630,17'd53331,17'd33801,17'd29829,17'd22328,17'd23573,17'd32344,17'd22506,17'd30276,17'd22325,17'd22326,17'd22500,17'd22680,17'd22856,17'd23926,17'd61501,17'd34882,17'd34759,17'd47159,17'd44591,17'd45492,17'd45379,17'd22329,17'd30277,17'd30277,17'd23215,17'd23215,17'd30277,17'd30277,17'd22329,17'd22331,17'd22856,17'd30276,17'd30276,17'd22332,17'd22856,17'd22500,17'd22329,17'd23217,17'd29826,17'd30879,17'd29533,17'd41730,17'd27511,17'd25438,17'd25438,17'd28850,17'd39591,17'd29970,17'd28600,17'd28721,17'd28253,17'd32658,17'd28594,17'd28597,17'd33008,17'd60988,17'd59213,17'd32211,17'd61631,17'd32374,17'd61632,17'd29252,17'd28731,17'd61633,17'd61634,17'd26080,17'd32205,17'd61635,17'd61636,17'd61637,17'd61638,17'd61639,17'd61640,17'd61641,17'd61642,17'd61643,17'd61644,17'd61645,17'd23752,17'd61646,17'd60604,17'd61647,17'd61648,17'd61649,17'd20340,17'd30153,17'd61650,17'd61651,17'd51009,17'd61652,17'd61653,17'd22056,17'd21585,17'd21585,17'd61654,17'd22924,17'd54592,17'd54496,17'd25996,17'd54672,17'd23110,17'd8911,17'd8289,17'd8289,17'd23628,17'd25999,17'd26827,17'd5150,17'd4841,17'd4839,17'd41891,17'd4998,17'd34657,17'd4526,17'd5157,17'd5329,17'd5167,17'd5166,17'd5010,17'd38318,17'd61655,17'd38847,17'd4527,17'd55254,17'd61656,17'd8309,17'd25229,17'd21007,17'd19095,17'd61657,17'd61658,17'd19232,17'd19232,17'd4213,17'd5347,17'd61394,17'd61659,17'd3546,17'd61660,17'd60023,17'd58851,17'd58357,17'd58484,17'd58733,17'd3690,17'd60266,17'd20857,17'd61661,17'd52911,17'd45652,17'd59236,17'd59236,17'd58492,17'd40095,17'd58616,17'd22602,17'd61662,17'd61663,17'd57098,17'd61664,17'd61665,17'd55755,17'd60509,17'd61539,17'd54084,17'd61666,17'd61667,17'd57242,17'd61668,17'd38070,17'd5935,17'd1680,17'd5372,17'd5372,17'd5372,17'd1946,17'd14178,17'd1383,17'd1383,17'd415,17'd1671,17'd1672,17'd2560,17'd2560,17'd2560,17'd26966,17'd26228,17'd29610,17'd27708,17'd29170,17'd29170,17'd29611,17'd35487,17'd7705,17'd6094,17'd6258,17'd6258,17'd36045,17'd60887,17'd16855,17'd13572,17'd60399,17'd12318,17'd39790,17'd61669,17'd61670,17'd61671,17'd61672,17'd61673,17'd61407,17'd61674,17'd61675,17'd61676,17'd32722,17'd57482,17'd2071,17'd2072,17'd61677,17'd61678,17'd61034,17'd61410
},
'{
17'd10547,17'd52621,17'd3429,17'd3429,17'd52621,17'd10547,17'd3252,17'd2422,17'd1127,17'd2,17'd2423,17'd8814,17'd2591,17'd2591,17'd1275,17'd3905,17'd1128,17'd1128,17'd16,17'd17187,17'd1415,17'd1415,17'd1414,17'd1414,17'd1688,17'd3252,17'd3427,17'd15877,17'd61679,17'd15877,17'd3251,17'd52621,17'd2258,17'd2258,17'd2597,17'd3752,17'd10669,17'd16011,17'd15878,17'd15118,17'd5204,17'd13943,17'd12504,17'd1279,17'd42,17'd61680,17'd61681,17'd61682,17'd60520,17'd61683,17'd57622,17'd1150,17'd1149,17'd70,17'd69,17'd838,17'd61036,17'd60893,17'd74,17'd74,17'd308,17'd670,17'd1710,17'd1288,17'd3265,17'd61684,17'd61685,17'd61686,17'd61687,17'd61688,17'd61689,17'd61690,17'd61691,17'd61692,17'd61297,17'd61693,17'd61694,17'd61695,17'd5687,17'd61696,17'd5850,17'd60910,17'd61697,17'd54625,17'd60909,17'd61698,17'd61431,17'd54262,17'd61699,17'd5852,17'd61055,17'd5546,17'd2299,17'd3960,17'd3480,17'd61436,17'd61700,17'd61701,17'd61702,17'd61703,17'd59655,17'd58409,17'd61704,17'd61705,17'd61706,17'd58653,17'd58157,17'd60306,17'd1034,17'd61707,17'd56811,17'd59401,17'd59273,17'd58769,17'd59525,17'd61708,17'd61709,17'd59399,17'd61710,17'd60545,17'd60308,17'd57649,17'd61711,17'd61712,17'd59526,17'd59284,17'd61713,17'd60668,17'd2687,17'd61714,17'd61715,17'd61716,17'd61717,17'd61718,17'd61719,17'd61720,17'd61721,17'd61722,17'd61723,17'd61724,17'd61725,17'd61726,17'd61727,17'd61728,17'd61729,17'd61463,17'd61730,17'd61464,17'd61731,17'd61732,17'd61733,17'd61734,17'd61734,17'd61603,17'd61735,17'd61736,17'd61734,17'd61215,17'd61737,17'd61608,17'd61609,17'd61738,17'd61739,17'd61740,17'd61475,17'd61741,17'd61742,17'd60958,17'd59827,17'd59554,17'd61743,17'd61744,17'd58193,17'd61745,17'd13507,17'd61746,17'd13758,17'd14672,17'd12860,17'd12415,17'd15811,17'd15687,17'd16560,17'd15571,17'd16558,17'd23855,17'd20452,17'd19408,17'd15185,17'd24029,17'd12423,17'd15176,17'd10603,17'd10603,17'd10606,17'd17839,17'd9478,17'd13887,17'd9039,17'd15684,17'd26498,17'd36625,17'd33404,17'd57186,17'd25678,17'd8419,17'd60710,17'd36204,17'd61747,17'd19034,17'd10341,17'd25930,17'd25930,17'd7457,17'd16075,17'd15194,17'd13894,17'd14939,17'd59978,17'd61748,17'd61749,17'd22140,17'd13529,17'd56167,17'd9351,17'd10860,17'd36204,17'd61750,17'd9887,17'd12865,17'd24042,17'd10608,17'd13649,17'd61751,17'd55125,17'd61752,17'd61753,17'd61754,17'd61755,17'd61756,17'd61757,17'd61758,17'd61759,17'd61760,17'd61761,17'd61762,17'd57710,17'd47332,17'd53562,17'd53203,17'd61763,17'd61764,17'd61765,17'd61766,17'd58212,17'd61767,17'd61768,17'd61769,17'd57325,17'd49976,17'd56966,17'd29376,17'd23216,17'd23038,17'd31343,17'd22160,17'd22324,17'd47457,17'd22326,17'd22330,17'd22680,17'd22856,17'd22324,17'd22324,17'd22325,17'd22500,17'd22500,17'd22500,17'd22326,17'd22327,17'd22502,17'd22501,17'd32191,17'd29828,17'd32191,17'd23215,17'd34453,17'd34882,17'd22333,17'd22681,17'd22856,17'd23038,17'd23038,17'd22678,17'd22331,17'd36986,17'd32191,17'd30275,17'd25032,17'd28850,17'd28369,17'd25438,17'd25179,17'd30432,17'd31034,17'd25317,17'd28600,17'd25566,17'd25565,17'd25565,17'd28720,17'd33000,17'd61770,17'd33345,17'd61364,17'd61771,17'd26066,17'd32212,17'd61772,17'd37912,17'd33326,17'd36560,17'd61634,17'd25188,17'd30600,17'd27043,17'd27656,17'd61773,17'd61774,17'd59469,17'd31378,17'd61775,17'd61776,17'd61777,17'd61778,17'd61779,17'd61780,17'd61781,17'd61782,17'd61783,17'd61648,17'd61784,17'd61785,17'd30610,17'd61786,17'd61787,17'd61788,17'd20813,17'd22073,17'd22211,17'd38051,17'd40981,17'd21592,17'd61789,17'd21904,17'd57588,17'd24943,17'd12443,17'd25768,17'd23110,17'd23110,17'd8607,17'd10881,17'd24645,17'd7325,17'd4994,17'd4842,17'd31716,17'd5000,17'd34157,17'd55350,17'd49804,17'd31552,17'd4842,17'd5158,17'd5329,17'd4849,17'd54498,17'd49996,17'd61790,17'd39015,17'd60387,17'd61791,17'd6397,17'd11860,17'd61792,17'd21778,17'd61793,17'd19096,17'd19096,17'd19233,17'd19233,17'd61794,17'd61795,17'd61796,17'd61797,17'd60753,17'd61396,17'd59232,17'd58483,17'd58731,17'd58850,17'd61533,17'd36038,17'd61798,17'd60504,17'd60268,17'd61799,17'd39479,17'd41767,17'd41767,17'd41767,17'd61800,17'd58856,17'd61801,17'd61802,17'd61400,17'd53864,17'd61803,17'd61804,17'd53865,17'd60882,17'd59903,17'd54084,17'd61805,17'd61806,17'd56108,17'd36453,17'd9246,17'd2558,17'd3246,17'd35907,17'd5630,17'd12496,17'd2393,17'd14178,17'd413,17'd15233,17'd15233,17'd2394,17'd1672,17'd2560,17'd29169,17'd32082,17'd27707,17'd27707,17'd27708,17'd27708,17'd28545,17'd29892,17'd29611,17'd35487,17'd7537,17'd6417,17'd6258,17'd16492,17'd16492,17'd37959,17'd13420,17'd12913,17'd61807,17'd12318,17'd41004,17'd61808,17'd61809,17'd10247,17'd61810,17'd61811,17'd61812,17'd54323,17'd54162,17'd55472,17'd32722,17'd59242,17'd57482,17'd61677,17'd61813,17'd61814,17'd54320,17'd61815
},
'{
17'd10547,17'd52621,17'd3429,17'd3429,17'd52621,17'd10547,17'd2935,17'd2422,17'd1689,17'd2,17'd2423,17'd8814,17'd4242,17'd2591,17'd283,17'd13,17'd1128,17'd1128,17'd16,17'd17187,17'd2936,17'd1415,17'd1416,17'd1414,17'd1688,17'd2422,17'd3427,17'd15496,17'd52704,17'd15877,17'd3428,17'd2935,17'd2258,17'd2425,17'd2597,17'd3752,17'd3593,17'd16501,17'd15878,17'd15118,17'd5204,17'd4086,17'd16392,17'd58016,17'd61816,17'd61817,17'd61818,17'd61035,17'd61819,17'd61820,17'd57622,17'd56114,17'd1429,17'd70,17'd69,17'd1291,17'd838,17'd60892,17'd56796,17'd56796,17'd308,17'd670,17'd1843,17'd1288,17'd1428,17'd55086,17'd61821,17'd61822,17'd61823,17'd61824,17'd61825,17'd61826,17'd61827,17'd61828,17'd61829,17'd61830,17'd61694,17'd61831,17'd6135,17'd61832,17'd61833,17'd60532,17'd60650,17'd53526,17'd60909,17'd61698,17'd61834,17'd53374,17'd61835,17'd5851,17'd53759,17'd61435,17'd4932,17'd54022,17'd3143,17'd3636,17'd3960,17'd61836,17'd61837,17'd61838,17'd57134,17'd59017,17'd61839,17'd61840,17'd57019,17'd61189,17'd59018,17'd59649,17'd61841,17'd61193,17'd56811,17'd59150,17'd59524,17'd60795,17'd61842,17'd61843,17'd61844,17'd61845,17'd61846,17'd61710,17'd60545,17'd59282,17'd59656,17'd59797,17'd61847,17'd56915,17'd61848,17'd59027,17'd61849,17'd61850,17'd61851,17'd61852,17'd61853,17'd61854,17'd61855,17'd61856,17'd61857,17'd61858,17'd61859,17'd61724,17'd61860,17'd61861,17'd61862,17'd61863,17'd61864,17'd61598,17'd61730,17'd61865,17'd61866,17'd61731,17'd61867,17'd61868,17'd61869,17'd61736,17'd61870,17'd61871,17'd61872,17'd61873,17'd61874,17'd61607,17'd61875,17'd61609,17'd61610,17'd61876,17'd61611,17'd61877,17'd61878,17'd61742,17'd60215,17'd61879,17'd61479,17'd59432,17'd58565,17'd61097,17'd13128,17'd56493,17'd61880,17'd16799,17'd12860,17'd18564,17'd12415,17'd14672,17'd14672,17'd14672,17'd18564,17'd12254,17'd22819,17'd18198,17'd19158,17'd10854,17'd11401,17'd19642,17'd10606,17'd17720,17'd17839,17'd9619,17'd13887,17'd9188,17'd9195,17'd9195,17'd36073,17'd61881,17'd24545,17'd21208,17'd7947,17'd17609,17'd15301,17'd23687,17'd41031,17'd15439,17'd8258,17'd8108,17'd26040,17'd7620,17'd23867,17'd7791,17'd14817,17'd18088,17'd59842,17'd61748,17'd60466,17'd19161,17'd14533,17'd14012,17'd9623,17'd7786,17'd23174,17'd61882,17'd8579,17'd8417,17'd61883,17'd14527,17'd53190,17'd61884,17'd59705,17'd61885,17'd61886,17'd61887,17'd61888,17'd61889,17'd61890,17'd61758,17'd61891,17'd61892,17'd61893,17'd61894,17'd61895,17'd47436,17'd46554,17'd53203,17'd61896,17'd61764,17'd61897,17'd61898,17'd58212,17'd61899,17'd61900,17'd61901,17'd50734,17'd61902,17'd53405,17'd31502,17'd29828,17'd22679,17'd22332,17'd22681,17'd22860,17'd22504,17'd22330,17'd22331,17'd22678,17'd22677,17'd22506,17'd22332,17'd22331,17'd36986,17'd22329,17'd22326,17'd22326,17'd22326,17'd22501,17'd32351,17'd32191,17'd29374,17'd32191,17'd30277,17'd45492,17'd39281,17'd22505,17'd22860,17'd22333,17'd22677,17'd22677,17'd23038,17'd22679,17'd23217,17'd29376,17'd32659,17'd29103,17'd25317,17'd25709,17'd25177,17'd32353,17'd33318,17'd28850,17'd28484,17'd28721,17'd32658,17'd25708,17'd27766,17'd27638,17'd28717,17'd25318,17'd59213,17'd33020,17'd61903,17'd35995,17'd34888,17'd38037,17'd31676,17'd29999,17'd36560,17'd32199,17'd25043,17'd26086,17'd28876,17'd61904,17'd35871,17'd61905,17'd61906,17'd61907,17'd61908,17'd61909,17'd61910,17'd61911,17'd60126,17'd61912,17'd61913,17'd61914,17'd61915,17'd61916,17'd61917,17'd61918,17'd25348,17'd61919,17'd61920,17'd24626,17'd20520,17'd22573,17'd61921,17'd61922,17'd29153,17'd61923,17'd21908,17'd61924,17'd23792,17'd54410,17'd53504,17'd25768,17'd25768,17'd23110,17'd23278,17'd10881,17'd7657,17'd24647,17'd4993,17'd31245,17'd28536,17'd4525,17'd61925,17'd61926,17'd39015,17'd31716,17'd61927,17'd5331,17'd5160,17'd4849,17'd50835,17'd55457,17'd54862,17'd60387,17'd61928,17'd36890,17'd11041,17'd12477,17'd61929,17'd61930,17'd61793,17'd61931,17'd61931,17'd61932,17'd61932,17'd10521,17'd6864,17'd61144,17'd49601,17'd3691,17'd61798,17'd59232,17'd58483,17'd58356,17'd58731,17'd58852,17'd36038,17'd60267,17'd20857,17'd59753,17'd46237,17'd61933,17'd61397,17'd40095,17'd22775,17'd42329,17'd39323,17'd36595,17'd61800,17'd56774,17'd61934,17'd61935,17'd61804,17'd56541,17'd60882,17'd59763,17'd61936,17'd61937,17'd61938,17'd56327,17'd36747,17'd9247,17'd5195,17'd3391,17'd49008,17'd12496,17'd2393,17'd16256,17'd16256,17'd12644,17'd12644,17'd15233,17'd2394,17'd1950,17'd1950,17'd32082,17'd27707,17'd27707,17'd29610,17'd29170,17'd29170,17'd27709,17'd29892,17'd35207,17'd38460,17'd6418,17'd36045,17'd37959,17'd16492,17'd16492,17'd37959,17'd13420,17'd13572,17'd61807,17'd45291,17'd41004,17'd61939,17'd61940,17'd61941,17'd61942,17'd5625,17'd61812,17'd2542,17'd41621,17'd55563,17'd32722,17'd59769,17'd59623,17'd55073,17'd61943,17'd61944,17'd61945,17'd61815
},
'{
17'd10802,17'd52621,17'd3429,17'd3429,17'd52621,17'd10802,17'd10669,17'd3429,17'd1689,17'd14,17'd2423,17'd8814,17'd2933,17'd2591,17'd283,17'd12,17'd1128,17'd1128,17'd18,17'd16,17'd17187,17'd1415,17'd1416,17'd1416,17'd2257,17'd3429,17'd2934,17'd15496,17'd5511,17'd15877,17'd3428,17'd3101,17'd2597,17'd2258,17'd2597,17'd3752,17'd3593,17'd12505,17'd57896,17'd15878,17'd5204,17'd5204,17'd16392,17'd14320,17'd15497,17'd60404,17'd61946,17'd59251,17'd61947,17'd61948,17'd60040,17'd56438,17'd61949,17'd1429,17'd69,17'd1291,17'd61037,17'd838,17'd1000,17'd839,17'd306,17'd486,17'd1843,17'd1709,17'd1288,17'd61950,17'd61951,17'd61952,17'd61953,17'd61954,17'd61294,17'd61423,17'd61690,17'd61955,17'd61956,17'd61957,17'd61958,17'd61695,17'd61428,17'd61959,17'd61960,17'd61961,17'd61962,17'd5852,17'd6009,17'd53818,17'd61963,17'd61964,17'd52852,17'd60904,17'd54354,17'd60163,17'd2657,17'd4931,17'd2989,17'd61965,17'd2978,17'd61966,17'd61967,17'd61968,17'd61703,17'd57134,17'd61969,17'd61970,17'd61971,17'd61189,17'd61972,17'd59519,17'd59932,17'd60425,17'd58661,17'd59147,17'd58887,17'd57518,17'd57397,17'd59521,17'd61973,17'd61580,17'd60793,17'd59796,17'd60427,17'd60427,17'd61449,17'd59276,17'd58773,17'd61974,17'd61975,17'd59286,17'd61976,17'd61977,17'd61978,17'd61979,17'd61980,17'd61981,17'd60437,17'd61982,17'd61983,17'd61984,17'd61985,17'd61986,17'd61987,17'd61988,17'd61989,17'd60945,17'd61990,17'd61991,17'd61730,17'd61865,17'd61992,17'd61993,17'd61867,17'd61994,17'd61995,17'd61996,17'd61870,17'd61997,17'd61735,17'd61998,17'd61215,17'd61737,17'd61999,17'd62000,17'd62001,17'd61739,17'd61876,17'd62002,17'd61345,17'd61878,17'd60958,17'd62003,17'd59555,17'd60826,17'd59060,17'd57680,17'd15171,17'd53896,17'd52484,17'd18684,17'd12997,17'd15434,17'd12418,17'd14523,17'd14930,17'd14930,17'd12254,17'd16203,17'd18198,17'd18917,17'd13762,17'd11131,17'd10331,17'd19642,17'd10479,17'd11134,17'd12116,17'd9480,17'd9038,17'd8723,17'd8724,17'd8570,17'd61881,17'd17729,17'd11967,17'd13005,17'd62004,17'd14136,17'd17241,17'd54378,17'd12266,17'd23689,17'd15572,17'd10747,17'd18921,17'd10342,17'd7622,17'd13528,17'd62005,17'd60969,17'd62006,17'd12269,17'd60100,17'd12268,17'd12430,17'd24045,17'd42228,17'd17238,17'd25289,17'd15301,17'd8580,17'd8418,17'd10608,17'd10745,17'd41031,17'd62007,17'd62008,17'd21677,17'd62009,17'd62010,17'd62011,17'd62012,17'd62013,17'd61758,17'd62014,17'd62015,17'd62016,17'd61894,17'd62017,17'd47436,17'd49880,17'd50264,17'd61896,17'd61764,17'd61897,17'd54568,17'd62018,17'd62019,17'd62020,17'd62021,17'd62022,17'd62023,17'd62024,17'd31032,17'd30128,17'd41273,17'd22330,17'd22325,17'd22325,17'd22326,17'd22326,17'd22329,17'd22331,17'd22680,17'd22856,17'd22680,17'd36986,17'd30277,17'd33158,17'd33158,17'd22502,17'd22502,17'd33158,17'd32351,17'd32191,17'd32191,17'd23215,17'd22329,17'd33311,17'd22681,17'd22860,17'd22333,17'd22159,17'd35292,17'd22159,17'd22677,17'd23389,17'd23386,17'd30431,17'd25031,17'd41730,17'd29244,17'd27637,17'd25178,17'd32353,17'd41730,17'd28369,17'd25435,17'd28253,17'd28253,17'd28723,17'd28130,17'd27882,17'd25320,17'd60989,17'd59869,17'd36268,17'd26066,17'd62025,17'd62026,17'd28733,17'd62027,17'd30453,17'd29698,17'd28732,17'd26196,17'd25854,17'd28747,17'd62028,17'd62029,17'd62030,17'd62031,17'd62032,17'd62033,17'd62034,17'd62035,17'd62036,17'd62037,17'd62038,17'd24768,17'd27538,17'd62039,17'd62040,17'd62041,17'd62042,17'd62043,17'd62044,17'd62045,17'd21890,17'd62046,17'd62047,17'd60749,17'd60749,17'd62048,17'd62049,17'd22064,17'd30792,17'd22932,17'd22586,17'd54956,17'd25768,17'd30636,17'd23110,17'd24644,17'd8289,17'd7659,17'd24648,17'd4993,17'd28418,17'd28536,17'd4999,17'd61925,17'd38848,17'd49995,17'd37153,17'd25627,17'd5335,17'd5166,17'd51663,17'd51326,17'd4370,17'd4370,17'd50587,17'd38193,17'd62050,17'd12009,17'd62051,17'd20554,17'd62052,17'd19095,17'd11583,17'd61931,17'd62053,17'd62054,17'd10521,17'd4546,17'd62055,17'd49601,17'd3691,17'd61660,17'd60619,17'd3543,17'd60756,17'd58852,17'd58732,17'd49004,17'd20857,17'd62056,17'd62057,17'd62058,17'd62059,17'd58857,17'd37039,17'd62060,17'd2879,17'd62061,17'd61662,17'd62062,17'd58620,17'd62063,17'd55877,17'd62064,17'd54971,17'd62065,17'd58874,17'd62066,17'd62067,17'd56216,17'd39626,17'd1942,17'd62068,17'd4424,17'd3391,17'd5630,17'd12496,17'd14178,17'd2098,17'd2098,17'd12644,17'd12644,17'd15233,17'd27094,17'd1950,17'd1950,17'd27707,17'd27707,17'd27708,17'd27708,17'd29170,17'd29170,17'd29892,17'd29610,17'd36602,17'd11061,17'd8186,17'd6095,17'd38459,17'd37959,17'd16492,17'd37959,17'd13176,17'd17546,17'd12635,17'd51098,17'd62069,17'd62069,17'd12317,17'd62070,17'd62071,17'd62072,17'd62073,17'd3059,17'd54162,17'd55563,17'd56101,17'd59130,17'd57482,17'd62074,17'd62075,17'd61944,17'd61945,17'd62076
},
'{
17'd10670,17'd10669,17'd3593,17'd3429,17'd10669,17'd10802,17'd10802,17'd10669,17'd3250,17'd1127,17'd12,17'd8814,17'd2933,17'd465,17'd283,17'd12,17'd1128,17'd1128,17'd18,17'd16,17'd17187,17'd1415,17'd17,17'd1414,17'd2597,17'd3429,17'd2593,17'd3592,17'd5511,17'd5511,17'd3592,17'd3427,17'd3752,17'd2258,17'd2258,17'd3752,17'd10546,17'd11071,17'd16501,17'd62077,17'd5204,17'd5511,17'd16392,17'd13944,17'd59381,17'd60519,17'd62078,17'd60774,17'd60280,17'd61947,17'd56672,17'd56892,17'd1150,17'd1429,17'd839,17'd69,17'd62079,17'd61037,17'd838,17'd70,17'd306,17'd487,17'd837,17'd55276,17'd54787,17'd62080,17'd61038,17'd62081,17'd62082,17'd2634,17'd62083,17'd61689,17'd62084,17'd62085,17'd62086,17'd62087,17'd61958,17'd62088,17'd15012,17'd62089,17'd62090,17'd62091,17'd62092,17'd6007,17'd62093,17'd61963,17'd43201,17'd52852,17'd6005,17'd62094,17'd62095,17'd60293,17'd5413,17'd2822,17'd2980,17'd59928,17'd62096,17'd61305,17'd62097,17'd62098,17'd61838,17'd62099,17'd62100,17'd62101,17'd62102,17'd55091,17'd62103,17'd56907,17'd59274,17'd62104,17'd60052,17'd62105,17'd59933,17'd60427,17'd60660,17'd62106,17'd62107,17'd62108,17'd62109,17'd59397,17'd60427,17'd59024,17'd61313,17'd60541,17'd59399,17'd62110,17'd62111,17'd62112,17'd62113,17'd2850,17'd62114,17'd62115,17'd62116,17'd62117,17'd62118,17'd62119,17'd62120,17'd62121,17'd62122,17'd62123,17'd61329,17'd62124,17'd62125,17'd61989,17'd62126,17'd62127,17'd62128,17'd62129,17'd62130,17'd62130,17'd61993,17'd62131,17'd62132,17'd61996,17'd61871,17'd62133,17'd62134,17'd61603,17'd61873,17'd61874,17'd62135,17'd61999,17'd62001,17'd62136,17'd61876,17'd61876,17'd62137,17'd60824,17'd62138,17'd62139,17'd60088,17'd61743,17'd59560,17'd60964,17'd62140,17'd13507,17'd52866,17'd12574,17'd12256,17'd15434,17'd12418,17'd12418,17'd12416,17'd12416,17'd12253,17'd15184,17'd15053,17'd12996,17'd11807,17'd11131,17'd11671,17'd16680,17'd17718,17'd16561,17'd17717,17'd10173,17'd16067,17'd8569,17'd12425,17'd24368,17'd26259,17'd26260,17'd24213,17'd17483,17'd62141,17'd62142,17'd10860,17'd10746,17'd61616,17'd23689,17'd10996,17'd18921,17'd19536,17'd17018,17'd8427,17'd19648,17'd19421,17'd55125,17'd62143,17'd21676,17'd12431,17'd8429,17'd19648,17'd9891,17'd24548,17'd14385,17'd17354,17'd21824,17'd8419,17'd53035,17'd7946,17'd10179,17'd62144,17'd62145,17'd62146,17'd11538,17'd62147,17'd62148,17'd62149,17'd62150,17'd62151,17'd61492,17'd62152,17'd62153,17'd62154,17'd61762,17'd62155,17'd55232,17'd50651,17'd57972,17'd61896,17'd61764,17'd62156,17'd62157,17'd62018,17'd62158,17'd62159,17'd62020,17'd62160,17'd55328,17'd62161,17'd54057,17'd23388,17'd23389,17'd36986,17'd22326,17'd45616,17'd51229,17'd22502,17'd22503,17'd22328,17'd22327,17'd45874,17'd22502,17'd22501,17'd32008,17'd23569,17'd29974,17'd37116,17'd36543,17'd29974,17'd32008,17'd32191,17'd37386,17'd23217,17'd36986,17'd22505,17'd22860,17'd22506,17'd30426,17'd22507,17'd22507,17'd22158,17'd22332,17'd30128,17'd24086,17'd29533,17'd25179,17'd25179,17'd25180,17'd29976,17'd30432,17'd29103,17'd27511,17'd28594,17'd25708,17'd28483,17'd33643,17'd28484,17'd27511,17'd29244,17'd30432,17'd62162,17'd39142,17'd25836,17'd62163,17'd62164,17'd29255,17'd27524,17'd30443,17'd31041,17'd30144,17'd62165,17'd25576,17'd25592,17'd28390,17'd35871,17'd62166,17'd62167,17'd62168,17'd62169,17'd62170,17'd62171,17'd62172,17'd62173,17'd62174,17'd62175,17'd24614,17'd62176,17'd28280,17'd23238,17'd62177,17'd62178,17'd30154,17'd62179,17'd62180,17'd62181,17'd22229,17'd21897,17'd62182,17'd60500,17'd58969,17'd21903,17'd22741,17'd62183,17'd24304,17'd22586,17'd26111,17'd25768,17'd30636,17'd23110,17'd24644,17'd24149,17'd62184,17'd5607,17'd4993,17'd28418,17'd5328,17'd41891,17'd55350,17'd54862,17'd38567,17'd5008,17'd5160,17'd5335,17'd5166,17'd51663,17'd61928,17'd38568,17'd60387,17'd51248,17'd36588,17'd10900,17'd17286,17'd20256,17'd12171,17'd62052,17'd19095,17'd11583,17'd61931,17'd62185,17'd62186,17'd61794,17'd6864,17'd62187,17'd49601,17'd3691,17'd61798,17'd3543,17'd49004,17'd58852,17'd58733,17'd59893,17'd36317,17'd60268,17'd62188,17'd62058,17'd62058,17'd62189,17'd46789,17'd53060,17'd39479,17'd62190,17'd62191,17'd62192,17'd57742,17'd62193,17'd62063,17'd62194,17'd55755,17'd28652,17'd62195,17'd62196,17'd61805,17'd61938,17'd56432,17'd38330,17'd62197,17'd62198,17'd3742,17'd5372,17'd3073,17'd2393,17'd2098,17'd6721,17'd6721,17'd12644,17'd12644,17'd2394,17'd29169,17'd1950,17'd1949,17'd27707,17'd27707,17'd27708,17'd29170,17'd29170,17'd29170,17'd29892,17'd35207,17'd11882,17'd7537,17'd6258,17'd38459,17'd38459,17'd38459,17'd16492,17'd37959,17'd13176,17'd17546,17'd12635,17'd62199,17'd62200,17'd62201,17'd62202,17'd62203,17'd62204,17'd62205,17'd4222,17'd2724,17'd53672,17'd55563,17'd56101,17'd62206,17'd56544,17'd62074,17'd53287,17'd62207,17'd54684,17'd62208
},
'{
17'd10925,17'd10802,17'd3593,17'd3593,17'd10669,17'd10802,17'd10924,17'd10669,17'd3429,17'd1414,17'd3905,17'd1128,17'd21,17'd10,17'd979,17'd18,17'd1128,17'd1128,17'd18,17'd16,17'd17187,17'd1415,17'd17,17'd1416,17'd1414,17'd3752,17'd2935,17'd3901,17'd5204,17'd5511,17'd15496,17'd3428,17'd52621,17'd52621,17'd2426,17'd3429,17'd3593,17'd11071,17'd16501,17'd62077,17'd5511,17'd5511,17'd5204,17'd13945,17'd62209,17'd42,17'd61680,17'd59913,17'd59627,17'd60280,17'd56672,17'd57002,17'd1151,17'd56795,17'd839,17'd839,17'd62210,17'd60894,17'd1291,17'd69,17'd69,17'd69,17'd488,17'd671,17'd62211,17'd62212,17'd54787,17'd62213,17'd62214,17'd62215,17'd62216,17'd62217,17'd62218,17'd62219,17'd62220,17'd62221,17'd47092,17'd61958,17'd47092,17'd47092,17'd61693,17'd62222,17'd62223,17'd3471,17'd6000,17'd62224,17'd62224,17'd6472,17'd6631,17'd6006,17'd62225,17'd60532,17'd62226,17'd62226,17'd2825,17'd62227,17'd3304,17'd2644,17'd62228,17'd61967,17'd61058,17'd61439,17'd59017,17'd1459,17'd58772,17'd57133,17'd56579,17'd57646,17'd59014,17'd62229,17'd59147,17'd60052,17'd59019,17'd60302,17'd60427,17'd62230,17'd60792,17'd61973,17'd62231,17'd58773,17'd61449,17'd62232,17'd62232,17'd59145,17'd60308,17'd56355,17'd61847,17'd62233,17'd58664,17'd1188,17'd62234,17'd62235,17'd62236,17'd62237,17'd62238,17'd62239,17'd62240,17'd61180,17'd62241,17'd61723,17'd62242,17'd62243,17'd62244,17'd62245,17'd62246,17'd62247,17'd62128,17'd61865,17'd62248,17'd62249,17'd62250,17'd62251,17'd62132,17'd62132,17'd62252,17'd62133,17'd62253,17'd61735,17'd61604,17'd61215,17'd62254,17'd62255,17'd62256,17'd62257,17'd62258,17'd61739,17'd61610,17'd61610,17'd61222,17'd60958,17'd60087,17'd59429,17'd59431,17'd62259,17'd62260,17'd12706,17'd62261,17'd62262,17'd12257,17'd12253,17'd12414,17'd12856,17'd12417,17'd12417,17'd12414,17'd13882,17'd11806,17'd11962,17'd11807,17'd10854,17'd9883,17'd16549,17'd37607,17'd17232,17'd16552,17'd24212,17'd23861,17'd8730,17'd8731,17'd31760,17'd26260,17'd11967,17'd12867,17'd22648,17'd62263,17'd62264,17'd35090,17'd23177,17'd62265,17'd14011,17'd16567,17'd18921,17'd15691,17'd15194,17'd16692,17'd15306,17'd12268,17'd23348,17'd62266,17'd23875,17'd13008,17'd8429,17'd13894,17'd9891,17'd18451,17'd16802,17'd8255,17'd33716,17'd17483,17'd8251,17'd7947,17'd10995,17'd62267,17'd15062,17'd62268,17'd62269,17'd62270,17'd62271,17'd62272,17'd62273,17'd62274,17'd62275,17'd62152,17'd62152,17'd62276,17'd61762,17'd62277,17'd57570,17'd51075,17'd54840,17'd62278,17'd62279,17'd62280,17'd62281,17'd61628,17'd62282,17'd62283,17'd62284,17'd62285,17'd62286,17'd62287,17'd62288,17'd44715,17'd34277,17'd41273,17'd22329,17'd33158,17'd36543,17'd33158,17'd22502,17'd22502,17'd22502,17'd51229,17'd45616,17'd36543,17'd23569,17'd29829,17'd29974,17'd29974,17'd23569,17'd29974,17'd23569,17'd29828,17'd37386,17'd23216,17'd36986,17'd30276,17'd22681,17'd30426,17'd22158,17'd22162,17'd22162,17'd30427,17'd30425,17'd23918,17'd28977,17'd33483,17'd25178,17'd25032,17'd25031,17'd38667,17'd33483,17'd29101,17'd27765,17'd27766,17'd25565,17'd28483,17'd42749,17'd28850,17'd30432,17'd32668,17'd33802,17'd62289,17'd59343,17'd61631,17'd39915,17'd38161,17'd30594,17'd30146,17'd30290,17'd29543,17'd30452,17'd26540,17'd26297,17'd25449,17'd62290,17'd23410,17'd62291,17'd62292,17'd62293,17'd62294,17'd62295,17'd62296,17'd62297,17'd62298,17'd62299,17'd62300,17'd62301,17'd62302,17'd20946,17'd24280,17'd62303,17'd62304,17'd22895,17'd62305,17'd24626,17'd20369,17'd62306,17'd62307,17'd21586,17'd62308,17'd22225,17'd22064,17'd23622,17'd62309,17'd24304,17'd22758,17'd22758,17'd26111,17'd26111,17'd23628,17'd25223,17'd7324,17'd7008,17'd5608,17'd4840,17'd5328,17'd40397,17'd55350,17'd54765,17'd49895,17'd50586,17'd5162,17'd5166,17'd5166,17'd5010,17'd51663,17'd61928,17'd38568,17'd38320,17'd57868,17'd6397,17'd25772,17'd12629,17'd22947,17'd62310,17'd62311,17'd62312,17'd29885,17'd29742,17'd11324,17'd62313,17'd4215,17'd61272,17'd62314,17'd49601,17'd3691,17'd61396,17'd60504,17'd58732,17'd58852,17'd62315,17'd49106,17'd20857,17'd59754,17'd50921,17'd62316,17'd62317,17'd62317,17'd62318,17'd46789,17'd37039,17'd62319,17'd62320,17'd62321,17'd56097,17'd62322,17'd56209,17'd56320,17'd62323,17'd62324,17'd62325,17'd62326,17'd62327,17'd62328,17'd19361,17'd1665,17'd7850,17'd2765,17'd6407,17'd6415,17'd14178,17'd2393,17'd2098,17'd779,17'd779,17'd12644,17'd12644,17'd33847,17'd1950,17'd1950,17'd26228,17'd26228,17'd26228,17'd27708,17'd29170,17'd29170,17'd29170,17'd29612,17'd35207,17'd11061,17'd8507,17'd6095,17'd4867,17'd4867,17'd38072,17'd14060,17'd13933,17'd43596,17'd43596,17'd62329,17'd62330,17'd62331,17'd14434,17'd17913,17'd18269,17'd62332,17'd62333,17'd4707,17'd41903,17'd41476,17'd62334,17'd62335,17'd56425,17'd62336,17'd62074,17'd25889,17'd62337,17'd54684,17'd62338
},
'{
17'd10925,17'd10924,17'd3593,17'd3593,17'd10669,17'd10802,17'd10924,17'd11071,17'd10669,17'd2597,17'd3905,17'd1128,17'd11,17'd10,17'd979,17'd19,17'd18,17'd18,17'd16,17'd16,17'd17187,17'd1415,17'd17,17'd1414,17'd2596,17'd10268,17'd2784,17'd2934,17'd15496,17'd5511,17'd15877,17'd15496,17'd10802,17'd52621,17'd2426,17'd2258,17'd3429,17'd11071,17'd16501,17'd62077,17'd5511,17'd5511,17'd5204,17'd4737,17'd14189,17'd61816,17'd62339,17'd60037,17'd60279,17'd60039,17'd60039,17'd56672,17'd56892,17'd1430,17'd56795,17'd839,17'd60894,17'd60894,17'd485,17'd1981,17'd69,17'd1291,17'd489,17'd62340,17'd62341,17'd62342,17'd2437,17'd62343,17'd62344,17'd2282,17'd62345,17'd62346,17'd62347,17'd62348,17'd62349,17'd62350,17'd62351,17'd47092,17'd61564,17'd47092,17'd31269,17'd61693,17'd62352,17'd62353,17'd3470,17'd6006,17'd44863,17'd6150,17'd5841,17'd5999,17'd6308,17'd62354,17'd5412,17'd60293,17'd2825,17'd4930,17'd59640,17'd53609,17'd62355,17'd62097,17'd61837,17'd61838,17'd61439,17'd55778,17'd58406,17'd62356,17'd56454,17'd55582,17'd58041,17'd57393,17'd58888,17'd60051,17'd60308,17'd58038,17'd56697,17'd59938,17'd61846,17'd62357,17'd61973,17'd62358,17'd62359,17'd57918,17'd59275,17'd59024,17'd59273,17'd59272,17'd60793,17'd62360,17'd58665,17'd62361,17'd62362,17'd62363,17'd62364,17'd62365,17'd62366,17'd62367,17'd62368,17'd60786,17'd61455,17'd62369,17'd62370,17'd61329,17'd61595,17'd61080,17'd60944,17'd62371,17'd62372,17'd62373,17'd62374,17'd62249,17'd62375,17'd62376,17'd62377,17'd62132,17'd61996,17'd61997,17'd62253,17'd62133,17'd61736,17'd61339,17'd62378,17'd62379,17'd62380,17'd62381,17'd62382,17'd62383,17'd62136,17'd61610,17'd61221,17'd61742,17'd60215,17'd60088,17'd61743,17'd62384,17'd62385,17'd57815,17'd22470,17'd21501,17'd15808,17'd12253,17'd12109,17'd12109,17'd12995,17'd16321,17'd15184,17'd13761,17'd20313,17'd16797,17'd11395,17'd10990,17'd11134,17'd9480,17'd9743,17'd26498,17'd16317,17'd16205,17'd8730,17'd8575,17'd24711,17'd24545,17'd11811,17'd53107,17'd8580,17'd14676,17'd7787,17'd23518,17'd62386,17'd7955,17'd23689,17'd62387,17'd18921,17'd16567,17'd15442,17'd15304,17'd62388,17'd62389,17'd18690,17'd62390,17'd62391,17'd8431,17'd55030,17'd23180,17'd24552,17'd10342,17'd18451,17'd11534,17'd13140,17'd12427,17'd18203,17'd17241,17'd11968,17'd15193,17'd62392,17'd8430,17'd62393,17'd17978,17'd62394,17'd62395,17'd62396,17'd62273,17'd62397,17'd62275,17'd61891,17'd62398,17'd62399,17'd61762,17'd62277,17'd57570,17'd51075,17'd54840,17'd62278,17'd52982,17'd62400,17'd62281,17'd62160,17'd62158,17'd62401,17'd62402,17'd62159,17'd58095,17'd62403,17'd62404,17'd36414,17'd37673,17'd23569,17'd32008,17'd23388,17'd23388,17'd29974,17'd50732,17'd37116,17'd37116,17'd36543,17'd36543,17'd29974,17'd30579,17'd23567,17'd23567,17'd37511,17'd29974,17'd32008,17'd32351,17'd23215,17'd23218,17'd36986,17'd22680,17'd22506,17'd22161,17'd32660,17'd32660,17'd32660,17'd30427,17'd39131,17'd29530,17'd33482,17'd53720,17'd29976,17'd25030,17'd28977,17'd38808,17'd38667,17'd29103,17'd28369,17'd28723,17'd25833,17'd25833,17'd32658,17'd28484,17'd29103,17'd32668,17'd33793,17'd34113,17'd62405,17'd59869,17'd26662,17'd32370,17'd30444,17'd33169,17'd36418,17'd30756,17'd27265,17'd27664,17'd28152,17'd25967,17'd28624,17'd24109,17'd62406,17'd62407,17'd62408,17'd62409,17'd62410,17'd62411,17'd62412,17'd62413,17'd25202,17'd61784,17'd62414,17'd62415,17'd62040,17'd21559,17'd62416,17'd62417,17'd62418,17'd62419,17'd62420,17'd21576,17'd62421,17'd28771,17'd61524,17'd62422,17'd22069,17'd22224,17'd22223,17'd23971,17'd24304,17'd24305,17'd30793,17'd22758,17'd26111,17'd26111,17'd23628,17'd62423,17'd7007,17'd4994,17'd32552,17'd32552,17'd4841,17'd5155,17'd39470,17'd54673,17'd4527,17'd5006,17'd5163,17'd5011,17'd5010,17'd52271,17'd52095,17'd38444,17'd60387,17'd38193,17'd62424,17'd8004,17'd25633,17'd24806,17'd12909,17'd62425,17'd62426,17'd62426,17'd18978,17'd29885,17'd62427,17'd11324,17'd5176,17'd62428,17'd62429,17'd49601,17'd3691,17'd62430,17'd3543,17'd36038,17'd62431,17'd62315,17'd59893,17'd36594,17'd62432,17'd50921,17'd62317,17'd3367,17'd3367,17'd3367,17'd46990,17'd38576,17'd62433,17'd62434,17'd62435,17'd62436,17'd62437,17'd55878,17'd56541,17'd62438,17'd62439,17'd58376,17'd62440,17'd62441,17'd62442,17'd62443,17'd451,17'd794,17'd4084,17'd2409,17'd12496,17'd2098,17'd14178,17'd2098,17'd779,17'd1383,17'd15233,17'd15233,17'd2560,17'd1949,17'd26228,17'd26228,17'd26228,17'd27580,17'd27708,17'd29170,17'd29170,17'd29170,17'd29612,17'd35487,17'd7537,17'd6258,17'd13933,17'd13933,17'd13420,17'd38072,17'd14060,17'd14060,17'd43596,17'd62444,17'd62445,17'd62446,17'd62447,17'd62448,17'd62449,17'd62450,17'd62451,17'd62452,17'd8480,17'd54324,17'd41476,17'd54513,17'd62453,17'd2360,17'd62454,17'd62074,17'd62455,17'd62456,17'd54684,17'd62457
},
'{
17'd16501,17'd10924,17'd10669,17'd3593,17'd10802,17'd10802,17'd10924,17'd10802,17'd52621,17'd2597,17'd17,17'd1128,17'd11,17'd10,17'd979,17'd19,17'd3905,17'd18,17'd16,17'd16,17'd16,17'd17,17'd17,17'd1416,17'd1414,17'd10268,17'd2592,17'd2934,17'd3592,17'd15877,17'd5511,17'd15877,17'd10670,17'd10547,17'd2258,17'd2258,17'd3429,17'd3593,17'd10925,17'd59133,17'd52704,17'd5511,17'd4086,17'd13944,17'd813,17'd15362,17'd58505,17'd60278,17'd59913,17'd59001,17'd60039,17'd56672,17'd57622,17'd1430,17'd56795,17'd1429,17'd69,17'd1981,17'd484,17'd485,17'd60894,17'd838,17'd61167,17'd61167,17'd62458,17'd62459,17'd62460,17'd54787,17'd62461,17'd62462,17'd62463,17'd62464,17'd62465,17'd61689,17'd62466,17'd3775,17'd62467,17'd62468,17'd61564,17'd47092,17'd16412,17'd6622,17'd61299,17'd62469,17'd3780,17'd5999,17'd44863,17'd44863,17'd7091,17'd5839,17'd3470,17'd5999,17'd62470,17'd5412,17'd62226,17'd2981,17'd62471,17'd3478,17'd2644,17'd62472,17'd56694,17'd61702,17'd62473,17'd58042,17'd57396,17'd61189,17'd60656,17'd55282,17'd58159,17'd62474,17'd57274,17'd59647,17'd60052,17'd57778,17'd62475,17'd59024,17'd60427,17'd58661,17'd62476,17'd62477,17'd60920,17'd60059,17'd58042,17'd55778,17'd59655,17'd59144,17'd56459,17'd62478,17'd62479,17'd59286,17'd62480,17'd4636,17'd62481,17'd62482,17'd62483,17'd62484,17'd62485,17'd62486,17'd60936,17'd62487,17'd62488,17'd62489,17'd62490,17'd62491,17'd62492,17'd62493,17'd62494,17'd62495,17'd62496,17'd62497,17'd62498,17'd62499,17'd62251,17'd62500,17'd62501,17'd62502,17'd62253,17'd62503,17'd61870,17'd62504,17'd62505,17'd62506,17'd62507,17'd62508,17'd62509,17'd62510,17'd62509,17'd62136,17'd61610,17'd61877,17'd61094,17'd60087,17'd59429,17'd62511,17'd62512,17'd62513,17'd21665,17'd14924,17'd12410,17'd12417,17'd12109,17'd12110,17'd12419,17'd11958,17'd11959,17'd19920,17'd13885,17'd29331,17'd29341,17'd10852,17'd10479,17'd23679,17'd9045,17'd8569,17'd22473,17'd8731,17'd8575,17'd8577,17'd21987,17'd25147,17'd13257,17'd23343,17'd16072,17'd12120,17'd15694,17'd9890,17'd24216,17'd12428,17'd8258,17'd24714,17'd16567,17'd10747,17'd17018,17'd62514,17'd25683,17'd14939,17'd8740,17'd62143,17'd11536,17'd23526,17'd14394,17'd54045,17'd15573,17'd18921,17'd7790,17'd14932,17'd7953,17'd8421,17'd9622,17'd11968,17'd12726,17'd14140,17'd62515,17'd23875,17'd62516,17'd15311,17'd62517,17'd62518,17'd62519,17'd62520,17'd62521,17'd62522,17'd62523,17'd62524,17'd62525,17'd62526,17'd62527,17'd52163,17'd51075,17'd54751,17'd43155,17'd53563,17'd62400,17'd62157,17'd61498,17'd62528,17'd62529,17'd62530,17'd62283,17'd62531,17'd62532,17'd62533,17'd62534,17'd34298,17'd23736,17'd23736,17'd24421,17'd24421,17'd31341,17'd31341,17'd62535,17'd62536,17'd30579,17'd30579,17'd38806,17'd23736,17'd23736,17'd23567,17'd37511,17'd29974,17'd22501,17'd30277,17'd22329,17'd22331,17'd30276,17'd22506,17'd22162,17'd30580,17'd32497,17'd32660,17'd31656,17'd29973,17'd29099,17'd33482,17'd40964,17'd33793,17'd28851,17'd29688,17'd38978,17'd48987,17'd32668,17'd25438,17'd27765,17'd27766,17'd25833,17'd25708,17'd28600,17'd31034,17'd38667,17'd33802,17'd34113,17'd33793,17'd62537,17'd33182,17'd62538,17'd38546,17'd62539,17'd37394,17'd36275,17'd26911,17'd26669,17'd29123,17'd28387,17'd30450,17'd24438,17'd22703,17'd62540,17'd62541,17'd62542,17'd62543,17'd62544,17'd62545,17'd62546,17'd62547,17'd27279,17'd62548,17'd23238,17'd62549,17'd21559,17'd62550,17'd62551,17'd62552,17'd29714,17'd62553,17'd48064,17'd19969,17'd42906,17'd62554,17'd33983,17'd62555,17'd22224,17'd62556,17'd23623,17'd24304,17'd30793,17'd24305,17'd30793,17'd22758,17'd24794,17'd22935,17'd24479,17'd26217,17'd4993,17'd5150,17'd4841,17'd4686,17'd4689,17'd41459,17'd34657,17'd4526,17'd4846,17'd5162,17'd5011,17'd5011,17'd37944,17'd62557,17'd62558,17'd38444,17'd61928,17'd62559,17'd6071,17'd12168,17'd13415,17'd13567,17'd22256,17'd62560,17'd62561,17'd62561,17'd62562,17'd30034,17'd62563,17'd62185,17'd5176,17'd61272,17'd62055,17'd49601,17'd3691,17'd61396,17'd60504,17'd58732,17'd58733,17'd58733,17'd58732,17'd61661,17'd3366,17'd62318,17'd62564,17'd62565,17'd21620,17'd62566,17'd62567,17'd62568,17'd62569,17'd61665,17'd62570,17'd54870,17'd56097,17'd55266,17'd62438,17'd62571,17'd30644,17'd58013,17'd62572,17'd62573,17'd19361,17'd1665,17'd7850,17'd1823,17'd6868,17'd2393,17'd14178,17'd14178,17'd2575,17'd2575,17'd1383,17'd1383,17'd15233,17'd2394,17'd2560,17'd1949,17'd26228,17'd26228,17'd27708,17'd27708,17'd29170,17'd29170,17'd29170,17'd29170,17'd29611,17'd33051,17'd8507,17'd4868,17'd4867,17'd38072,17'd12636,17'd12636,17'd13176,17'd13176,17'd16855,17'd16132,17'd62574,17'd62575,17'd15348,17'd17291,17'd62449,17'd62576,17'd14309,17'd11865,17'd46883,17'd51760,17'd61674,17'd40858,17'd2079,17'd60632,17'd56213,17'd62577,17'd62455,17'd62456,17'd60517,17'd62578
},
'{
17'd16501,17'd10924,17'd10669,17'd3593,17'd10802,17'd10802,17'd10924,17'd10802,17'd10669,17'd2597,17'd17,17'd18,17'd11,17'd10,17'd979,17'd19,17'd3905,17'd17,17'd16,17'd16,17'd16,17'd17,17'd17,17'd1414,17'd2596,17'd2596,17'd3250,17'd2935,17'd3428,17'd15877,17'd5511,17'd15877,17'd10925,17'd10669,17'd3429,17'd2258,17'd3429,17'd3593,17'd10924,17'd16011,17'd52704,17'd5511,17'd4086,17'd13943,17'd13944,17'd59381,17'd62579,17'd60404,17'd60037,17'd59251,17'd59627,17'd60039,17'd62580,17'd62581,17'd57005,17'd1429,17'd70,17'd1981,17'd484,17'd1980,17'd485,17'd61037,17'd61167,17'd62582,17'd62583,17'd62584,17'd62460,17'd1144,17'd62585,17'd61419,17'd62586,17'd62587,17'd62588,17'd61689,17'd62466,17'd62589,17'd62350,17'd62590,17'd61957,17'd62089,17'd17323,17'd14476,17'd61693,17'd4921,17'd59643,17'd3470,17'd6151,17'd62591,17'd7257,17'd5839,17'd5839,17'd6316,17'd6308,17'd6007,17'd53371,17'd2982,17'd3141,17'd3635,17'd3292,17'd61183,17'd62592,17'd61440,17'd58892,17'd62593,17'd57279,17'd58886,17'd62594,17'd62595,17'd55582,17'd56239,17'd58768,17'd58888,17'd59647,17'd61063,17'd59274,17'd58524,17'd60176,17'd57644,17'd62596,17'd62597,17'd1035,17'd61578,17'd55911,17'd59017,17'd58409,17'd57022,17'd61449,17'd59937,17'd62598,17'd62599,17'd62600,17'd2173,17'd62114,17'd62601,17'd62602,17'd62603,17'd62604,17'd62605,17'd61433,17'd62606,17'd62607,17'd62608,17'd62609,17'd62610,17'd62611,17'd62612,17'd62613,17'd62614,17'd62615,17'd62616,17'd62617,17'd62499,17'd62251,17'd62618,17'd62619,17'd62620,17'd62253,17'd62621,17'd62622,17'd62623,17'd62624,17'd62625,17'd62626,17'd62627,17'd62509,17'd62510,17'd62257,17'd62136,17'd61610,17'd61345,17'd61742,17'd62139,17'd62628,17'd62629,17'd62630,17'd62631,17'd15556,17'd62632,17'd62262,17'd12856,17'd12110,17'd12577,17'd12111,17'd13135,17'd21361,17'd16325,17'd13885,17'd43219,17'd42810,17'd10852,17'd12863,17'd23853,17'd15297,17'd8728,17'd8575,17'd8575,17'd8576,17'd24862,17'd25147,17'd24713,17'd8579,17'd50418,17'd25288,17'd7787,17'd10341,17'd12428,17'd13767,17'd16335,17'd22135,17'd24714,17'd14938,17'd14938,17'd17018,17'd24553,17'd62633,17'd17732,17'd23348,17'd62634,17'd21676,17'd8740,17'd13142,17'd10997,17'd14009,17'd15439,17'd15439,17'd12266,17'd7954,17'd7953,17'd17238,17'd25152,17'd21210,17'd59844,17'd62635,17'd62636,17'd62637,17'd62638,17'd62639,17'd62640,17'd62641,17'd62642,17'd62643,17'd62644,17'd62645,17'd62646,17'd62647,17'd61768,17'd62527,17'd55045,17'd51075,17'd54291,17'd53262,17'd50068,17'd62400,17'd62157,17'd55626,17'd62648,17'd62649,17'd62650,17'd62651,17'd62531,17'd62652,17'd62653,17'd53330,17'd33673,17'd29376,17'd23733,17'd29528,17'd33950,17'd33794,17'd31190,17'd62654,17'd62654,17'd24421,17'd31502,17'd24421,17'd35865,17'd23387,17'd23388,17'd32008,17'd36543,17'd22501,17'd22329,17'd33311,17'd22681,17'd22159,17'd22507,17'd30727,17'd23040,17'd30580,17'd22857,17'd29973,17'd29242,17'd35159,17'd33653,17'd29533,17'd24742,17'd34883,17'd62655,17'd62656,17'd34459,17'd32353,17'd29101,17'd28723,17'd25708,17'd25708,17'd28723,17'd25317,17'd29103,17'd33653,17'd54061,17'd33802,17'd59090,17'd59213,17'd29701,17'd60364,17'd36134,17'd33325,17'd30603,17'd31201,17'd27268,17'd26192,17'd62657,17'd62658,17'd29847,17'd35031,17'd23586,17'd62659,17'd62660,17'd62661,17'd62662,17'd62544,17'd62663,17'd62664,17'd62665,17'd62666,17'd62667,17'd62668,17'd62669,17'd62670,17'd62671,17'd62672,17'd62673,17'd62674,17'd62675,17'd62676,17'd21755,17'd62677,17'd42025,17'd62678,17'd62679,17'd22566,17'd62680,17'd62681,17'd55060,17'd30793,17'd22933,17'd30793,17'd22758,17'd24794,17'd22935,17'd9906,17'd60138,17'd5150,17'd5150,17'd4841,17'd4687,17'd4689,17'd5154,17'd5154,17'd4684,17'd4848,17'd5161,17'd5011,17'd5011,17'd37944,17'd62557,17'd61928,17'd38444,17'd61791,17'd36173,17'd62682,17'd27938,17'd18378,17'd18137,17'd13288,17'd62560,17'd62561,17'd62561,17'd62562,17'd62683,17'd30184,17'd62684,17'd62685,17'd62428,17'd62686,17'd21938,17'd3691,17'd61660,17'd60504,17'd49004,17'd62687,17'd3690,17'd60266,17'd50179,17'd3367,17'd62688,17'd62689,17'd62690,17'd62691,17'd62692,17'd53285,17'd53431,17'd56421,17'd62693,17'd54969,17'd62694,17'd53865,17'd60027,17'd60882,17'd62695,17'd61153,17'd62326,17'd59243,17'd2732,17'd62696,17'd52462,17'd1962,17'd604,17'd12496,17'd2098,17'd2098,17'd14178,17'd2575,17'd2575,17'd413,17'd1383,17'd15233,17'd2394,17'd1950,17'd26228,17'd27580,17'd27580,17'd27708,17'd29170,17'd29170,17'd28793,17'd28793,17'd60625,17'd36903,17'd7705,17'd6258,17'd39328,17'd38203,17'd38072,17'd12636,17'd12636,17'd13176,17'd16855,17'd16132,17'd62697,17'd62698,17'd62699,17'd16959,17'd62700,17'd62701,17'd17415,17'd62702,17'd11441,17'd62703,17'd41905,17'd62704,17'd2539,17'd54873,17'd62705,17'd62706,17'd62577,17'd62707,17'd62456,17'd60517,17'd62708
},
'{
17'd16011,17'd11609,17'd10802,17'd3429,17'd52621,17'd12195,17'd10670,17'd10802,17'd10802,17'd3429,17'd1415,17'd18,17'd2423,17'd1275,17'd4732,17'd283,17'd0,17'd466,17'd17,17'd1277,17'd3905,17'd3905,17'd16,17'd17,17'd1414,17'd2596,17'd2781,17'd2935,17'd3427,17'd15877,17'd5511,17'd15877,17'd11609,17'd3593,17'd3429,17'd2426,17'd2258,17'd3429,17'd10670,17'd16501,17'd5511,17'd5511,17'd5204,17'd4086,17'd13944,17'd813,17'd14445,17'd62709,17'd59250,17'd59913,17'd59001,17'd56791,17'd57622,17'd57622,17'd1430,17'd20272,17'd70,17'd62710,17'd14451,17'd1980,17'd18151,17'd838,17'd490,17'd62582,17'd62711,17'd62712,17'd2612,17'd1428,17'd43879,17'd62713,17'd62714,17'd62715,17'd62716,17'd62717,17'd62466,17'd62718,17'd62719,17'd62720,17'd61297,17'd62721,17'd17323,17'd46708,17'd61693,17'd4921,17'd62722,17'd5839,17'd5841,17'd6150,17'd62723,17'd6774,17'd62724,17'd5839,17'd6774,17'd5999,17'd5842,17'd59786,17'd3142,17'd59640,17'd3635,17'd62096,17'd62725,17'd54802,17'd58276,17'd62726,17'd57279,17'd1459,17'd61837,17'd62727,17'd62594,17'd57133,17'd62728,17'd59274,17'd60052,17'd60051,17'd58887,17'd57512,17'd56129,17'd58768,17'd61846,17'd62729,17'd62730,17'd62731,17'd62732,17'd62733,17'd60176,17'd59523,17'd56697,17'd60424,17'd62734,17'd60926,17'd56813,17'd62735,17'd62736,17'd62737,17'd62738,17'd62739,17'd62740,17'd62741,17'd62742,17'd62743,17'd62744,17'd62745,17'd62746,17'd62747,17'd62748,17'd62611,17'd62749,17'd62613,17'd62750,17'd62751,17'd62752,17'd62753,17'd62754,17'd62618,17'd62619,17'd62620,17'd62755,17'd62756,17'd62757,17'd62758,17'd62759,17'd62760,17'd62761,17'd62762,17'd62763,17'd62257,17'd62509,17'd62136,17'd62258,17'd61611,17'd61223,17'd62764,17'd61879,17'd59556,17'd62765,17'd62766,17'd12699,17'd62767,17'd62768,17'd13518,17'd13365,17'd12857,17'd12861,17'd11806,17'd22472,17'd29488,17'd11666,17'd18915,17'd23336,17'd25278,17'd26037,17'd17965,17'd26874,17'd30672,17'd37334,17'd17481,17'd25147,17'd11967,17'd34206,17'd23173,17'd62769,17'd25288,17'd62770,17'd7618,17'd25004,17'd12590,17'd62771,17'd54382,17'd15303,17'd14011,17'd26040,17'd7621,17'd12728,17'd16692,17'd17356,17'd23872,17'd62772,17'd21676,17'd62773,17'd10032,17'd62774,17'd56734,17'd14938,17'd13766,17'd10861,17'd23176,17'd18085,17'd7954,17'd10746,17'd25929,17'd24871,17'd62775,17'd19040,17'd15310,17'd62776,17'd15200,17'd62777,17'd62778,17'd62779,17'd62780,17'd62781,17'd62782,17'd62783,17'd62646,17'd62784,17'd62526,17'd62277,17'd62785,17'd62786,17'd53263,17'd50068,17'd53333,17'd62787,17'd62281,17'd62788,17'd62018,17'd62789,17'd62790,17'd62791,17'd62283,17'd62792,17'd62793,17'd62794,17'd62795,17'd23918,17'd29528,17'd30578,17'd30578,17'd33801,17'd33950,17'd62796,17'd23211,17'd23733,17'd23918,17'd29376,17'd29376,17'd23387,17'd30128,17'd32351,17'd22501,17'd22500,17'd22325,17'd51306,17'd22683,17'd22861,17'd30880,17'd21848,17'd36691,17'd31343,17'd41273,17'd23918,17'd34621,17'd32353,17'd27637,17'd24744,17'd33482,17'd53556,17'd62797,17'd57076,17'd48987,17'd30432,17'd29970,17'd33643,17'd32658,17'd25435,17'd25317,17'd29244,17'd32353,17'd53720,17'd54061,17'd33653,17'd32353,17'd39138,17'd59998,17'd62798,17'd62799,17'd37394,17'd30757,17'd26911,17'd27523,17'd28277,17'd62800,17'd62801,17'd62802,17'd62803,17'd62804,17'd62805,17'd62806,17'd62807,17'd46006,17'd62808,17'd62809,17'd62810,17'd27540,17'd62041,17'd62811,17'd23948,17'd23764,17'd24281,17'd62812,17'd62813,17'd62814,17'd62815,17'd62816,17'd62817,17'd53729,17'd62818,17'd33983,17'd62819,17'd21903,17'd62820,17'd55740,17'd22934,17'd22586,17'd24306,17'd24306,17'd22586,17'd22758,17'd24794,17'd23628,17'd9906,17'd60138,17'd5150,17'd25770,17'd4841,17'd4686,17'd5156,17'd5154,17'd40397,17'd29024,17'd5002,17'd42031,17'd5012,17'd37697,17'd37945,17'd62821,17'd62822,17'd62823,17'd62824,17'd62825,17'd12008,17'd13286,17'd17908,17'd17909,17'd62826,17'd62827,17'd62828,17'd62827,17'd13053,17'd62683,17'd18978,17'd62684,17'd5021,17'd6078,17'd62829,17'd62830,17'd61017,17'd61145,17'd60266,17'd60267,17'd60022,17'd60022,17'd61145,17'd62831,17'd62832,17'd62833,17'd62834,17'd62835,17'd62836,17'd59610,17'd59237,17'd62837,17'd62838,17'd62839,17'd62840,17'd62841,17'd62842,17'd60027,17'd55470,17'd59249,17'd58630,17'd62066,17'd62843,17'd62844,17'd55882,17'd1944,17'd1680,17'd11062,17'd12496,17'd16256,17'd2098,17'd5940,17'd7027,17'd2575,17'd2589,17'd2589,17'd12644,17'd2394,17'd1950,17'd27580,17'd27580,17'd27581,17'd29170,17'd28793,17'd28793,17'd28793,17'd60625,17'd60625,17'd35487,17'd7537,17'd6095,17'd38459,17'd38072,17'd12483,17'd12483,17'd62845,17'd13176,17'd16855,17'd62846,17'd62847,17'd62848,17'd62849,17'd62850,17'd62851,17'd62852,17'd62853,17'd62854,17'd62855,17'd45787,17'd5024,17'd62856,17'd51182,17'd54085,17'd62857,17'd62858,17'd62859,17'd62707,17'd62455,17'd24492,17'd58253
},
'{
17'd16011,17'd11609,17'd10802,17'd3429,17'd52621,17'd10547,17'd10670,17'd10802,17'd10670,17'd52621,17'd1414,17'd17,17'd13,17'd3,17'd283,17'd1,17'd1830,17'd14,17'd16,17'd1277,17'd18,17'd18,17'd16,17'd1416,17'd1414,17'd2596,17'd2781,17'd2422,17'd3251,17'd15358,17'd5511,17'd52704,17'd15496,17'd11071,17'd3429,17'd2426,17'd2258,17'd3429,17'd10802,17'd11888,17'd5511,17'd5511,17'd5204,17'd4086,17'd13945,17'd13944,17'd59773,17'd62860,17'd60278,17'd60037,17'd59251,17'd59001,17'd56791,17'd57622,17'd57005,17'd20272,17'd69,17'd62710,17'd14451,17'd1980,17'd62861,17'd60894,17'd490,17'd62582,17'd62862,17'd62863,17'd1144,17'd3266,17'd32886,17'd62864,17'd62865,17'd62866,17'd62867,17'd62868,17'd62348,17'd62466,17'd62869,17'd62870,17'd61957,17'd62721,17'd15388,17'd62871,17'd61958,17'd62872,17'd62873,17'd3781,17'd5841,17'd6472,17'd62874,17'd62874,17'd6936,17'd3626,17'd3626,17'd6774,17'd5840,17'd2986,17'd2988,17'd60418,17'd62875,17'd3478,17'd54620,17'd60298,17'd62876,17'd58653,17'd62473,17'd58277,17'd61970,17'd62877,17'd62727,17'd61440,17'd62103,17'd56810,17'd58038,17'd59147,17'd60302,17'd59393,17'd56129,17'd62878,17'd62879,17'd61578,17'd62360,17'd62880,17'd59657,17'd59651,17'd59018,17'd56810,17'd58893,17'd61449,17'd61846,17'd62881,17'd57281,17'd62882,17'd1467,17'd4637,17'd62883,17'd62884,17'd62885,17'd62886,17'd58781,17'd62887,17'd62888,17'd62889,17'd62890,17'd62891,17'd62892,17'd62893,17'd62894,17'd62895,17'd62896,17'd62897,17'd62898,17'd62899,17'd62376,17'd62251,17'd62619,17'd62620,17'd62755,17'd62900,17'd62901,17'd62622,17'd62902,17'd62903,17'd62904,17'd62905,17'd62256,17'd62257,17'd62509,17'd62136,17'd62258,17'd61611,17'd61877,17'd62906,17'd62907,17'd59429,17'd59432,17'd62908,17'd59185,17'd62909,17'd62910,17'd32603,17'd13365,17'd12420,17'd12861,17'd11667,17'd24858,17'd24363,17'd11667,17'd29331,17'd43363,17'd25278,17'd20610,17'd16561,17'd26874,17'd12723,17'd8414,17'd14135,17'd25147,17'd26261,17'd62911,17'd53478,17'd53836,17'd7787,17'd42228,17'd38903,17'd13893,17'd15436,17'd62912,17'd62913,17'd19536,17'd14011,17'd8258,17'd10342,17'd14266,17'd12592,17'd10483,17'd13008,17'd62914,17'd7798,17'd9625,17'd62915,17'd16449,17'd14678,17'd10996,17'd12727,17'd14682,17'd12727,17'd25004,17'd10609,17'd14932,17'd13377,17'd62916,17'd62917,17'd62918,17'd11972,17'd62919,17'd15312,17'd62920,17'd62921,17'd62922,17'd62923,17'd62924,17'd62925,17'd62926,17'd62927,17'd62928,17'd61768,17'd62277,17'd62929,17'd51474,17'd51828,17'd52817,17'd53333,17'd62787,17'd62281,17'd62930,17'd62931,17'd62932,17'd62933,17'd62933,17'd62789,17'd62934,17'd62935,17'd62936,17'd54057,17'd23918,17'd31033,17'd29375,17'd30424,17'd30424,17'd33801,17'd44244,17'd23209,17'd23733,17'd31502,17'd29530,17'd23388,17'd30128,17'd32351,17'd30277,17'd22328,17'd22680,17'd32344,17'd22507,17'd35153,17'd22156,17'd22163,17'd30727,17'd22159,17'd22328,17'd23734,17'd50364,17'd32668,17'd25178,17'd24898,17'd28851,17'd38978,17'd57839,17'd62797,17'd33644,17'd40964,17'd31034,17'd43977,17'd28721,17'd42749,17'd29101,17'd31034,17'd33483,17'd53720,17'd53720,17'd33653,17'd33483,17'd59457,17'd59341,17'd32681,17'd38824,17'd62937,17'd35027,17'd29990,17'd27034,17'd26912,17'd62938,17'd62939,17'd32035,17'd62940,17'd62941,17'd22185,17'd62942,17'd62943,17'd21095,17'd46006,17'd62944,17'd61132,17'd24926,17'd62945,17'd62946,17'd62947,17'd23415,17'd62948,17'd62949,17'd62950,17'd62951,17'd62952,17'd62953,17'd62954,17'd21446,17'd62955,17'd62956,17'd33983,17'd62957,17'd23271,17'd23103,17'd54593,17'd22758,17'd26111,17'd62958,17'd24643,17'd22758,17'd25878,17'd22759,17'd62423,17'd24650,17'd26827,17'd5478,17'd25770,17'd4686,17'd4686,17'd4526,17'd28778,17'd4685,17'd4848,17'd5329,17'd42031,17'd5012,17'd37697,17'd62557,17'd62959,17'd62960,17'd62823,17'd62961,17'd10781,17'd12628,17'd28781,17'd18265,17'd27431,17'd62826,17'd62827,17'd62828,17'd62827,17'd13053,17'd62683,17'd18978,17'd11439,17'd19097,17'd5176,17'd62962,17'd62963,17'd21938,17'd3691,17'd20392,17'd60267,17'd3544,17'd20392,17'd60753,17'd21460,17'd62964,17'd49300,17'd62965,17'd3368,17'd21462,17'd47854,17'd42643,17'd60271,17'd62966,17'd62967,17'd55262,17'd62968,17'd53865,17'd53740,17'd56212,17'd2070,17'd53433,17'd57885,17'd59495,17'd19997,17'd6083,17'd3745,17'd445,17'd12026,17'd16382,17'd16256,17'd6889,17'd5940,17'd412,17'd412,17'd413,17'd413,17'd15233,17'd28916,17'd26966,17'd26228,17'd27581,17'd27581,17'd29170,17'd28793,17'd28793,17'd28793,17'd60625,17'd36904,17'd9261,17'd6418,17'd38459,17'd38203,17'd38580,17'd12483,17'd12483,17'd12913,17'd16855,17'd15735,17'd62847,17'd62969,17'd62849,17'd62970,17'd62971,17'd62972,17'd62973,17'd62974,17'd62975,17'd62976,17'd62977,17'd7680,17'd62978,17'd54323,17'd37302,17'd55359,17'd62858,17'd62979,17'd62980,17'd53218,17'd24492,17'd58253
},
'{
17'd16501,17'd11609,17'd3101,17'd3252,17'd3252,17'd14070,17'd3251,17'd2934,17'd2934,17'd2935,17'd1689,17'd14,17'd2,17'd1,17'd4884,17'd3749,17'd62981,17'd1830,17'd0,17'd0,17'd18,17'd18,17'd16,17'd1416,17'd1414,17'd1414,17'd1689,17'd2422,17'd3101,17'd15358,17'd4891,17'd52704,17'd5511,17'd3751,17'd10669,17'd12194,17'd2258,17'd2258,17'd10669,17'd10925,17'd15877,17'd5204,17'd5204,17'd4086,17'd12653,17'd13945,17'd473,17'd62982,17'd62983,17'd59250,17'd59498,17'd58256,17'd62984,17'd57003,17'd56795,17'd20272,17'd62985,17'd19500,17'd14451,17'd1980,17'd62341,17'd62458,17'd61037,17'd838,17'd67,17'd18151,17'd2950,17'd32731,17'd54608,17'd62986,17'd62987,17'd62714,17'd62988,17'd62989,17'd62717,17'd62990,17'd62991,17'd62992,17'd62993,17'd62994,17'd62089,17'd15141,17'd62995,17'd62996,17'd62997,17'd62998,17'd5839,17'd5841,17'd6151,17'd6775,17'd6477,17'd62999,17'd6471,17'd6471,17'd3781,17'd3297,17'd63000,17'd3141,17'd4771,17'd3789,17'd59141,17'd63001,17'd58401,17'd55906,17'd61968,17'd61058,17'd61704,17'd60915,17'd62877,17'd61440,17'd58159,17'd63002,17'd62475,17'd59933,17'd55905,17'd57391,17'd63003,17'd56350,17'd63004,17'd57644,17'd63005,17'd63006,17'd63007,17'd59399,17'd60923,17'd58651,17'd60176,17'd62475,17'd61449,17'd63008,17'd63009,17'd63010,17'd62735,17'd63011,17'd63012,17'd63013,17'd63014,17'd63015,17'd63016,17'd63017,17'd61433,17'd63018,17'd63019,17'd61985,17'd63020,17'd63021,17'd63022,17'd62894,17'd63023,17'd63024,17'd63025,17'd63026,17'd63027,17'd62251,17'd62619,17'd63028,17'd63029,17'd62900,17'd62901,17'd63030,17'd63031,17'd63032,17'd63033,17'd63034,17'd62627,17'd62381,17'd62257,17'd62136,17'd63035,17'd61474,17'd61611,17'd63036,17'd63037,17'd60700,17'd63038,17'd63039,17'd57308,17'd63040,17'd56269,17'd63041,17'd30684,17'd12420,17'd12861,17'd11807,17'd25143,17'd24706,17'd11667,17'd29331,17'd32590,17'd10852,17'd11524,17'd12585,17'd8883,17'd15568,17'd9349,17'd17126,17'd24213,17'd11405,17'd61750,17'd23174,17'd13140,17'd16565,17'd63042,17'd63043,17'd7293,17'd21059,17'd24870,17'd61618,17'd21059,17'd7621,17'd7621,17'd13769,17'd14678,17'd54045,17'd18810,17'd18691,17'd63044,17'd63044,17'd11143,17'd63045,17'd20616,17'd13378,17'd14269,17'd18921,17'd15572,17'd16567,17'd13007,17'd25004,17'd7790,17'd14679,17'd53039,17'd55950,17'd63046,17'd12125,17'd63047,17'd10870,17'd63048,17'd63049,17'd63050,17'd63051,17'd63052,17'd63053,17'd63054,17'd63055,17'd63056,17'd58457,17'd59332,17'd63057,17'd51154,17'd52426,17'd53333,17'd61114,17'd51736,17'd51308,17'd63058,17'd62022,17'd63059,17'd63060,17'd63061,17'd63062,17'd63063,17'd63064,17'd63065,17'd63066,17'd29241,17'd24086,17'd23731,17'd24087,17'd32186,17'd24087,17'd23732,17'd31502,17'd23567,17'd29974,17'd22501,17'd36986,17'd32827,17'd32827,17'd23572,17'd35158,17'd34107,17'd46958,17'd32660,17'd37659,17'd31657,17'd35429,17'd22677,17'd23389,17'd23733,17'd34621,17'd33802,17'd25031,17'd24745,17'd28851,17'd30733,17'd33644,17'd62656,17'd50364,17'd48987,17'd33653,17'd42148,17'd43977,17'd43977,17'd39591,17'd30432,17'd38667,17'd54061,17'd59863,17'd54061,17'd33483,17'd41730,17'd29970,17'd63067,17'd63068,17'd63069,17'd37663,17'd30592,17'd30747,17'd31042,17'd29395,17'd63070,17'd63071,17'd26798,17'd63072,17'd63073,17'd22030,17'd63074,17'd63075,17'd20941,17'd63076,17'd63077,17'd63078,17'd63079,17'd63080,17'd63081,17'd63082,17'd23762,17'd63083,17'd63084,17'd62813,17'd63085,17'd19055,17'd20215,17'd19335,17'd21915,17'd63086,17'd62048,17'd61923,17'd21749,17'd30791,17'd57588,17'd53577,17'd22586,17'd25767,17'd60137,17'd24643,17'd23110,17'd23110,17'd7658,17'd7324,17'd24649,17'd4994,17'd4687,17'd4686,17'd5157,17'd4846,17'd40397,17'd34791,17'd29024,17'd5009,17'd5166,17'd5167,17'd37697,17'd52603,17'd62821,17'd62823,17'd63087,17'd62824,17'd7185,17'd12474,17'd18747,17'd16378,17'd18748,17'd14057,17'd13568,17'd63088,17'd63088,17'd63088,17'd63089,17'd12910,17'd63090,17'd11439,17'd62684,17'd4215,17'd61796,17'd62314,17'd62830,17'd60753,17'd3545,17'd60753,17'd63091,17'd60392,17'd60392,17'd63092,17'd63093,17'd62830,17'd62965,17'd63094,17'd63095,17'd2879,17'd63096,17'd63097,17'd63098,17'd63099,17'd55752,17'd63100,17'd63101,17'd63102,17'd56322,17'd58872,17'd53144,17'd56780,17'd63103,17'd18757,17'd8314,17'd5629,17'd3391,17'd5630,17'd4714,17'd4714,17'd6889,17'd5630,17'd2409,17'd412,17'd413,17'd1383,17'd2394,17'd29169,17'd27707,17'd27707,17'd27708,17'd29170,17'd29170,17'd28793,17'd60625,17'd60625,17'd31251,17'd36904,17'd7705,17'd6258,17'd4867,17'd38203,17'd38580,17'd44019,17'd12913,17'd13572,17'd15104,17'd62846,17'd63104,17'd63105,17'd63106,17'd63107,17'd62972,17'd63108,17'd63109,17'd63109,17'd63110,17'd17543,17'd63111,17'd46021,17'd63112,17'd53516,17'd63113,17'd53061,17'd63114,17'd63115,17'd62980,17'd53218,17'd2072,17'd57756
},
'{
17'd16501,17'd16501,17'd3251,17'd3252,17'd3252,17'd3101,17'd2934,17'd2593,17'd2782,17'd6424,17'd9815,17'd63116,17'd1830,17'd3749,17'd14069,17'd14069,17'd63117,17'd63118,17'd1830,17'd0,17'd18,17'd19,17'd16,17'd22965,17'd1414,17'd1414,17'd1689,17'd1688,17'd3252,17'd3428,17'd4891,17'd5646,17'd5511,17'd3592,17'd10802,17'd10547,17'd2426,17'd2258,17'd10669,17'd10924,17'd5204,17'd5204,17'd5204,17'd5204,17'd12504,17'd12653,17'd16392,17'd59773,17'd60519,17'd63119,17'd60037,17'd59498,17'd63120,17'd56559,17'd56223,17'd20272,17'd55892,17'd62985,17'd62710,17'd1980,17'd62341,17'd62341,17'd62210,17'd1291,17'd68,17'd485,17'd998,17'd32886,17'd54693,17'd63121,17'd63122,17'd63123,17'd63124,17'd63125,17'd63126,17'd62990,17'd62991,17'd63127,17'd63128,17'd63129,17'd62089,17'd63130,17'd63131,17'd63132,17'd63133,17'd63134,17'd3781,17'd5841,17'd5841,17'd6318,17'd63135,17'd63136,17'd3949,17'd6772,17'd62998,17'd63137,17'd63138,17'd3624,17'd3299,17'd5257,17'd63139,17'd60652,17'd63140,17'd63141,17'd63142,17'd58772,17'd63143,17'd63144,17'd56353,17'd55779,17'd60657,17'd56132,17'd57517,17'd59523,17'd57131,17'd57391,17'd63145,17'd63146,17'd62726,17'd58042,17'd59651,17'd59283,17'd62357,17'd63147,17'd63148,17'd59400,17'd59018,17'd59024,17'd56697,17'd57644,17'd60794,17'd63149,17'd63150,17'd63151,17'd63152,17'd63153,17'd62884,17'd63154,17'd62238,17'd63155,17'd61718,17'd63156,17'd63157,17'd63158,17'd63159,17'd63160,17'd62892,17'd63161,17'd63162,17'd63163,17'd63164,17'd63165,17'd63166,17'd62250,17'd63167,17'd63028,17'd63029,17'd63168,17'd63169,17'd62901,17'd62622,17'd63170,17'd63171,17'd63172,17'd62627,17'd62256,17'd62381,17'd62509,17'd63173,17'd63035,17'd61611,17'd63174,17'd63175,17'd63176,17'd60217,17'd61744,17'd57946,17'd15171,17'd63177,17'd58075,17'd32603,17'd12106,17'd11962,17'd13762,17'd23169,17'd36348,17'd11521,17'd11666,17'd32590,17'd10988,17'd11399,17'd16200,17'd10175,17'd11404,17'd12865,17'd8417,17'd8580,17'd11674,17'd63178,17'd63179,17'd63180,17'd63181,17'd63182,17'd63183,17'd18086,17'd10342,17'd15442,17'd20613,17'd15442,17'd14391,17'd8259,17'd14141,17'd22478,17'd7627,17'd17854,17'd55218,17'd61101,17'd23526,17'd63184,17'd63185,17'd10997,17'd13378,17'd17018,17'd19646,17'd63186,17'd24716,17'd23867,17'd62387,17'd15191,17'd22138,17'd20182,17'd63187,17'd16698,17'd63188,17'd13144,17'd16456,17'd63189,17'd63190,17'd63191,17'd63192,17'd63193,17'd63194,17'd63195,17'd63055,17'd63196,17'd63197,17'd59332,17'd63198,17'd53986,17'd52426,17'd52817,17'd61114,17'd51736,17'd53986,17'd63199,17'd63200,17'd62528,17'd63201,17'd63202,17'd63203,17'd63062,17'd63204,17'd63205,17'd63206,17'd55228,17'd31033,17'd23732,17'd24086,17'd24087,17'd31033,17'd30275,17'd29376,17'd29974,17'd22328,17'd22680,17'd22332,17'd22332,17'd22677,17'd33795,17'd33795,17'd40523,17'd34107,17'd30427,17'd39911,17'd35018,17'd36426,17'd30128,17'd34137,17'd28851,17'd29533,17'd29533,17'd28851,17'd35159,17'd38978,17'd50364,17'd50364,17'd48987,17'd34276,17'd32668,17'd38406,17'd42302,17'd43553,17'd41730,17'd33483,17'd40964,17'd34282,17'd63207,17'd59863,17'd53720,17'd33318,17'd29825,17'd59340,17'd63208,17'd63209,17'd41869,17'd37519,17'd30592,17'd30747,17'd31042,17'd35028,17'd63210,17'd62801,17'd25722,17'd63211,17'd23588,17'd22352,17'd29854,17'd63212,17'd63213,17'd63214,17'd63215,17'd63216,17'd63217,17'd63218,17'd63219,17'd63218,17'd63220,17'd63221,17'd63222,17'd63223,17'd63224,17'd63225,17'd21271,17'd20236,17'd28054,17'd34915,17'd60871,17'd21590,17'd63226,17'd22221,17'd23792,17'd22758,17'd22758,17'd63227,17'd62958,17'd26111,17'd24794,17'd23628,17'd6702,17'd7324,17'd24649,17'd5326,17'd4686,17'd4841,17'd5157,17'd4847,17'd34791,17'd4685,17'd5008,17'd5163,17'd5167,17'd5012,17'd5171,17'd36587,17'd63228,17'd62823,17'd63229,17'd63230,17'd11857,17'd13051,17'd25231,17'd15100,17'd18266,17'd63231,17'd63088,17'd63088,17'd13568,17'd13568,17'd63089,17'd63232,17'd63090,17'd11439,17'd62684,17'd63233,17'd63234,17'd62686,17'd62187,17'd49601,17'd49500,17'd3545,17'd20260,17'd21154,17'd7845,17'd7845,17'd62963,17'd3546,17'd62835,17'd63235,17'd35902,17'd63236,17'd60145,17'd63237,17'd63098,17'd63101,17'd58241,17'd58740,17'd63238,17'd63102,17'd62336,17'd63239,17'd63240,17'd57106,17'd37954,17'd9101,17'd5775,17'd11721,17'd4085,17'd5940,17'd5183,17'd4714,17'd3073,17'd5630,17'd2409,17'd2409,17'd413,17'd15233,17'd28916,17'd29169,17'd29610,17'd27708,17'd29170,17'd29170,17'd29170,17'd28793,17'd60625,17'd60625,17'd31251,17'd36903,17'd8507,17'd37959,17'd38203,17'd38203,17'd38580,17'd44019,17'd12913,17'd14584,17'd62846,17'd62847,17'd63241,17'd63242,17'd63107,17'd63243,17'd63108,17'd63244,17'd63245,17'd63246,17'd63247,17'd63248,17'd62203,17'd63249,17'd63250,17'd62704,17'd63251,17'd63252,17'd63253,17'd63115,17'd35484,17'd53218,17'd2070,17'd57756
},
'{
17'd13943,17'd3592,17'd3251,17'd2935,17'd3252,17'd3101,17'd2934,17'd63254,17'd63255,17'd11454,17'd63256,17'd63257,17'd12929,17'd63117,17'd63258,17'd14867,17'd63259,17'd63260,17'd1830,17'd2,17'd18,17'd19,17'd17,17'd1416,17'd1414,17'd1414,17'd1127,17'd1688,17'd3252,17'd3251,17'd3902,17'd5646,17'd5203,17'd4086,17'd10670,17'd12194,17'd57493,17'd2426,17'd52621,17'd10925,17'd5204,17'd5203,17'd5511,17'd5511,17'd3592,17'd12505,17'd11888,17'd15118,17'd63261,17'd62983,17'd63262,17'd63263,17'd58380,17'd56114,17'd56795,17'd20272,17'd55892,17'd62985,17'd19500,17'd305,17'd18391,17'd17791,17'd18151,17'd1981,17'd69,17'd486,17'd1290,17'd63264,17'd62212,17'd63265,17'd63266,17'd63267,17'd63268,17'd63269,17'd63270,17'd62990,17'd62991,17'd63271,17'd63272,17'd61957,17'd63129,17'd63273,17'd63274,17'd63275,17'd61429,17'd60903,17'd62998,17'd6773,17'd6152,17'd5999,17'd6775,17'd62998,17'd6772,17'd3950,17'd60783,17'd62873,17'd63276,17'd3945,17'd53234,17'd3476,17'd5257,17'd53524,17'd60536,17'd60538,17'd63277,17'd55906,17'd58659,17'd58659,17'd61188,17'd56457,17'd55183,17'd63278,17'd57390,17'd57783,17'd63279,17'd63280,17'd63281,17'd58771,17'd58160,17'd58277,17'd62099,17'd59282,17'd61443,17'd63282,17'd58527,17'd60545,17'd63283,17'd59018,17'd61190,17'd57918,17'd59282,17'd63284,17'd63285,17'd57400,17'd63286,17'd63287,17'd63288,17'd63289,17'd63290,17'd63291,17'd63292,17'd63293,17'd63294,17'd53883,17'd63295,17'd63296,17'd63297,17'd63298,17'd63299,17'd63300,17'd63024,17'd63301,17'd62899,17'd62250,17'd63302,17'd63303,17'd63304,17'd63168,17'd63169,17'd63305,17'd63030,17'd61870,17'd63306,17'd62904,17'd62905,17'd62508,17'd62508,17'd63307,17'd63173,17'd63035,17'd61739,17'd61611,17'd61741,17'd60086,17'd60342,17'd63308,17'd62512,17'd63309,17'd63310,17'd63311,17'd52796,17'd15685,17'd12260,17'd13762,17'd21985,17'd18327,17'd13762,17'd11520,17'd11665,17'd10737,17'd12584,17'd63312,17'd57063,17'd25147,17'd8250,17'd14676,17'd10860,17'd15693,17'd53710,17'd63313,17'd16206,17'd8426,17'd63314,17'd63315,17'd9891,17'd21059,17'd21059,17'd22301,17'd14139,17'd12591,17'd8891,17'd11281,17'd7793,17'd54281,17'd8740,17'd54121,17'd21676,17'd63316,17'd63317,17'd17486,17'd63318,17'd14266,17'd14387,17'd15304,17'd63319,17'd63320,17'd7622,17'd7293,17'd55949,17'd19782,17'd63321,17'd57825,17'd62269,17'd14015,17'd11149,17'd63322,17'd63323,17'd63049,17'd63324,17'd63325,17'd63326,17'd63327,17'd63328,17'd63055,17'd63329,17'd63330,17'd62526,17'd57842,17'd51308,17'd53559,17'd54845,17'd61114,17'd51736,17'd50900,17'd56969,17'd63331,17'd63332,17'd63333,17'd63334,17'd63335,17'd63203,17'd63336,17'd63337,17'd57564,17'd50730,17'd29527,17'd23733,17'd23920,17'd29528,17'd29241,17'd23564,17'd29827,17'd30277,17'd22677,17'd35296,17'd31343,17'd36566,17'd36566,17'd34107,17'd23391,17'd45492,17'd35158,17'd31194,17'd35017,17'd32667,17'd30278,17'd24902,17'd28977,17'd32353,17'd30432,17'd28368,17'd34883,17'd62655,17'd62797,17'd50363,17'd34621,17'd34276,17'd29533,17'd33318,17'd42302,17'd42302,17'd53720,17'd38667,17'd33793,17'd34113,17'd50156,17'd34113,17'd59863,17'd63338,17'd43553,17'd43022,17'd28253,17'd27028,17'd37135,17'd63339,17'd63340,17'd35027,17'd27380,17'd31042,17'd30755,17'd63210,17'd63341,17'd24607,17'd63342,17'd63343,17'd63344,17'd63345,17'd63346,17'd20943,17'd63347,17'd25205,17'd63348,17'd63349,17'd62551,17'd63350,17'd22888,17'd23065,17'd24115,17'd23067,17'd63351,17'd63352,17'd18005,17'd19201,17'd63353,17'd53923,17'd22226,17'd63354,17'd23100,17'd22740,17'd22222,17'd22933,17'd11984,17'd24643,17'd57470,17'd25625,17'd54956,17'd61528,17'd22935,17'd7324,17'd24479,17'd5323,17'd24944,17'd32552,17'd4840,17'd5157,17'd4684,17'd61529,17'd38567,17'd5009,17'd37030,17'd5012,17'd5013,17'd36172,17'd63355,17'd63229,17'd62824,17'd62961,17'd7185,17'd17176,17'd15099,17'd63356,17'd63357,17'd63358,17'd17541,17'd63088,17'd13568,17'd63359,17'd63359,17'd63089,17'd63232,17'd63090,17'd11716,17'd29602,17'd62053,17'd63234,17'd63360,17'd62686,17'd62830,17'd7845,17'd63092,17'd7845,17'd62963,17'd62830,17'd62830,17'd3547,17'd63361,17'd63362,17'd63363,17'd63364,17'd63365,17'd63366,17'd63098,17'd63367,17'd58740,17'd63368,17'd59241,17'd58859,17'd59488,17'd53219,17'd63369,17'd58629,17'd19600,17'd57747,17'd1943,17'd63370,17'd2240,17'd4085,17'd5958,17'd4559,17'd3073,17'd5776,17'd8185,17'd2409,17'd412,17'd14178,17'd14586,17'd28916,17'd29037,17'd29892,17'd28793,17'd29170,17'd29039,17'd60625,17'd60625,17'd60625,17'd31251,17'd36903,17'd12923,17'd8186,17'd4883,17'd37709,17'd38203,17'd38580,17'd12635,17'd62444,17'd14584,17'd17180,17'd63371,17'd63372,17'd63373,17'd63243,17'd63374,17'd63375,17'd63376,17'd63246,17'd63377,17'd63378,17'd63379,17'd63380,17'd63381,17'd63382,17'd20262,17'd54513,17'd63383,17'd63253,17'd63115,17'd35484,17'd53218,17'd2070,17'd57757
},
'{
17'd13943,17'd5204,17'd3428,17'd3101,17'd2935,17'd3101,17'd3751,17'd63384,17'd63385,17'd63385,17'd12332,17'd11608,17'd63386,17'd9684,17'd63387,17'd10543,17'd10923,17'd63258,17'd62981,17'd2,17'd3905,17'd18,17'd17,17'd1416,17'd1414,17'd1414,17'd1127,17'd4247,17'd1831,17'd3251,17'd3902,17'd4426,17'd5203,17'd5204,17'd10670,17'd10547,17'd12194,17'd2426,17'd52621,17'd10925,17'd5204,17'd5203,17'd52704,17'd52704,17'd15496,17'd3901,17'd11888,17'd14320,17'd15243,17'd63388,17'd63389,17'd47,17'd63390,17'd56675,17'd56223,17'd20272,17'd55892,17'd55892,17'd62985,17'd15366,17'd18391,17'd17791,17'd995,17'd484,17'd1981,17'd487,17'd1148,17'd39038,17'd1288,17'd62212,17'd61289,17'd63391,17'd63392,17'd63393,17'd63394,17'd63395,17'd62869,17'd63396,17'd63397,17'd63398,17'd63399,17'd62994,17'd63274,17'd63400,17'd6464,17'd63401,17'd63134,17'd6774,17'd5841,17'd3469,17'd63402,17'd62998,17'd6772,17'd3950,17'd4463,17'd4922,17'd4289,17'd53165,17'd3475,17'd3474,17'd3476,17'd3464,17'd53687,17'd60653,17'd56574,17'd63403,17'd63404,17'd63405,17'd55906,17'd56457,17'd55907,17'd63406,17'd63403,17'd55378,17'd57018,17'd61190,17'd56807,17'd57918,17'd58160,17'd58406,17'd57396,17'd56810,17'd63407,17'd63408,17'd61192,17'd63409,17'd60795,17'd59650,17'd62232,17'd58768,17'd59524,17'd59272,17'd63410,17'd63411,17'd63412,17'd63413,17'd4960,17'd63414,17'd63415,17'd63416,17'd63417,17'd63418,17'd63419,17'd63420,17'd51949,17'd63421,17'd63422,17'd63423,17'd63424,17'd63425,17'd63426,17'd63301,17'd62899,17'd63427,17'd63428,17'd63429,17'd63430,17'd63431,17'd63432,17'd63305,17'd63433,17'd62622,17'd63032,17'd63434,17'd63172,17'd62762,17'd63435,17'd63436,17'd63437,17'd63173,17'd62382,17'd63035,17'd63438,17'd62764,17'd63439,17'd61613,17'd63440,17'd61480,17'd22129,17'd63441,17'd63442,17'd12417,17'd12260,17'd13762,17'd14673,17'd11523,17'd11521,17'd13762,17'd15186,17'd10736,17'd12584,17'd63443,17'd63444,17'd18202,17'd57690,17'd63445,17'd63446,17'd63447,17'd8890,17'd21058,17'd25681,17'd62387,17'd14011,17'd26040,17'd16567,17'd19536,17'd14679,17'd17852,17'd15438,17'd63448,17'd24552,17'd63449,17'd11676,17'd54650,17'd63450,17'd21676,17'd25007,17'd63316,17'd63317,17'd17486,17'd17131,17'd14392,17'd22138,17'd53711,17'd63451,17'd15573,17'd9052,17'd63452,17'd23868,17'd24370,17'd55322,17'd63453,17'd12272,17'd63454,17'd63455,17'd63322,17'd63323,17'd63456,17'd63457,17'd63458,17'd63459,17'd63460,17'd63461,17'd63462,17'd63463,17'd63464,17'd61768,17'd63465,17'd50820,17'd52585,17'd54845,17'd55330,17'd63466,17'd50900,17'd58587,17'd63199,17'd63467,17'd63468,17'd63469,17'd63470,17'd63471,17'd63472,17'd50727,17'd58463,17'd63473,17'd58091,17'd31029,17'd23920,17'd23920,17'd23918,17'd29972,17'd29830,17'd39278,17'd31656,17'd22858,17'd22506,17'd39441,17'd39441,17'd48913,17'd30428,17'd44702,17'd45754,17'd23572,17'd30582,17'd38979,17'd29377,17'd24416,17'd32353,17'd30432,17'd25031,17'd30733,17'd56966,17'd57205,17'd57205,17'd62655,17'd34106,17'd29533,17'd32353,17'd39443,17'd38282,17'd38406,17'd32668,17'd38808,17'd34282,17'd52966,17'd57070,17'd49680,17'd59863,17'd53557,17'd43157,17'd32996,17'd35012,17'd63474,17'd28136,17'd63339,17'd63340,17'd36706,17'd32838,17'd26911,17'd30755,17'd63070,17'd34472,17'd22883,17'd24106,17'd63475,17'd26197,17'd31219,17'd63476,17'd20788,17'd30910,17'd63477,17'd63478,17'd63479,17'd63480,17'd63481,17'd22188,17'd23416,17'd63482,17'd23597,17'd63483,17'd63484,17'd19195,17'd63485,17'd63486,17'd63487,17'd63488,17'd23099,17'd23098,17'd22567,17'd23624,17'd63489,17'd61268,17'd62958,17'd60137,17'd25878,17'd26583,17'd11158,17'd26216,17'd24479,17'd7324,17'd4992,17'd5608,17'd4840,17'd4840,17'd4846,17'd40397,17'd61529,17'd38318,17'd5165,17'd51930,17'd37435,17'd5171,17'd63490,17'd63355,17'd63491,17'd62961,17'd63492,17'd12007,17'd63493,17'd15229,17'd63494,17'd63495,17'd63496,17'd63497,17'd17541,17'd63359,17'd18380,17'd63359,17'd63089,17'd63232,17'd30643,17'd30034,17'd29885,17'd62185,17'd63498,17'd62428,17'd63499,17'd61144,17'd7188,17'd7845,17'd63500,17'd62963,17'd62830,17'd63501,17'd3369,17'd63502,17'd52274,17'd63503,17'd63504,17'd60881,17'd63505,17'd55999,17'd63506,17'd63507,17'd63508,17'd58000,17'd57234,17'd53512,17'd63509,17'd52457,17'd23299,17'd2556,17'd37167,17'd1944,17'd4424,17'd12637,17'd4085,17'd5958,17'd4559,17'd5940,17'd49009,17'd49008,17'd2393,17'd2393,17'd16256,17'd14586,17'd28916,17'd27707,17'd29170,17'd28793,17'd29040,17'd29040,17'd60625,17'd60625,17'd60625,17'd31251,17'd35487,17'd7705,17'd6095,17'd4867,17'd38203,17'd38580,17'd12635,17'd13056,17'd62444,17'd15862,17'd63371,17'd62969,17'd63242,17'd63373,17'd63374,17'd63108,17'd63510,17'd63376,17'd63377,17'd63511,17'd63377,17'd63512,17'd17913,17'd63513,17'd4223,17'd45655,17'd63514,17'd33536,17'd2218,17'd63515,17'd23471,17'd53218,17'd2070,17'd57757
},
'{
17'd4737,17'd5511,17'd15358,17'd3101,17'd2935,17'd3251,17'd3751,17'd63384,17'd63516,17'd63516,17'd63517,17'd63518,17'd63519,17'd9814,17'd12783,17'd63520,17'd10543,17'd63521,17'd14319,17'd13,17'd26127,17'd3905,17'd17,17'd1415,17'd1414,17'd1414,17'd466,17'd4247,17'd1831,17'd3101,17'd4244,17'd4087,17'd15117,17'd5511,17'd54978,17'd12194,17'd63522,17'd12194,17'd52621,17'd10924,17'd5204,17'd6730,17'd4425,17'd4425,17'd15496,17'd3751,17'd10924,17'd12504,17'd14746,17'd43,17'd62339,17'd63523,17'd58379,17'd56112,17'd56795,17'd20272,17'd60775,17'd55892,17'd68,17'd15366,17'd1980,17'd17554,17'd2438,17'd995,17'd670,17'd488,17'd672,17'd1843,17'd2437,17'd2437,17'd63524,17'd63525,17'd63526,17'd63527,17'd63528,17'd62218,17'd62869,17'd63529,17'd63530,17'd63531,17'd63532,17'd15012,17'd14627,17'd63533,17'd63534,17'd6303,17'd63535,17'd6477,17'd63536,17'd6308,17'd63537,17'd61301,17'd60783,17'd3950,17'd3951,17'd60290,17'd52625,17'd59390,17'd3947,17'd63538,17'd63539,17'd3476,17'd63540,17'd63541,17'd63542,17'd55780,17'd63543,17'd55582,17'd63404,17'd59013,17'd55907,17'd56689,17'd63544,17'd63545,17'd63546,17'd61441,17'd58893,17'd57022,17'd57648,17'd58406,17'd56909,17'd63547,17'd63548,17'd63407,17'd63549,17'd63147,17'd62105,17'd57518,17'd63550,17'd62232,17'd58893,17'd57644,17'd59397,17'd63551,17'd58412,17'd63552,17'd63553,17'd5894,17'd61851,17'd63554,17'd63555,17'd63556,17'd63557,17'd63558,17'd44863,17'd63559,17'd63560,17'd63561,17'd63562,17'd63563,17'd63163,17'd63165,17'd62753,17'd63564,17'd63565,17'd63428,17'd63566,17'd63567,17'd63432,17'd63568,17'd63569,17'd63168,17'd63570,17'd62760,17'd63571,17'd63435,17'd63572,17'd63573,17'd63307,17'd63437,17'd63437,17'd63173,17'd61610,17'd60573,17'd60699,17'd60575,17'd63574,17'd63575,17'd63576,17'd60097,17'd63577,17'd13134,17'd11958,17'd11807,17'd14931,17'd14931,17'd13762,17'd13516,17'd13362,17'd11395,17'd11400,17'd63578,17'd63579,17'd63580,17'd63581,17'd63582,17'd63583,17'd63584,17'd22480,17'd58569,17'd14140,17'd25681,17'd15436,17'd22475,17'd12590,17'd12428,17'd13893,17'd7621,17'd63448,17'd17130,17'd10482,17'd20616,17'd60708,17'd63585,17'd63586,17'd59841,17'd63587,17'd24051,17'd60350,17'd63588,17'd17853,17'd16692,17'd16693,17'd63589,17'd54829,17'd17130,17'd7791,17'd63590,17'd63591,17'd7959,17'd54121,17'd63592,17'd11539,17'd63593,17'd63594,17'd63595,17'd25011,17'd63596,17'd63597,17'd63598,17'd63599,17'd63600,17'd63601,17'd63602,17'd63603,17'd63604,17'd63605,17'd58094,17'd61363,17'd50069,17'd61114,17'd55330,17'd57071,17'd50900,17'd58587,17'd63606,17'd63607,17'd63608,17'd63609,17'd63610,17'd63611,17'd63612,17'd50894,17'd59721,17'd57564,17'd51074,17'd56973,17'd33794,17'd30127,17'd23565,17'd29689,17'd23385,17'd23923,17'd32008,17'd22501,17'd22503,17'd31500,17'd31500,17'd31500,17'd31500,17'd45492,17'd31500,17'd30428,17'd32015,17'd32191,17'd29528,17'd34106,17'd29533,17'd28851,17'd30733,17'd53405,17'd60361,17'd50563,17'd57839,17'd62655,17'd34459,17'd38667,17'd33483,17'd39443,17'd33318,17'd32668,17'd38808,17'd48987,17'd50156,17'd57070,17'd57070,17'd63613,17'd53193,17'd42438,17'd43836,17'd43978,17'd32995,17'd63614,17'd63615,17'd63616,17'd63617,17'd36706,17'd32838,17'd26911,17'd27523,17'd62938,17'd63618,17'd63619,17'd63620,17'd63621,17'd63622,17'd63623,17'd63624,17'd63625,17'd25347,17'd19667,17'd63626,17'd23066,17'd63627,17'd63628,17'd63629,17'd62950,17'd63630,17'd63631,17'd63632,17'd63633,17'd19678,17'd20103,17'd21916,17'd22747,17'd43179,17'd22571,17'd63634,17'd23097,17'd23792,17'd9502,17'd10881,17'd23455,17'd24306,17'd54956,17'd54956,17'd22759,17'd26216,17'd24479,17'd7007,17'd5607,17'd5607,17'd5757,17'd4529,17'd4847,17'd40397,17'd63635,17'd38059,17'd5170,17'd51930,17'd37435,17'd35198,17'd6070,17'd63636,17'd63636,17'd62961,17'd63637,17'd63638,17'd15615,17'd15481,17'd63639,17'd63640,17'd25488,17'd63641,17'd13568,17'd18380,17'd18380,17'd63359,17'd12910,17'd63232,17'd62683,17'd30492,17'd30034,17'd29602,17'd31720,17'd61795,17'd7021,17'd62686,17'd19725,17'd19725,17'd63642,17'd62055,17'd62314,17'd3547,17'd63643,17'd63644,17'd37952,17'd63645,17'd63646,17'd63647,17'd56209,17'd56542,17'd63648,17'd63648,17'd23985,17'd63649,17'd56001,17'd54511,17'd63650,17'd52275,17'd37820,17'd2904,17'd235,17'd2739,17'd4424,17'd6885,17'd4423,17'd7211,17'd6889,17'd5630,17'd63651,17'd63651,17'd2393,17'd2393,17'd14586,17'd5777,17'd29169,17'd29610,17'd29170,17'd28793,17'd27822,17'd29040,17'd60625,17'd60625,17'd63652,17'd36905,17'd33051,17'd11336,17'd7365,17'd3896,17'd37709,17'd38203,17'd44019,17'd13056,17'd63653,17'd16381,17'd62848,17'd63372,17'd63373,17'd63654,17'd63655,17'd63655,17'd63656,17'd63378,17'd63511,17'd63657,17'd63658,17'd63512,17'd17913,17'd63659,17'd8786,17'd3379,17'd41475,17'd63660,17'd2217,17'd63661,17'd63662,17'd63663,17'd2072,17'd57757
},
'{
17'd4737,17'd5511,17'd15877,17'd2934,17'd2593,17'd3427,17'd3751,17'd63384,17'd63664,17'd63664,17'd63665,17'd12035,17'd63666,17'd63667,17'd63668,17'd11607,17'd14441,17'd6273,17'd63669,17'd2,17'd4089,17'd3905,17'd17,17'd17187,17'd1414,17'd1414,17'd1127,17'd4247,17'd1831,17'd3101,17'd4892,17'd4087,17'd5203,17'd15359,17'd11609,17'd10547,17'd12194,17'd12194,17'd52621,17'd10924,17'd4086,17'd5204,17'd4891,17'd4425,17'd15496,17'd3751,17'd12196,17'd12653,17'd14989,17'd63670,17'd63671,17'd60278,17'd58379,17'd56440,17'd56009,17'd55892,17'd55892,17'd61413,17'd68,17'd1981,17'd1980,17'd17554,17'd41628,17'd2438,17'd670,17'd488,17'd488,17'd63672,17'd2438,17'd41628,17'd63673,17'd63674,17'd63675,17'd63676,17'd63677,17'd62868,17'd62869,17'd63396,17'd63530,17'd63531,17'd62994,17'd63678,17'd14476,17'd46140,17'd63534,17'd63679,17'd63680,17'd63681,17'd63682,17'd63536,17'd6151,17'd63683,17'd63134,17'd4125,17'd4292,17'd4768,17'd4769,17'd52625,17'd4289,17'd3300,17'd63684,17'd63685,17'd63686,17'd63687,17'd63688,17'd56021,17'd55676,17'd59013,17'd63689,17'd54890,17'd56351,17'd54892,17'd55780,17'd63690,17'd63691,17'd56237,17'd55778,17'd63692,17'd63693,17'd61058,17'd57782,17'd60916,17'd63694,17'd63695,17'd61582,17'd61447,17'd60303,17'd59279,17'd63696,17'd59519,17'd59024,17'd57022,17'd61449,17'd63697,17'd60926,17'd63698,17'd63699,17'd63700,17'd63701,17'd63702,17'd63703,17'd63704,17'd63705,17'd63706,17'd62094,17'd63707,17'd63708,17'd63709,17'd63710,17'd63711,17'd63163,17'd63165,17'd62375,17'd63712,17'd63713,17'd63714,17'd63715,17'd63716,17'd63717,17'd63718,17'd63719,17'd63720,17'd63721,17'd63722,17'd63723,17'd63724,17'd63725,17'd63726,17'd63436,17'd63307,17'd63307,17'd63437,17'd61610,17'd61742,17'd59828,17'd61479,17'd63727,17'd63728,17'd13243,17'd63729,17'd63730,17'd45547,17'd13763,17'd11963,17'd10990,17'd13886,17'd11274,17'd11275,17'd10989,17'd14673,17'd19280,17'd14383,17'd63731,17'd53252,17'd63732,17'd63733,17'd63583,17'd55949,17'd14679,17'd19536,17'd24869,17'd20318,17'd54465,17'd54382,17'd13767,17'd12590,17'd7457,17'd9891,17'd24553,17'd63734,17'd17853,17'd7627,17'd54650,17'd63735,17'd11536,17'd63736,17'd63737,17'd14395,17'd63738,17'd63588,17'd17853,17'd8586,17'd10997,17'd63739,17'd63740,17'd61234,17'd14816,17'd7460,17'd53981,17'd63741,17'd63742,17'd63743,17'd11287,17'd63744,17'd14541,17'd63745,17'd63323,17'd63746,17'd63747,17'd63748,17'd63749,17'd63750,17'd63751,17'd63752,17'd60716,17'd59199,17'd63753,17'd63754,17'd51233,17'd56746,17'd58953,17'd50562,17'd57200,17'd53986,17'd58587,17'd63606,17'd63755,17'd63756,17'd63757,17'd63758,17'd63759,17'd63760,17'd63761,17'd50813,17'd59721,17'd59205,17'd58951,17'd51232,17'd33794,17'd29241,17'd24087,17'd24087,17'd29241,17'd23734,17'd30579,17'd23217,17'd50989,17'd34277,17'd34277,17'd37533,17'd45154,17'd43843,17'd32513,17'd43986,17'd51160,17'd60361,17'd50364,17'd29688,17'd34883,17'd62655,17'd57205,17'd57839,17'd57839,17'd50363,17'd50364,17'd48987,17'd53720,17'd38406,17'd33318,17'd32668,17'd34276,17'd34106,17'd53642,17'd63762,17'd57706,17'd57070,17'd53331,17'd54394,17'd53643,17'd43694,17'd47438,17'd42147,17'd63763,17'd63764,17'd63765,17'd30134,17'd36862,17'd32838,17'd26911,17'd63766,17'd26793,17'd25048,17'd63767,17'd63768,17'd63769,17'd63770,17'd63771,17'd20201,17'd63772,17'd63773,17'd27908,17'd63774,17'd62813,17'd63775,17'd63776,17'd63777,17'd63778,17'd23950,17'd63779,17'd63780,17'd18838,17'd63781,17'd63353,17'd63782,17'd63783,17'd23099,17'd63784,17'd22220,17'd23621,17'd22932,17'd61268,17'd23278,17'd60137,17'd24643,17'd26583,17'd30636,17'd26216,17'd26216,17'd9906,17'd6545,17'd5608,17'd4839,17'd39166,17'd34656,17'd4847,17'd37433,17'd38567,17'd5010,17'd51930,17'd34336,17'd52833,17'd37436,17'd63636,17'd63492,17'd63492,17'd63785,17'd11857,17'd16620,17'd63786,17'd63787,17'd63788,17'd63789,17'd63790,17'd17541,17'd63359,17'd18380,17'd18138,17'd18380,17'd63791,17'd63232,17'd12910,17'd13053,17'd12314,17'd29885,17'd63792,17'd63793,17'd32554,17'd63794,17'd63642,17'd63642,17'd62314,17'd63795,17'd49404,17'd63643,17'd63796,17'd20859,17'd63797,17'd63798,17'd63799,17'd57743,17'd53798,17'd63800,17'd63801,17'd63802,17'd63803,17'd63804,17'd63805,17'd54238,17'd37041,17'd40714,17'd57749,17'd63806,17'd795,17'd2777,17'd1810,17'd4728,17'd4423,17'd16003,17'd4559,17'd5630,17'd63651,17'd16382,17'd12496,17'd16382,17'd14586,17'd33050,17'd27707,17'd29892,17'd29170,17'd29170,17'd27822,17'd29040,17'd60625,17'd60625,17'd63652,17'd36903,17'd33051,17'd8507,17'd4730,17'd37709,17'd38203,17'd38580,17'd44019,17'd62445,17'd14735,17'd63371,17'd63372,17'd63106,17'd63807,17'd63655,17'd63655,17'd63244,17'd63808,17'd63378,17'd63657,17'd63809,17'd63658,17'd63512,17'd63810,17'd63659,17'd63811,17'd41903,17'd41768,17'd33694,17'd53003,17'd26590,17'd63812,17'd63663,17'd56002,17'd58253
},
'{
17'd4893,17'd5204,17'd15877,17'd15358,17'd2934,17'd3427,17'd3751,17'd63813,17'd63814,17'd63815,17'd63816,17'd63817,17'd63818,17'd63819,17'd63820,17'd63821,17'd63821,17'd63822,17'd6101,17'd3749,17'd8971,17'd12,17'd2595,17'd1830,17'd1967,17'd1127,17'd1127,17'd1127,17'd1689,17'd2422,17'd3427,17'd15496,17'd5203,17'd5511,17'd15496,17'd3427,17'd3101,17'd3252,17'd2935,17'd2934,17'd3592,17'd5204,17'd5511,17'd52704,17'd5511,17'd3592,17'd3751,17'd63254,17'd14320,17'd14322,17'd63388,17'd63823,17'd63824,17'd63825,17'd56332,17'd56010,17'd19500,17'd1981,17'd1981,17'd485,17'd1980,17'd17554,17'd2789,17'd62,17'd669,17'd2615,17'd488,17'd672,17'd62341,17'd62211,17'd54787,17'd61950,17'd63826,17'd63827,17'd63828,17'd63125,17'd63829,17'd63830,17'd63831,17'd63832,17'd63833,17'd63834,17'd63835,17'd63836,17'd63837,17'd63838,17'd63839,17'd63840,17'd63136,17'd6774,17'd6151,17'd6775,17'd63134,17'd60290,17'd4291,17'd63841,17'd63842,17'd59513,17'd4288,17'd3138,17'd63843,17'd59642,17'd3634,17'd58395,17'd63844,17'd63845,17'd54892,17'd56582,17'd63846,17'd63846,17'd63141,17'd56351,17'd55380,17'd57510,17'd57639,17'd56579,17'd57783,17'd63847,17'd63847,17'd58886,17'd58772,17'd58041,17'd56913,17'd58651,17'd61449,17'd59647,17'd60658,17'd58527,17'd63848,17'd60428,17'd57922,17'd59281,17'd62475,17'd61313,17'd59649,17'd63849,17'd63850,17'd63851,17'd63852,17'd63701,17'd63853,17'd63854,17'd63855,17'd63856,17'd54099,17'd53451,17'd63857,17'd63858,17'd63859,17'd63424,17'd63860,17'd63861,17'd62376,17'd63862,17'd63716,17'd63863,17'd63863,17'd63864,17'd63865,17'd63866,17'd63867,17'd63569,17'd62757,17'd63868,17'd63869,17'd63172,17'd63435,17'd63726,17'd63870,17'd63870,17'd63871,17'd63872,17'd63035,17'd63873,17'd60215,17'd63874,17'd63875,17'd63876,17'd62140,17'd22809,17'd63877,17'd63878,17'd45093,17'd13365,17'd20910,17'd10991,17'd11670,17'd11670,17'd13886,17'd10605,17'd15176,17'd11671,17'd50112,17'd29919,17'd8105,17'd14680,17'd15303,17'd25681,17'd12428,17'd15949,17'd53109,17'd21058,17'd16078,17'd15436,17'd14531,17'd7620,17'd63879,17'd11969,17'd12267,17'd18087,17'd14142,17'd12268,17'd18454,17'd11816,17'd9489,17'd7634,17'd63880,17'd18924,17'd63185,17'd63881,17'd63739,17'd63882,17'd54045,17'd21509,17'd63883,17'd53191,17'd10482,17'd8428,17'd63884,17'd63885,17'd24875,17'd17859,17'd63886,17'd16087,17'd23014,17'd63744,17'd63887,17'd43115,17'd63888,17'd63889,17'd63890,17'd63891,17'd63892,17'd63893,17'd63894,17'd63895,17'd63896,17'd57970,17'd63897,17'd52162,17'd50461,17'd49171,17'd56968,17'd50820,17'd53986,17'd51554,17'd63898,17'd63899,17'd63900,17'd63901,17'd63902,17'd63903,17'd63904,17'd63905,17'd63906,17'd50813,17'd51914,17'd58707,17'd56507,17'd30578,17'd29375,17'd32186,17'd29528,17'd30127,17'd29827,17'd48257,17'd29531,17'd29374,17'd23387,17'd35865,17'd24421,17'd23388,17'd30128,17'd31190,17'd56507,17'd63907,17'd60361,17'd57839,17'd63907,17'd50563,17'd57205,17'd57839,17'd62655,17'd50364,17'd34459,17'd33793,17'd33802,17'd33793,17'd40964,17'd34106,17'd63908,17'd63909,17'd63910,17'd63911,17'd63911,17'd57707,17'd55722,17'd63912,17'd63913,17'd43550,17'd63914,17'd29824,17'd33477,17'd37135,17'd29541,17'd63915,17'd30888,17'd26909,17'd30747,17'd27270,17'd28871,17'd63916,17'd63917,17'd63918,17'd63919,17'd63920,17'd63921,17'd63922,17'd63923,17'd63924,17'd63925,17'd63926,17'd63927,17'd63928,17'd63929,17'd63930,17'd21100,17'd63931,17'd63932,17'd63933,17'd63934,17'd19581,17'd63935,17'd63936,17'd63783,17'd22069,17'd21903,17'd22741,17'd63937,17'd24304,17'd30793,17'd24306,17'd24643,17'd26111,17'd61528,17'd22759,17'd6544,17'd7324,17'd24798,17'd5607,17'd4840,17'd32552,17'd32552,17'd4841,17'd4684,17'd37153,17'd5007,17'd5011,17'd37435,17'd8474,17'd37698,17'd63490,17'd5484,17'd6071,17'd62825,17'd12166,17'd13804,17'd63938,17'd63939,17'd63940,17'd63941,17'd63942,17'd63943,17'd63944,17'd63945,17'd63946,17'd63946,17'd18030,17'd17910,17'd17910,17'd13568,17'd19229,17'd18750,17'd12631,17'd63947,17'd19231,17'd63948,17'd4214,17'd61272,17'd33045,17'd49501,17'd63949,17'd33535,17'd63950,17'd46133,17'd63951,17'd63952,17'd63953,17'd63954,17'd63955,17'd63956,17'd62192,17'd63957,17'd23985,17'd63649,17'd25778,17'd62705,17'd63958,17'd52458,17'd3067,17'd57891,17'd54777,17'd1402,17'd2096,17'd4422,17'd4423,17'd6415,17'd5940,17'd5940,17'd5630,17'd8185,17'd8185,17'd5776,17'd4714,17'd2906,17'd33050,17'd27707,17'd27708,17'd28793,17'd28792,17'd28793,17'd28793,17'd29611,17'd29611,17'd36904,17'd58864,17'd7537,17'd6095,17'd5028,17'd37957,17'd38580,17'd44019,17'd63959,17'd63960,17'd63961,17'd62969,17'd63106,17'd63962,17'd63963,17'd63963,17'd63655,17'd63244,17'd63964,17'd63965,17'd63657,17'd63809,17'd63966,17'd63967,17'd63968,17'd12174,17'd62072,17'd49902,17'd41902,17'd63969,17'd63970,17'd63971,17'd2214,17'd63972,17'd56002,17'd58135
},
'{
17'd6730,17'd6730,17'd52704,17'd15496,17'd3901,17'd3901,17'd3901,17'd63384,17'd63814,17'd63973,17'd63974,17'd63975,17'd63976,17'd63977,17'd63978,17'd63979,17'd13433,17'd63980,17'd6267,17'd63118,17'd2595,17'd0,17'd1127,17'd1830,17'd1967,17'd1689,17'd1127,17'd1127,17'd1689,17'd2422,17'd3251,17'd15496,17'd5511,17'd5511,17'd15496,17'd3901,17'd2934,17'd2935,17'd2935,17'd2934,17'd3592,17'd15496,17'd5511,17'd52704,17'd5511,17'd5204,17'd3901,17'd2783,17'd12504,17'd15629,17'd63261,17'd63981,17'd63982,17'd63983,17'd57109,17'd56116,17'd21473,17'd14451,17'd486,17'd486,17'd1980,17'd17791,17'd2789,17'd2789,17'd1843,17'd1148,17'd488,17'd489,17'd63984,17'd63985,17'd54787,17'd32886,17'd61039,17'd63986,17'd63987,17'd63988,17'd63989,17'd63990,17'd63831,17'd63832,17'd63839,17'd8847,17'd63991,17'd63992,17'd63993,17'd63838,17'd63994,17'd63401,17'd63995,17'd61301,17'd6151,17'd63537,17'd63136,17'd5083,17'd44521,17'd59011,17'd63996,17'd63997,17'd4288,17'd63138,17'd3136,17'd4466,17'd63998,17'd63999,17'd58027,17'd53880,17'd64000,17'd55584,17'd61967,17'd61576,17'd54801,17'd56351,17'd55675,17'd55380,17'd55676,17'd55282,17'd64001,17'd64002,17'd64003,17'd64003,17'd57921,17'd58653,17'd56913,17'd64004,17'd58893,17'd59019,17'd58894,17'd60922,17'd64005,17'd59145,17'd60428,17'd58893,17'd58768,17'd58768,17'd56697,17'd61707,17'd64006,17'd64007,17'd64008,17'd64009,17'd64010,17'd64011,17'd64012,17'd64013,17'd64014,17'd43887,17'd64015,17'd64016,17'd64017,17'd64018,17'd64019,17'd64020,17'd62376,17'd63862,17'd64021,17'd64022,17'd64023,17'd64024,17'd64025,17'd63866,17'd63718,17'd63719,17'd62901,17'd61870,17'd61214,17'd63723,17'd63724,17'd63726,17'd64026,17'd64027,17'd63871,17'd64028,17'd63035,17'd63873,17'd60958,17'd63176,17'd64029,17'd64030,17'd64031,17'd17959,17'd64032,17'd54278,17'd17015,17'd12575,17'd18560,17'd19282,17'd10479,17'd11528,17'd12863,17'd13886,17'd14134,17'd10330,17'd26034,17'd26626,17'd16916,17'd12726,17'd21508,17'd15946,17'd16447,17'd16447,17'd21508,17'd64033,17'd14390,17'd16078,17'd13893,17'd14011,17'd9052,17'd13770,17'd13529,17'd15444,17'd17732,17'd12730,17'd62390,17'd12269,17'd15698,17'd64034,17'd64035,17'd18924,17'd54735,17'd20457,17'd21825,17'd21825,17'd10863,17'd7627,17'd17356,17'd16695,17'd24873,17'd7627,17'd64036,17'd64037,17'd64038,17'd11976,17'd24561,17'd19542,17'd22145,17'd64039,17'd64040,17'd64041,17'd64042,17'd64043,17'd64044,17'd64045,17'd64046,17'd64047,17'd64048,17'd64049,17'd64050,17'd63605,17'd63897,17'd57325,17'd56746,17'd64051,17'd63466,17'd50992,17'd53986,17'd51554,17'd61769,17'd50645,17'd64052,17'd64053,17'd63901,17'd64054,17'd63903,17'd63904,17'd64055,17'd63761,17'd64056,17'd64057,17'd58824,17'd58091,17'd33652,17'd30424,17'd29527,17'd29241,17'd23733,17'd23918,17'd23918,17'd23733,17'd23920,17'd29241,17'd23734,17'd31502,17'd23734,17'd56973,17'd56285,17'd50563,17'd63907,17'd63907,17'd50730,17'd50563,17'd57839,17'd62655,17'd38978,17'd48987,17'd33793,17'd33802,17'd33793,17'd34282,17'd33644,17'd50363,17'd64058,17'd64058,17'd64059,17'd64060,17'd64061,17'd61902,17'd64062,17'd64063,17'd64064,17'd44359,17'd64065,17'd29824,17'd33154,17'd42444,17'd29541,17'd64066,17'd29543,17'd29698,17'd30290,17'd30891,17'd24910,17'd64067,17'd64068,17'd64069,17'd64070,17'd25060,17'd64071,17'd25061,17'd64072,17'd64073,17'd64074,17'd22536,17'd64075,17'd64075,17'd64076,17'd23419,17'd64077,17'd22363,17'd64078,17'd64079,17'd64080,17'd64081,17'd64082,17'd22577,17'd64083,17'd64084,17'd22064,17'd64085,17'd23791,17'd24304,17'd24642,17'd64086,17'd25767,17'd26111,17'd22759,17'd11158,17'd6544,17'd7324,17'd24649,17'd4993,17'd32552,17'd4687,17'd4687,17'd4686,17'd37153,17'd29024,17'd4849,17'd5013,17'd52833,17'd52762,17'd35479,17'd6396,17'd5341,17'd7185,17'd10900,17'd17069,17'd14055,17'd64087,17'd64088,17'd64089,17'd64090,17'd63942,17'd63943,17'd64091,17'd63945,17'd63946,17'd63945,17'd18030,17'd17783,17'd17910,17'd63231,17'd14057,17'd18506,17'd64092,17'd62311,17'd64093,17'd19231,17'd63948,17'd63234,17'd64094,17'd64095,17'd64096,17'd64097,17'd64098,17'd21621,17'd64099,17'd64100,17'd64101,17'd64102,17'd64103,17'd61398,17'd53359,17'd63957,17'd23985,17'd63803,17'd23640,17'd64104,17'd61032,17'd40714,17'd19360,17'd58372,17'd5627,17'd5629,17'd2240,17'd4728,17'd4423,17'd5940,17'd5940,17'd5940,17'd8185,17'd35907,17'd35907,17'd8186,17'd6416,17'd11061,17'd27949,17'd27708,17'd29170,17'd28793,17'd28792,17'd28793,17'd29170,17'd29611,17'd36904,17'd64105,17'd58865,17'd6418,17'd38459,17'd5028,17'd38334,17'd38580,17'd62329,17'd64106,17'd64107,17'd64108,17'd63105,17'd63106,17'd63962,17'd63963,17'd63963,17'd63108,17'd63244,17'd64109,17'd64110,17'd64111,17'd63809,17'd64112,17'd63967,17'd63968,17'd18269,17'd62205,17'd49902,17'd41902,17'd63969,17'd33995,17'd64113,17'd2214,17'd64114,17'd59488,17'd64115
},
'{
17'd64116,17'd5203,17'd52704,17'd15877,17'd3592,17'd3592,17'd3901,17'd64117,17'd63664,17'd64118,17'd63975,17'd64119,17'd64120,17'd64121,17'd64122,17'd13815,17'd64123,17'd64124,17'd9683,17'd64125,17'd1127,17'd2,17'd1127,17'd15,17'd1415,17'd1414,17'd1416,17'd1416,17'd1414,17'd2597,17'd14070,17'd3428,17'd15496,17'd5511,17'd15496,17'd3428,17'd3101,17'd2935,17'd2935,17'd3101,17'd3427,17'd3592,17'd5511,17'd52704,17'd5511,17'd5204,17'd3901,17'd3751,17'd12505,17'd58016,17'd15243,17'd64126,17'd64127,17'd63824,17'd56789,17'd56011,17'd21473,17'd14451,17'd486,17'd486,17'd18151,17'd17791,17'd2789,17'd2789,17'd1709,17'd1843,17'd488,17'd489,17'd62210,17'd62341,17'd54787,17'd54693,17'd61684,17'd61555,17'd64128,17'd64129,17'd64130,17'd64131,17'd64132,17'd63272,17'd64133,17'd63839,17'd64134,17'd64134,17'd64135,17'd64136,17'd63994,17'd63401,17'd64137,17'd64138,17'd64139,17'd6308,17'd6316,17'd64140,17'd5083,17'd4768,17'd8688,17'd59011,17'd4462,17'd3945,17'd53303,17'd4771,17'd64141,17'd59142,17'd58027,17'd64142,17'd63001,17'd54704,17'd64143,17'd54801,17'd63277,17'd64144,17'd55675,17'd55184,17'd55902,17'd64145,17'd54890,17'd63405,17'd64146,17'd64147,17'd56237,17'd61059,17'd58653,17'd57396,17'd57279,17'd64148,17'd58769,17'd59647,17'd64149,17'd60541,17'd60663,17'd64150,17'd59024,17'd57022,17'd58660,17'd57397,17'd64151,17'd64152,17'd3023,17'd64153,17'd64154,17'd64155,17'd64156,17'd5423,17'd5855,17'd64157,17'd6635,17'd64158,17'd64159,17'd32113,17'd64160,17'd64161,17'd64162,17'd64163,17'd63712,17'd64024,17'd64164,17'd64164,17'd64165,17'd64166,17'd64167,17'd64168,17'd64169,17'd63721,17'd61468,17'd62904,17'd63724,17'd63726,17'd64026,17'd64026,17'd64170,17'd64028,17'd63035,17'd63438,17'd61742,17'd60087,17'd64171,17'd64172,17'd64173,17'd13995,17'd64174,17'd53706,17'd45209,17'd13513,17'd16797,17'd16555,17'd10741,17'd10479,17'd11134,17'd11527,17'd12721,17'd11670,17'd11134,17'd18080,17'd8579,17'd12589,17'd25929,17'd15060,17'd16802,17'd15440,17'd10180,17'd19036,17'd19536,17'd18921,17'd21059,17'd13769,17'd24552,17'd12868,17'd15444,17'd13772,17'd18811,17'd64175,17'd62772,17'd23875,17'd15577,17'd23874,17'd8116,17'd25537,17'd22827,17'd64176,17'd60101,17'd10863,17'd7628,17'd7628,17'd14939,17'd64177,17'd14818,17'd17854,17'd10033,17'd8121,17'd9754,17'd11007,17'd23883,17'd64178,17'd9755,17'd19043,17'd14274,17'd64179,17'd64180,17'd64181,17'd64182,17'd64183,17'd64184,17'd64185,17'd64186,17'd64187,17'd64188,17'd64189,17'd64190,17'd50734,17'd52162,17'd56967,17'd57071,17'd64191,17'd64192,17'd58711,17'd58826,17'd64193,17'd59581,17'd64194,17'd64195,17'd64196,17'd64197,17'd64198,17'd64199,17'd64200,17'd64201,17'd60360,17'd58707,17'd60480,17'd58091,17'd53556,17'd55228,17'd55228,17'd55228,17'd56973,17'd56973,17'd56973,17'd55228,17'd35430,17'd33950,17'd35430,17'd58091,17'd56285,17'd56285,17'd50563,17'd63907,17'd50563,17'd56285,17'd56285,17'd57205,17'd50363,17'd33644,17'd34459,17'd33802,17'd54061,17'd48987,17'd48987,17'd50364,17'd50363,17'd64058,17'd64202,17'd64203,17'd64204,17'd64205,17'd64206,17'd52584,17'd64207,17'd64208,17'd45036,17'd64209,17'd29824,17'd33478,17'd64210,17'd29541,17'd34130,17'd30900,17'd36560,17'd28272,17'd64211,17'd64212,17'd64213,17'd64214,17'd25595,17'd64215,17'd64216,17'd64071,17'd25061,17'd63477,17'd64217,17'd19947,17'd64218,17'd64219,17'd64220,17'd20344,17'd23419,17'd64221,17'd64222,17'd64223,17'd64224,17'd20805,17'd26932,17'd26442,17'd22749,17'd22743,17'd23098,17'd22742,17'd57727,17'd23791,17'd24304,17'd24642,17'd64086,17'd25878,17'd54956,17'd11158,17'd11158,17'd6544,17'd7324,17'd24649,17'd4994,17'd4688,17'd4687,17'd4687,17'd4842,17'd29024,17'd4848,17'd5011,17'd53353,17'd52833,17'd34923,17'd5483,17'd6396,17'd34795,17'd34659,17'd12007,17'd16852,17'd15731,17'd64225,17'd64226,17'd64227,17'd63640,17'd63788,17'd64091,17'd63945,17'd63946,17'd63946,17'd63945,17'd18030,17'd18030,17'd18030,17'd14057,17'd17177,17'd18379,17'd18505,17'd62426,17'd64228,17'd62053,17'd62685,17'd61394,17'd64229,17'd49602,17'd64230,17'd64231,17'd64232,17'd64233,17'd64234,17'd43191,17'd42330,17'd35612,17'd64235,17'd64236,17'd64237,17'd64238,17'd63803,17'd27944,17'd54871,17'd64104,17'd61162,17'd64239,17'd58373,17'd54975,17'd64240,17'd11589,17'd2096,17'd4423,17'd4423,17'd4423,17'd4728,17'd4423,17'd3391,17'd3391,17'd4729,17'd9123,17'd4714,17'd5030,17'd36602,17'd29892,17'd28792,17'd27822,17'd27822,17'd28793,17'd29170,17'd29611,17'd58990,17'd58864,17'd7878,17'd6258,17'd39328,17'd37957,17'd38334,17'd38580,17'd44019,17'd43596,17'd15735,17'd62847,17'd63105,17'd63807,17'd63807,17'd63963,17'd63963,17'd63108,17'd63244,17'd64109,17'd63965,17'd63809,17'd64241,17'd64242,17'd64243,17'd64244,17'd18269,17'd64245,17'd49902,17'd46475,17'd64246,17'd33843,17'd64247,17'd64248,17'd64249,17'd24492,17'd64250
},
'{
17'd64116,17'd15117,17'd15359,17'd52704,17'd5204,17'd5204,17'd4086,17'd64251,17'd64252,17'd63973,17'd63975,17'd63975,17'd64120,17'd64253,17'd64121,17'd64254,17'd64255,17'd64256,17'd9270,17'd10923,17'd1967,17'd14,17'd14,17'd14,17'd1415,17'd1414,17'd1416,17'd1416,17'd1414,17'd2597,17'd3252,17'd3427,17'd15496,17'd5204,17'd15496,17'd3428,17'd3251,17'd2935,17'd2935,17'd2934,17'd3901,17'd3592,17'd5204,17'd5511,17'd5511,17'd5204,17'd3592,17'd3901,17'd12196,17'd16392,17'd15361,17'd64257,17'd64258,17'd64259,17'd64260,17'd64261,17'd15248,17'd14872,17'd1981,17'd486,17'd485,17'd18391,17'd17554,17'd995,17'd17554,17'd1843,17'd62340,17'd489,17'd60894,17'd18391,17'd54787,17'd54693,17'd64262,17'd64263,17'd64264,17'd64265,17'd64266,17'd64267,17'd64268,17'd64269,17'd64270,17'd63992,17'd64271,17'd64272,17'd64273,17'd64274,17'd9985,17'd64275,17'd60903,17'd62223,17'd64139,17'd64276,17'd6006,17'd64277,17'd63134,17'd4126,17'd7088,17'd4766,17'd5082,17'd4461,17'd3623,17'd3477,17'd53954,17'd53448,17'd58027,17'd64278,17'd64279,17'd64280,17'd60299,17'd64281,17'd57389,17'd64282,17'd55280,17'd64283,17'd60170,17'd60422,17'd56580,17'd54890,17'd57782,17'd64284,17'd64285,17'd64286,17'd58653,17'd57132,17'd58892,17'd62473,17'd60427,17'd59150,17'd64287,17'd58038,17'd64288,17'd64289,17'd58654,17'd56244,17'd54898,17'd61579,17'd63008,17'd64290,17'd64291,17'd64292,17'd64293,17'd64294,17'd4792,17'd64295,17'd64296,17'd53689,17'd6473,17'd8378,17'd15536,17'd18422,17'd34024,17'd64297,17'd64298,17'd64163,17'd64299,17'd63865,17'd64165,17'd64165,17'd64300,17'd64166,17'd64167,17'd64301,17'd64302,17'd62503,17'd64303,17'd64304,17'd63034,17'd63572,17'd64305,17'd64026,17'd64170,17'd64028,17'd63173,17'd63438,17'd61742,17'd64306,17'd64307,17'd64308,17'd58071,17'd14250,17'd57312,17'd13510,17'd61482,17'd13361,17'd15564,17'd10853,17'd10328,17'd16796,17'd17719,17'd10479,17'd10478,17'd12863,17'd9883,17'd49324,17'd24711,17'd8734,17'd25152,17'd10995,17'd14385,17'd7789,17'd7619,17'd22135,17'd18921,17'd21059,17'd12429,17'd14266,17'd10343,17'd18922,17'd15696,17'd18924,17'd18571,17'd59706,17'd61748,17'd55708,17'd23875,17'd8431,17'd23526,17'd18691,17'd64309,17'd22827,17'd19038,17'd7628,17'd64310,17'd54650,17'd64311,17'd15063,17'd55125,17'd64312,17'd8591,17'd64313,17'd7976,17'd15069,17'd64314,17'd64314,17'd13533,17'd22839,17'd64315,17'd64316,17'd64317,17'd64318,17'd64319,17'd64320,17'd64321,17'd62274,17'd64322,17'd64323,17'd64324,17'd64325,17'd59084,17'd64326,17'd52162,17'd56967,17'd57200,17'd64327,17'd64328,17'd64192,17'd61500,17'd57841,17'd50728,17'd59860,17'd64329,17'd64330,17'd64331,17'd64332,17'd64199,17'd64333,17'd64334,17'd64335,17'd64336,17'd51473,17'd60480,17'd56507,17'd55228,17'd55228,17'd56973,17'd63907,17'd63907,17'd63907,17'd56973,17'd55228,17'd56973,17'd63907,17'd56285,17'd56285,17'd63907,17'd63907,17'd50563,17'd56285,17'd57967,17'd57205,17'd50363,17'd33644,17'd34459,17'd34282,17'd33802,17'd34113,17'd34621,17'd38978,17'd62655,17'd57205,17'd64202,17'd64059,17'd64337,17'd64061,17'd64205,17'd64338,17'd64339,17'd64063,17'd64208,17'd64340,17'd46095,17'd45749,17'd64341,17'd64342,17'd64343,17'd38030,17'd36862,17'd30136,17'd64344,17'd37672,17'd64345,17'd64346,17'd23754,17'd64347,17'd64348,17'd64349,17'd64071,17'd64350,17'd64351,17'd64352,17'd64353,17'd64354,17'd64355,17'd64356,17'd64218,17'd64218,17'd64357,17'd64358,17'd64359,17'd64360,17'd20963,17'd64361,17'd64362,17'd64363,17'd64364,17'd22220,17'd22921,17'd23622,17'd24142,17'd24305,17'd24943,17'd64365,17'd26111,17'd26215,17'd22587,17'd10196,17'd6702,17'd24650,17'd5324,17'd5326,17'd4687,17'd5005,17'd5005,17'd4842,17'd4848,17'd5007,17'd5013,17'd5617,17'd52762,17'd34923,17'd5483,17'd9784,17'd34795,17'd11580,17'd17069,17'd14973,17'd64366,17'd64367,17'd64368,17'd64369,17'd63640,17'd64370,17'd14432,17'd63946,17'd63946,17'd63946,17'd63945,17'd63945,17'd18030,17'd63945,17'd17177,17'd16622,17'd18379,17'd27431,17'd64092,17'd62312,17'd64228,17'd63233,17'd31246,17'd64371,17'd64372,17'd49301,17'd64373,17'd64374,17'd64375,17'd64376,17'd64377,17'd64378,17'd64379,17'd64380,17'd64381,17'd24160,17'd63649,17'd25778,17'd64382,17'd64383,17'd54873,17'd64384,17'd21322,17'd18981,17'd7025,17'd64385,17'd11589,17'd50843,17'd3423,17'd3391,17'd4085,17'd4423,17'd4423,17'd4085,17'd4085,17'd4713,17'd4714,17'd4714,17'd5030,17'd35207,17'd28793,17'd27711,17'd31410,17'd27822,17'd28793,17'd31251,17'd36903,17'd58864,17'd58865,17'd6418,17'd37959,17'd38203,17'd38202,17'd38334,17'd38580,17'd62329,17'd63960,17'd63961,17'd63241,17'd64386,17'd63807,17'd64387,17'd63963,17'd63655,17'd63244,17'd63808,17'd64109,17'd64110,17'd64388,17'd63809,17'd64112,17'd64389,17'd64390,17'd18269,17'd64245,17'd49902,17'd46475,17'd2529,17'd33995,17'd64247,17'd64391,17'd64114,17'd59488,17'd24320
},
'{
17'd64392,17'd64116,17'd15359,17'd52704,17'd5511,17'd5511,17'd5204,17'd4737,17'd64393,17'd64394,17'd64395,17'd64395,17'd64396,17'd63976,17'd63977,17'd64397,17'd64398,17'd64255,17'd64399,17'd9967,17'd64400,17'd14,17'd1415,17'd1415,17'd17,17'd1416,17'd4089,17'd3905,17'd17,17'd1414,17'd2258,17'd10802,17'd3592,17'd5204,17'd15496,17'd15358,17'd3251,17'd3101,17'd3101,17'd3101,17'd3427,17'd3592,17'd5204,17'd5511,17'd5511,17'd5204,17'd4086,17'd3901,17'd12505,17'd36,17'd14989,17'd63670,17'd64401,17'd59912,17'd299,17'd57001,17'd55660,17'd15248,17'd62710,17'd1981,17'd670,17'd63672,17'd55276,17'd995,17'd2438,17'd17554,17'd671,17'd489,17'd670,17'd669,17'd1709,17'd63265,17'd64402,17'd64403,17'd64404,17'd64405,17'd64406,17'd64407,17'd64408,17'd64409,17'd64410,17'd64411,17'd64412,17'd64413,17'd64414,17'd8220,17'd9842,17'd63994,17'd5687,17'd64415,17'd62092,17'd6007,17'd62093,17'd64416,17'd6477,17'd5084,17'd6306,17'd4464,17'd4125,17'd4609,17'd64417,17'd63686,17'd53448,17'd53448,17'd57910,17'd53522,17'd53758,17'd64418,17'd59930,17'd56688,17'd56689,17'd57637,17'd56449,17'd64419,17'd57506,17'd60170,17'd59516,17'd64420,17'd64421,17'd64422,17'd64423,17'd64423,17'd58041,17'd57021,17'd57021,17'd58406,17'd57275,17'd58893,17'd55905,17'd58038,17'd63407,17'd63848,17'd64148,17'd64424,17'd58660,17'd59524,17'd61313,17'd64425,17'd64426,17'd64427,17'd64428,17'd64429,17'd64430,17'd64431,17'd64432,17'd64433,17'd6631,17'd7100,17'd12822,17'd10124,17'd15149,17'd64434,17'd64435,17'd64436,17'd64437,17'd64025,17'd64300,17'd64300,17'd64438,17'd64439,17'd64167,17'd64167,17'd64440,17'd64441,17'd64442,17'd62505,17'd63571,17'd63572,17'd64305,17'd64026,17'd64170,17'd63871,17'd64443,17'd62258,17'd63438,17'd62764,17'd64444,17'd59831,17'd64445,17'd64446,17'd23845,17'd62910,17'd61615,17'd13884,17'd64447,17'd16797,17'd27864,17'd24542,17'd9885,17'd11277,17'd10479,17'd20756,17'd10169,17'd17473,17'd64448,17'd11674,17'd8254,17'd7787,17'd9485,17'd63445,17'd63446,17'd7620,17'd7458,17'd7791,17'd24369,17'd24550,17'd10863,17'd19161,17'd61230,17'd62914,17'd62390,17'd55708,17'd61748,17'd61748,17'd21372,17'd25007,17'd61233,17'd64449,17'd64450,17'd64451,17'd23871,17'd7630,17'd64452,17'd7631,17'd15196,17'd13895,17'd59841,17'd12871,17'd64453,17'd9357,17'd64454,17'd9495,17'd64178,17'd64455,17'd9755,17'd23014,17'd16577,17'd64456,17'd64457,17'd64458,17'd64459,17'd64460,17'd64461,17'd64462,17'd64463,17'd64464,17'd64465,17'd59714,17'd64466,17'd58208,17'd50646,17'd56967,17'd57326,17'd50646,17'd57708,17'd61500,17'd64467,17'd63897,17'd58208,17'd64468,17'd60113,17'd63337,17'd64330,17'd64188,17'd64469,17'd64470,17'd64471,17'd64471,17'd64472,17'd60360,17'd64473,17'd60480,17'd59453,17'd59453,17'd51232,17'd56507,17'd58334,17'd50730,17'd50563,17'd50563,17'd50563,17'd56285,17'd56285,17'd50563,17'd60361,17'd57839,17'd62797,17'd62797,17'd62797,17'd62797,17'd57076,17'd50156,17'd34282,17'd34282,17'd34459,17'd48987,17'd38978,17'd62655,17'd57839,17'd56285,17'd64202,17'd64203,17'd64474,17'd64475,17'd64206,17'd64476,17'd64477,17'd64207,17'd53051,17'd64478,17'd46095,17'd46095,17'd64479,17'd64480,17'd64481,17'd62937,17'd29985,17'd30758,17'd28733,17'd24102,17'd64482,17'd24268,17'd64483,17'd64484,17'd27395,17'd64485,17'd64486,17'd64487,17'd64488,17'd64489,17'd64490,17'd64491,17'd64492,17'd64493,17'd64494,17'd64494,17'd64495,17'd64496,17'd64497,17'd28628,17'd19208,17'd64498,17'd64499,17'd64500,17'd64501,17'd22568,17'd57727,17'd63937,17'd22932,17'd30793,17'd24943,17'd25997,17'd54956,17'd26327,17'd11294,17'd8608,17'd6544,17'd24649,17'd4993,17'd5479,17'd5478,17'd4843,17'd5005,17'd30637,17'd5009,17'd5010,17'd5013,17'd53353,17'd52762,17'd8937,17'd64502,17'd10239,17'd64503,17'd12310,17'd13565,17'd15731,17'd64504,17'd64505,17'd64506,17'd64507,17'd63788,17'd64508,17'd18138,17'd18138,17'd14432,17'd14432,17'd63944,17'd63944,17'd63944,17'd14432,17'd64509,17'd15230,17'd14172,17'd18266,17'd13288,17'd12631,17'd11716,17'd19097,17'd64510,17'd4217,17'd4548,17'd64511,17'd64512,17'd64513,17'd64514,17'd64515,17'd64516,17'd64517,17'd64518,17'd64519,17'd24160,17'd64520,17'd64521,17'd35203,17'd63253,17'd2528,17'd64522,17'd37818,17'd52533,17'd64523,17'd5352,17'd64524,17'd17786,17'd5357,17'd3246,17'd3246,17'd3897,17'd4575,17'd3897,17'd3423,17'd4085,17'd4728,17'd6889,17'd5183,17'd33050,17'd29611,17'd28792,17'd31410,17'd31410,17'd27822,17'd60625,17'd29611,17'd58990,17'd58864,17'd64525,17'd6258,17'd4867,17'd37958,17'd38202,17'd38334,17'd44019,17'd63959,17'd62574,17'd63371,17'd64386,17'd64526,17'd64387,17'd64387,17'd63655,17'd63655,17'd63244,17'd64527,17'd63658,17'd64528,17'd63809,17'd64241,17'd64529,17'd64530,17'd64531,17'd64532,17'd64245,17'd41904,17'd46475,17'd64533,17'd64534,17'd52529,17'd64391,17'd2215,17'd59623,17'd24320
},
'{
17'd64392,17'd64116,17'd5203,17'd15359,17'd5511,17'd5511,17'd5203,17'd4893,17'd64535,17'd64536,17'd63974,17'd63974,17'd64396,17'd64396,17'd63977,17'd64537,17'd64538,17'd64538,17'd64399,17'd63668,17'd63260,17'd1967,17'd1415,17'd1415,17'd17,17'd1416,17'd4089,17'd3905,17'd17,17'd1414,17'd2597,17'd3593,17'd3901,17'd3592,17'd15358,17'd15358,17'd34512,17'd3251,17'd3101,17'd2934,17'd3901,17'd3592,17'd5204,17'd5511,17'd5511,17'd5204,17'd4086,17'd13943,17'd10924,17'd294,17'd14320,17'd15361,17'd43,17'd64539,17'd45,17'd299,17'd50,17'd55660,17'd19500,17'd1981,17'd837,17'd63672,17'd63672,17'd669,17'd2438,17'd17554,17'd64540,17'd62340,17'd670,17'd2439,17'd1843,17'd63673,17'd64402,17'd63674,17'd64541,17'd64542,17'd64543,17'd64544,17'd64545,17'd64546,17'd63397,17'd64547,17'd64548,17'd64413,17'd39646,17'd7917,17'd8847,17'd9985,17'd63401,17'd63995,17'd64549,17'd6310,17'd53305,17'd61834,17'd62723,17'd63681,17'd4924,17'd6306,17'd4292,17'd52625,17'd3621,17'd64550,17'd53302,17'd58396,17'd57910,17'd59143,17'd64142,17'd64551,17'd64552,17'd57506,17'd64283,17'd64553,17'd56449,17'd64419,17'd57506,17'd59930,17'd54803,17'd56689,17'd64554,17'd64555,17'd64422,17'd64284,17'd56909,17'd55091,17'd64556,17'd58772,17'd57783,17'd64004,17'd59523,17'd64557,17'd59932,17'd62359,17'd1320,17'd59650,17'd59024,17'd62475,17'd56807,17'd56583,17'd64558,17'd56814,17'd3328,17'd64292,17'd64559,17'd64560,17'd64561,17'd64562,17'd54261,17'd7915,17'd24524,17'd10124,17'd64563,17'd33391,17'd64564,17'd64565,17'd64566,17'd64567,17'd64568,17'd64439,17'd64300,17'd64439,17'd64569,17'd64569,17'd64301,17'd64570,17'd64571,17'd64572,17'd63723,17'd64573,17'd63726,17'd64026,17'd64170,17'd63871,17'd64443,17'd62382,17'd61474,17'd64574,17'd63176,17'd64575,17'd63440,17'd64576,17'd20602,17'd64577,17'd12716,17'd12415,17'd13514,17'd13364,17'd22647,17'd24542,17'd10992,17'd11809,17'd12116,17'd15688,17'd12116,17'd14674,17'd28583,17'd12588,17'd34040,17'd35371,17'd7954,17'd7955,17'd13893,17'd7458,17'd7956,17'd8586,17'd22300,17'd60101,17'd63738,17'd13008,17'd64578,17'd64312,17'd23875,17'd55708,17'd61748,17'd25007,17'd25007,17'd60830,17'd60830,17'd64579,17'd64580,17'd64581,17'd8430,17'd54463,17'd59193,17'd64582,17'd64583,17'd13143,17'd13655,17'd64584,17'd10349,17'd64585,17'd64586,17'd18928,17'd23533,17'd23533,17'd10621,17'd14692,17'd23533,17'd52880,17'd52146,17'd64587,17'd64588,17'd64589,17'd64590,17'd64591,17'd64592,17'd64593,17'd59574,17'd64594,17'd64595,17'd50645,17'd57325,17'd56967,17'd60842,17'd50646,17'd64596,17'd64326,17'd64192,17'd57708,17'd64326,17'd59085,17'd50814,17'd64597,17'd64053,17'd64598,17'd64330,17'd64599,17'd50813,17'd64056,17'd59456,17'd59456,17'd59990,17'd64057,17'd58824,17'd56507,17'd56507,17'd58334,17'd50730,17'd51074,17'd56285,17'd57967,17'd56285,17'd56285,17'd56285,17'd56285,17'd62797,17'd62797,17'd62797,17'd62797,17'd62797,17'd57076,17'd50156,17'd50156,17'd34282,17'd34459,17'd48987,17'd50364,17'd50363,17'd57205,17'd56285,17'd58823,17'd64600,17'd64601,17'd64602,17'd64603,17'd64206,17'd55967,17'd64604,17'd64605,17'd64606,17'd64478,17'd46095,17'd46095,17'd64607,17'd64608,17'd64481,17'd38029,17'd64609,17'd29999,17'd64610,17'd29399,17'd64611,17'd26088,17'd64612,17'd64613,17'd64614,17'd64615,17'd62810,17'd64616,17'd23421,17'd63632,17'd64617,17'd64618,17'd64619,17'd64358,17'd23241,17'd64620,17'd21259,17'd20345,17'd64621,17'd64622,17'd25071,17'd26577,17'd64623,17'd64501,17'd22740,17'd22392,17'd23622,17'd23971,17'd30793,17'd22934,17'd54410,17'd53504,17'd26584,17'd26448,17'd8608,17'd7008,17'd5323,17'd5324,17'd4994,17'd5609,17'd4843,17'd4843,17'd30637,17'd5008,17'd5010,17'd5011,17'd5013,17'd53426,17'd34923,17'd64624,17'd10239,17'd7332,17'd11319,17'd64625,17'd14429,17'd64626,17'd64627,17'd64628,17'd64629,17'd64630,17'd64631,17'd64508,17'd64632,17'd18506,17'd17177,17'd63944,17'd63944,17'd63944,17'd14432,17'd64509,17'd15230,17'd15861,17'd16622,17'd14172,17'd27431,17'd13288,17'd30643,17'd64633,17'd10787,17'd10069,17'd64634,17'd64634,17'd64635,17'd64636,17'd64513,17'd64637,17'd2882,17'd40257,17'd2714,17'd24319,17'd64382,17'd64638,17'd64639,17'd64640,17'd52529,17'd64641,17'd64642,17'd64643,17'd64644,17'd64645,17'd64646,17'd64524,17'd64647,17'd50843,17'd5939,17'd3246,17'd3897,17'd3897,17'd3423,17'd3423,17'd4085,17'd4713,17'd4714,17'd11061,17'd27949,17'd60625,17'd27822,17'd31410,17'd27822,17'd35770,17'd31251,17'd36905,17'd64648,17'd58865,17'd6094,17'd37959,17'd38203,17'd37958,17'd38202,17'd38580,17'd63959,17'd64649,17'd62697,17'd62969,17'd64526,17'd64650,17'd64387,17'd64387,17'd63655,17'd64651,17'd64652,17'd64109,17'd63658,17'd63657,17'd64388,17'd64653,17'd64654,17'd64655,17'd64656,17'd64532,17'd64657,17'd64658,17'd38855,17'd64533,17'd64534,17'd64659,17'd64391,17'd2215,17'd59623,17'd61033
},
'{
17'd64116,17'd64660,17'd5203,17'd15359,17'd5511,17'd5511,17'd6730,17'd4893,17'd64661,17'd64662,17'd63816,17'd64663,17'd64253,17'd64396,17'd63977,17'd64396,17'd64664,17'd64665,17'd64666,17'd64667,17'd64668,17'd3249,17'd17187,17'd17,17'd3905,17'd4089,17'd4089,17'd3905,17'd17,17'd1415,17'd2596,17'd3429,17'd2934,17'd3427,17'd15358,17'd15358,17'd34512,17'd3251,17'd3427,17'd2934,17'd3751,17'd3901,17'd4086,17'd5511,17'd5511,17'd5511,17'd6730,17'd16392,17'd656,17'd33,17'd12653,17'd14321,17'd63670,17'd43,17'd61286,17'd45,17'd662,17'd50,17'd64669,17'd15366,17'd18151,17'd63672,17'd999,17'd2614,17'd1145,17'd1709,17'd64540,17'd64670,17'd41162,17'd14604,17'd1148,17'd39038,17'd63265,17'd60895,17'd64671,17'd64672,17'd64673,17'd64674,17'd64675,17'd64676,17'd64677,17'd64678,17'd64679,17'd64413,17'd49112,17'd64414,17'd8072,17'd63834,17'd63834,17'd64680,17'd63683,17'd52852,17'd53305,17'd53305,17'd52852,17'd64681,17'd43069,17'd4924,17'd3952,17'd3954,17'd52782,17'd52471,17'd53302,17'd53448,17'd54173,17'd53607,17'd53522,17'd64142,17'd53811,17'd55776,17'd60171,17'd64682,17'd56574,17'd57387,17'd59789,17'd54618,17'd64000,17'd55184,17'd64683,17'd64684,17'd64685,17'd57646,17'd58652,17'd57278,17'd55091,17'd55091,17'd56909,17'd56237,17'd58404,17'd58893,17'd57778,17'd57649,17'd59282,17'd60428,17'd59275,17'd64686,17'd63281,17'd58887,17'd55784,17'd64687,17'd64688,17'd64689,17'd64690,17'd64691,17'd64692,17'd64693,17'd64694,17'd6774,17'd8544,17'd20890,17'd64695,17'd64696,17'd64697,17'd64698,17'd64566,17'd64699,17'd64568,17'd64439,17'd64439,17'd64166,17'd64700,17'd64701,17'd64702,17'd64703,17'd62253,17'd61469,17'd64704,17'd63034,17'd63572,17'd64305,17'd64170,17'd63871,17'd64028,17'd62509,17'd62258,17'd63174,17'd61226,17'd61479,17'd63574,17'd64705,17'd12848,17'd54040,17'd64706,17'd12416,17'd12256,17'd30682,17'd11395,17'd37852,17'd9340,17'd9346,17'd16554,17'd34204,17'd22131,17'd13887,17'd47406,17'd8580,17'd16800,17'd8423,17'd10341,17'd14531,17'd10342,17'd14266,17'd8586,17'd23180,17'd10612,17'd64707,17'd8740,17'd63450,17'd64312,17'd59841,17'd25007,17'd25007,17'd21372,17'd25007,17'd61617,17'd64708,17'd64708,17'd64708,17'd64709,17'd64710,17'd64711,17'd13895,17'd64712,17'd64713,17'd7471,17'd64714,17'd64715,17'd14398,17'd11007,17'd64716,17'd9359,17'd64717,17'd12274,17'd14399,17'd12874,17'd12274,17'd64455,17'd64718,17'd64719,17'd64720,17'd64721,17'd64722,17'd64723,17'd64724,17'd64725,17'd64323,17'd64726,17'd64727,17'd64728,17'd64729,17'd50460,17'd64051,17'd50561,17'd57325,17'd57456,17'd58092,17'd51233,17'd51233,17'd64326,17'd64730,17'd51993,17'd50814,17'd64731,17'd63337,17'd63900,17'd64330,17'd64599,17'd64732,17'd64732,17'd64733,17'd64734,17'd59721,17'd59205,17'd58706,17'd58951,17'd58951,17'd58951,17'd58706,17'd58823,17'd58823,17'd57967,17'd56285,17'd57967,17'd57967,17'd51735,17'd62797,17'd62797,17'd62797,17'd62656,17'd57076,17'd50156,17'd53642,17'd33644,17'd50364,17'd50364,17'd50363,17'd62797,17'd57967,17'd64735,17'd64736,17'd64737,17'd64738,17'd64739,17'd64740,17'd64741,17'd64742,17'd64743,17'd64744,17'd64606,17'd64478,17'd44230,17'd44230,17'd64606,17'd64745,17'd64746,17'd64747,17'd33817,17'd33326,17'd64748,17'd36147,17'd64749,17'd64750,17'd64484,17'd27395,17'd64751,17'd64615,17'd19799,17'd64752,17'd23242,17'd64753,17'd64754,17'd64755,17'd64618,17'd21875,17'd20793,17'd64756,17'd64757,17'd20076,17'd64758,17'd64759,17'd64760,17'd64761,17'd64762,17'd63634,17'd22567,17'd23621,17'd23623,17'd24304,17'd25483,17'd22758,17'd54410,17'd29590,17'd26826,17'd10196,17'd7325,17'd7008,17'd5323,17'd5325,17'd5326,17'd5609,17'd5005,17'd5005,17'd5008,17'd5163,17'd5170,17'd35197,17'd52762,17'd52762,17'd6225,17'd6396,17'd64503,17'd12006,17'd13283,17'd64763,17'd64764,17'd64765,17'd64505,17'd64766,17'd64767,17'd64630,17'd64631,17'd64508,17'd26004,17'd18506,17'd14057,17'd63944,17'd63944,17'd14432,17'd64768,17'd64768,17'd64769,17'd64769,17'd64769,17'd15230,17'd17177,17'd63359,17'd64770,17'd64771,17'd64772,17'd10904,17'd64773,17'd64774,17'd64775,17'd64776,17'd64777,17'd48470,17'd64778,17'd64779,17'd64780,17'd64781,17'd64782,17'd64783,17'd64784,17'd64785,17'd39787,17'd2367,17'd2541,17'd2893,17'd51252,17'd53292,17'd64786,17'd10524,17'd52020,17'd4400,17'd4712,17'd50843,17'd37821,17'd37708,17'd3423,17'd3246,17'd3897,17'd4728,17'd6889,17'd5777,17'd30942,17'd29612,17'd28792,17'd27822,17'd64787,17'd35770,17'd31101,17'd36903,17'd9261,17'd7364,17'd6258,17'd4867,17'd37957,17'd5938,17'd38860,17'd12635,17'd63959,17'd62574,17'd64788,17'd63372,17'd63962,17'd64387,17'd64387,17'd64387,17'd63655,17'd64651,17'd64527,17'd64109,17'd63657,17'd63809,17'd64388,17'd64789,17'd64790,17'd64791,17'd64531,17'd64532,17'd64657,17'd64658,17'd38855,17'd64792,17'd2529,17'd37817,17'd52529,17'd2215,17'd59623,17'd60772
},
'{
17'd64116,17'd64116,17'd5203,17'd15359,17'd5511,17'd5204,17'd6730,17'd4737,17'd64793,17'd64393,17'd64794,17'd63816,17'd64795,17'd63976,17'd63977,17'd64121,17'd64796,17'd64797,17'd64798,17'd64799,17'd10923,17'd3249,17'd17187,17'd17,17'd3905,17'd4089,17'd4089,17'd3905,17'd17,17'd1415,17'd1414,17'd3752,17'd2935,17'd3427,17'd15358,17'd15358,17'd37047,17'd34512,17'd3427,17'd3427,17'd3751,17'd3901,17'd4086,17'd5204,17'd5511,17'd5511,17'd6730,17'd5204,17'd10924,17'd33,17'd12784,17'd58016,17'd14322,17'd63670,17'd43,17'd64401,17'd60036,17'd662,17'd55660,17'd64669,17'd18151,17'd63672,17'd2616,17'd14604,17'd996,17'd1709,17'd64800,17'd64540,17'd41162,17'd15631,17'd2615,17'd999,17'd63265,17'd999,17'd64801,17'd64802,17'd64803,17'd64804,17'd64805,17'd64806,17'd64132,17'd64807,17'd64808,17'd64809,17'd49112,17'd64810,17'd8072,17'd64811,17'd64812,17'd64813,17'd64814,17'd64815,17'd54262,17'd64816,17'd61834,17'd62591,17'd64814,17'd5084,17'd4127,17'd7912,17'd63841,17'd58641,17'd64817,17'd53448,17'd54173,17'd53522,17'd53370,17'd64818,17'd64819,17'd64820,17'd64821,17'd60171,17'd64822,17'd64823,17'd64824,17'd59930,17'd54893,17'd64825,17'd55380,17'd64826,17'd57639,17'd58035,17'd55378,17'd63405,17'd55091,17'd57133,17'd58159,17'd64827,17'd58525,17'd63550,17'd59144,17'd59150,17'd64828,17'd60177,17'd58771,17'd63146,17'd63280,17'd59024,17'd58526,17'd58410,17'd64829,17'd64830,17'd709,17'd64831,17'd64832,17'd64833,17'd64834,17'd5690,17'd7917,17'd13104,17'd20890,17'd14489,17'd64835,17'd64836,17'd64837,17'd64699,17'd64838,17'd64568,17'd64568,17'd64700,17'd64839,17'd64701,17'd64840,17'd64440,17'd64841,17'd61736,17'd64842,17'd64843,17'd64844,17'd64305,17'd64170,17'd64170,17'd63871,17'd64028,17'd62382,17'd63438,17'd61095,17'd59690,17'd63308,17'd64845,17'd14251,17'd56268,17'd64846,17'd12418,17'd12856,17'd64447,17'd15175,17'd19532,17'd15295,17'd9189,17'd25525,17'd25407,17'd24037,17'd9192,17'd50526,17'd11138,17'd8421,17'd57820,17'd20456,17'd14139,17'd15574,17'd12430,17'd14271,17'd10612,17'd64707,17'd61230,17'd62773,17'd64847,17'd16338,17'd61232,17'd60830,17'd25007,17'd59841,17'd61100,17'd64848,17'd21830,17'd64849,17'd64850,17'd64708,17'd64851,17'd56058,17'd61233,17'd11816,17'd64852,17'd64853,17'd64854,17'd22834,17'd64855,17'd52731,17'd12275,17'd12275,17'd18211,17'd12274,17'd64856,17'd11977,17'd18458,17'd64857,17'd64858,17'd64859,17'd64860,17'd64861,17'd64862,17'd64863,17'd64864,17'd64865,17'd64866,17'd64867,17'd64866,17'd64868,17'd64869,17'd64596,17'd60842,17'd50465,17'd57325,17'd52075,17'd64870,17'd64870,17'd64326,17'd64871,17'd64872,17'd58462,17'd59205,17'd58584,17'd59580,17'd64731,17'd64329,17'd64329,17'd63337,17'd64873,17'd64733,17'd64733,17'd64874,17'd58584,17'd59083,17'd58951,17'd58706,17'd64875,17'd64875,17'd50819,17'd50819,17'd52887,17'd57967,17'd56285,17'd57967,17'd62797,17'd57205,17'd57205,17'd62797,17'd62656,17'd57076,17'd57076,17'd33644,17'd50364,17'd62655,17'd62655,17'd57205,17'd56285,17'd51074,17'd64876,17'd64736,17'd64877,17'd64878,17'd64879,17'd64880,17'd64881,17'd64742,17'd64743,17'd64744,17'd61764,17'd64606,17'd43286,17'd53051,17'd64208,17'd64882,17'd64883,17'd64747,17'd33817,17'd28731,17'd64884,17'd23584,17'd60491,17'd64885,17'd64886,17'd64887,17'd64751,17'd64888,17'd64889,17'd26423,17'd64890,17'd64891,17'd64892,17'd64893,17'd64618,17'd22035,17'd64894,17'd64757,17'd20794,17'd64895,17'd18601,17'd18731,17'd64896,17'd23094,17'd64897,17'd54671,17'd23621,17'd56875,17'd23792,17'd30793,17'd11829,17'd54956,17'd64898,17'd10359,17'd9503,17'd10196,17'd6545,17'd7008,17'd5324,17'd5151,17'd5478,17'd4844,17'd5002,17'd30637,17'd5009,17'd5170,17'd37435,17'd52762,17'd52762,17'd9093,17'd9396,17'd64899,17'd11182,17'd13283,17'd64625,17'd64900,17'd64901,17'd64627,17'd64902,17'd64903,17'd64630,17'd64904,17'd64905,17'd64508,17'd26004,17'd18506,17'd14057,17'd63944,17'd14432,17'd14432,17'd64768,17'd64769,17'd64769,17'd64769,17'd63494,17'd64769,17'd64509,17'd63945,17'd63791,17'd11863,17'd11584,17'd64772,17'd64906,17'd5348,17'd3860,17'd64907,17'd3050,17'd64908,17'd64909,17'd64910,17'd64911,17'd22776,17'd24949,17'd64912,17'd52529,17'd64913,17'd2370,17'd53672,17'd51182,17'd64914,17'd51412,17'd53006,17'd64915,17'd18142,17'd38579,17'd5937,17'd5937,17'd4400,17'd5939,17'd37821,17'd37821,17'd3423,17'd4575,17'd5958,17'd4714,17'd5030,17'd29611,17'd64916,17'd27822,17'd35770,17'd64787,17'd64917,17'd37168,17'd64648,17'd58865,17'd14858,17'd13933,17'd38203,17'd5938,17'd39948,17'd39182,17'd64918,17'd62444,17'd62574,17'd64788,17'd63106,17'd64387,17'd64387,17'd64919,17'd64387,17'd63655,17'd64651,17'd64527,17'd63965,17'd63657,17'd64388,17'd64920,17'd64921,17'd64922,17'd64923,17'd64656,17'd64924,17'd64925,17'd64658,17'd2891,17'd64792,17'd2529,17'd41620,17'd64926,17'd2215,17'd59623,17'd60772
},
'{
17'd6730,17'd6730,17'd5203,17'd5203,17'd5511,17'd5511,17'd5204,17'd5204,17'd4893,17'd64117,17'd64927,17'd64928,17'd64928,17'd64121,17'd64121,17'd64928,17'd64929,17'd63978,17'd11070,17'd64667,17'd64930,17'd10668,17'd1414,17'd17,17'd3905,17'd20404,17'd4089,17'd4089,17'd17,17'd17187,17'd1415,17'd2596,17'd3252,17'd3101,17'd3251,17'd34512,17'd34512,17'd34512,17'd3427,17'd3427,17'd3427,17'd3427,17'd3592,17'd15496,17'd5204,17'd5204,17'd6730,17'd5204,17'd10924,17'd11071,17'd12196,17'd12504,17'd14989,17'd15360,17'd63261,17'd61286,17'd60036,17'd662,17'd55660,17'd15248,17'd1981,17'd63672,17'd2616,17'd14196,17'd2614,17'd1290,17'd39038,17'd61289,17'd64931,17'd64932,17'd16266,17'd1148,17'd63673,17'd64800,17'd64933,17'd64934,17'd64935,17'd64936,17'd61825,17'd64937,17'd64938,17'd64939,17'd64940,17'd64941,17'd6778,17'd6938,17'd7755,17'd64811,17'd8847,17'd8073,17'd6778,17'd53376,17'd64416,17'd61053,17'd64816,17'd64942,17'd63135,17'd64943,17'd4127,17'd7252,17'd64944,17'd58267,17'd58642,17'd53233,17'd63139,17'd58028,17'd53232,17'd56343,17'd64945,17'd64946,17'd63845,17'd64821,17'd64419,17'd59516,17'd54799,17'd60171,17'd54893,17'd64947,17'd56020,17'd60171,17'd64553,17'd58152,17'd54890,17'd55378,17'd58159,17'd56132,17'd56450,17'd55486,17'd58404,17'd63550,17'd58042,17'd58526,17'd58657,17'd58890,17'd56453,17'd63550,17'd56810,17'd61190,17'd56807,17'd59939,17'd57280,17'd64948,17'd64949,17'd64950,17'd64951,17'd1599,17'd64952,17'd64953,17'd6778,17'd17818,17'd20890,17'd64954,17'd64955,17'd64956,17'd64957,17'd64567,17'd64958,17'd64839,17'd63866,17'd63866,17'd64958,17'd64959,17'd64960,17'd64301,17'd64961,17'd62133,17'd61468,17'd64962,17'd64963,17'd64964,17'd64965,17'd63870,17'd64966,17'd64967,17'd64443,17'd64968,17'd64969,17'd59829,17'd59970,17'd64970,17'd64971,17'd53973,17'd14128,17'd64972,17'd13760,17'd12575,17'd64973,17'd17236,17'd13370,17'd17600,17'd24039,17'd17964,17'd18195,17'd16318,17'd29919,17'd64974,17'd8256,17'd10747,17'd64975,17'd64976,17'd17133,17'd64977,17'd15063,17'd55125,17'd63044,17'd7798,17'd8266,17'd64847,17'd59841,17'd64978,17'd54468,17'd64979,17'd16452,17'd12432,17'd64980,17'd11537,17'd11537,17'd64981,17'd64982,17'd16452,17'd16924,17'd61232,17'd64983,17'd10866,17'd64984,17'd64985,17'd11975,17'd64986,17'd16458,17'd64987,17'd22664,17'd18211,17'd18928,17'd11977,17'd12275,17'd18211,17'd17616,17'd64988,17'd64989,17'd64990,17'd64991,17'd64992,17'd64993,17'd64994,17'd64995,17'd64996,17'd64997,17'd64998,17'd63895,17'd64999,17'd64880,17'd65000,17'd65001,17'd65002,17'd50734,17'd51553,17'd51553,17'd65003,17'd64872,17'd64730,17'd59207,17'd59861,17'd52502,17'd64597,17'd64731,17'd60113,17'd60113,17'd64873,17'd64873,17'd60113,17'd64597,17'd64597,17'd65004,17'd65004,17'd57564,17'd57564,17'd57564,17'd59205,17'd58706,17'd58706,17'd58823,17'd58823,17'd56285,17'd56285,17'd57967,17'd57967,17'd51735,17'd51735,17'd57706,17'd51735,17'd62797,17'd57839,17'd65005,17'd65005,17'd65006,17'd65007,17'd64876,17'd65008,17'd65009,17'd64877,17'd65010,17'd64879,17'd65011,17'd65012,17'd64881,17'd65013,17'd50562,17'd53487,17'd65014,17'd64208,17'd64208,17'd65015,17'd61764,17'd65016,17'd65017,17'd65018,17'd65019,17'd65020,17'd65021,17'd26071,17'd65022,17'd64484,17'd64887,17'd65023,17'd65024,17'd64888,17'd65025,17'd65026,17'd65027,17'd65028,17'd65029,17'd65030,17'd64620,17'd23241,17'd65031,17'd65028,17'd65032,17'd65033,17'd25611,17'd19705,17'd21297,17'd22407,17'd22391,17'd22567,17'd22931,17'd65034,17'd22933,17'd11984,17'd54309,17'd22759,17'd26327,17'd10627,17'd8608,17'd26449,17'd7008,17'd7008,17'd4993,17'd5150,17'd5150,17'd4843,17'd5005,17'd5004,17'd5166,17'd5170,17'd37435,17'd8473,17'd8305,17'd8782,17'd10518,17'd12006,17'd12006,17'd13284,17'd13927,17'd65035,17'd65036,17'd65037,17'd65038,17'd65039,17'd64630,17'd65040,17'd15482,17'd64508,17'd18506,17'd26004,17'd14432,17'd63790,17'd25488,17'd64768,17'd64769,17'd63494,17'd65041,17'd65041,17'd63495,17'd63639,17'd65042,17'd65043,17'd65044,17'd65045,17'd65046,17'd65047,17'd3860,17'd4549,17'd47669,17'd65048,17'd65049,17'd65050,17'd37301,17'd65051,17'd65052,17'd64781,17'd62707,17'd63812,17'd52529,17'd64785,17'd2220,17'd55654,17'd51016,17'd52019,17'd3703,17'd53006,17'd54014,17'd59619,17'd5496,17'd38717,17'd4558,17'd4558,17'd5938,17'd37821,17'd37821,17'd4575,17'd5789,17'd6581,17'd5183,17'd36602,17'd29612,17'd64916,17'd65053,17'd35770,17'd31900,17'd36906,17'd36905,17'd38460,17'd7364,17'd16623,17'd4867,17'd37957,17'd37957,17'd41481,17'd13056,17'd62445,17'd62444,17'd15862,17'd62848,17'd63962,17'd64387,17'd64387,17'd65054,17'd65054,17'd64651,17'd64651,17'd64527,17'd63965,17'd63657,17'd63809,17'd65055,17'd65056,17'd64529,17'd64530,17'd65057,17'd65058,17'd65059,17'd46594,17'd2892,17'd64792,17'd65060,17'd41620,17'd65061,17'd65062,17'd57482,17'd60772
},
'{
17'd6730,17'd6730,17'd6730,17'd5203,17'd5511,17'd5511,17'd5204,17'd5204,17'd4086,17'd64251,17'd65063,17'd65064,17'd64928,17'd63977,17'd64121,17'd65065,17'd65066,17'd65067,17'd65068,17'd65068,17'd12783,17'd63386,17'd2936,17'd1416,17'd3905,17'd4089,17'd4089,17'd1416,17'd1415,17'd1415,17'd1414,17'd1414,17'd3252,17'd2935,17'd3251,17'd3251,17'd34512,17'd34512,17'd3427,17'd3427,17'd3427,17'd3427,17'd3592,17'd15496,17'd5204,17'd5204,17'd6730,17'd5204,17'd10925,17'd10924,17'd11071,17'd11888,17'd58016,17'd14322,17'd63261,17'd65069,17'd61286,17'd60036,17'd50,17'd55660,17'd15366,17'd62861,17'd672,17'd65070,17'd14604,17'd1290,17'd39038,17'd64402,17'd63266,17'd64932,17'd16266,17'd38867,17'd39038,17'd63673,17'd61168,17'd65071,17'd65072,17'd65073,17'd62083,17'd65074,17'd64938,17'd65075,17'd65076,17'd65077,17'd64809,17'd6778,17'd7755,17'd8073,17'd8220,17'd8074,17'd7261,17'd6636,17'd65078,17'd60904,17'd53305,17'd53884,17'd65079,17'd63681,17'd44521,17'd7252,17'd4611,17'd8539,17'd58762,17'd64817,17'd58396,17'd54094,17'd53232,17'd56343,17'd58648,17'd57382,17'd54093,17'd65080,17'd65081,17'd59516,17'd64682,17'd64283,17'd54992,17'd64947,17'd65082,17'd54618,17'd54529,17'd56904,17'd57508,17'd57395,17'd57277,17'd57277,17'd58035,17'd57390,17'd62474,17'd58651,17'd64004,17'd59275,17'd63848,17'd63407,17'd56578,17'd59024,17'd56810,17'd63003,17'd58771,17'd60183,17'd65083,17'd65084,17'd65085,17'd58285,17'd65086,17'd65087,17'd65088,17'd65089,17'd6774,17'd65090,17'd10125,17'd21658,17'd65091,17'd65092,17'd65093,17'd65094,17'd65095,17'd65096,17'd65097,17'd65098,17'd64839,17'd65099,17'd65100,17'd65101,17'd65102,17'd65103,17'd63170,17'd65104,17'd65105,17'd64964,17'd64965,17'd65106,17'd65107,17'd65108,17'd64028,17'd63035,17'd61742,17'd60699,17'd65109,17'd65110,17'd65111,17'd65112,17'd17961,17'd65113,17'd13518,17'd12575,17'd14808,17'd15432,17'd10169,17'd53474,17'd8873,17'd65114,17'd15180,17'd9347,17'd8723,17'd61099,17'd8106,17'd65115,17'd13771,17'd65116,17'd55322,17'd15309,17'd23526,17'd23875,17'd8266,17'd8266,17'd8266,17'd8266,17'd59841,17'd64978,17'd16924,17'd16452,17'd60232,17'd11284,17'd65117,17'd65118,17'd65118,17'd21993,17'd65119,17'd15065,17'd65120,17'd58810,17'd65121,17'd9627,17'd7475,17'd65122,17'd14541,17'd16458,17'd23536,17'd65123,17'd65124,17'd22664,17'd18211,17'd18211,17'd8444,17'd13899,17'd65125,17'd65126,17'd65127,17'd65128,17'd65129,17'd65130,17'd65131,17'd65132,17'd65133,17'd65134,17'd64865,17'd65135,17'd65136,17'd65137,17'd65011,17'd64206,17'd57199,17'd65002,17'd57456,17'd58092,17'd65138,17'd65139,17'd59085,17'd59085,17'd59207,17'd51993,17'd65004,17'd52502,17'd65004,17'd64874,17'd64597,17'd60113,17'd64731,17'd58708,17'd58708,17'd58463,17'd65004,17'd65004,17'd59205,17'd59205,17'd59205,17'd59205,17'd58706,17'd58706,17'd50819,17'd58823,17'd56285,17'd56285,17'd56285,17'd57967,17'd62797,17'd57205,17'd62797,17'd57205,17'd57205,17'd50563,17'd65006,17'd65006,17'd65007,17'd65008,17'd65140,17'd65009,17'd64877,17'd64878,17'd64739,17'd64879,17'd65011,17'd64880,17'd65141,17'd65142,17'd52425,17'd53841,17'd64744,17'd65143,17'd65015,17'd61764,17'd65144,17'd65145,17'd65146,17'd28375,17'd65147,17'd65148,17'd65149,17'd65150,17'd65151,17'd64613,17'd65023,17'd63217,17'd63079,17'd65152,17'd26309,17'd65153,17'd21414,17'd20794,17'd65154,17'd65155,17'd64358,17'd64620,17'd21101,17'd65156,17'd65157,17'd65158,17'd17770,17'd65159,17'd23966,17'd22564,17'd22928,17'd23097,17'd65034,17'd55643,17'd24643,17'd26583,17'd22587,17'd8912,17'd30330,17'd10627,17'd26449,17'd26449,17'd7008,17'd26827,17'd5480,17'd5150,17'd25770,17'd4843,17'd30637,17'd5165,17'd5170,17'd37435,17'd8474,17'd8305,17'd8157,17'd8634,17'd11319,17'd13283,17'd13411,17'd16375,17'd65160,17'd65161,17'd65162,17'd65163,17'd65164,17'd65039,17'd64507,17'd63789,17'd15482,17'd64508,17'd17177,17'd18379,17'd64768,17'd63790,17'd25488,17'd64768,17'd64769,17'd63494,17'd65041,17'd65165,17'd63639,17'd63639,17'd65042,17'd65166,17'd18381,17'd65167,17'd65168,17'd65169,17'd8010,17'd3374,17'd65170,17'd65171,17'd65172,17'd65173,17'd65174,17'd65175,17'd65176,17'd65177,17'd23125,17'd62980,17'd34341,17'd65178,17'd2371,17'd55654,17'd53870,17'd51581,17'd4552,17'd5493,17'd39179,17'd18383,17'd5355,17'd38579,17'd5937,17'd4558,17'd5938,17'd37957,17'd37708,17'd4883,17'd5958,17'd6416,17'd11061,17'd35207,17'd60625,17'd64916,17'd65053,17'd64917,17'd65179,17'd65180,17'd64648,17'd58865,17'd14858,17'd13176,17'd12636,17'd38334,17'd38334,17'd38580,17'd62445,17'd62445,17'd62574,17'd64788,17'd63372,17'd63807,17'd64387,17'd64387,17'd65181,17'd65181,17'd64651,17'd65182,17'd64109,17'd64110,17'd63809,17'd64921,17'd64921,17'd64921,17'd64654,17'd64655,17'd65183,17'd65058,17'd65059,17'd46594,17'd2892,17'd65184,17'd65060,17'd41620,17'd65185,17'd65062,17'd57482,17'd60772
},
'{
17'd5204,17'd5204,17'd5204,17'd5204,17'd15496,17'd15877,17'd15877,17'd15877,17'd3592,17'd4738,17'd65186,17'd64927,17'd65187,17'd65065,17'd64795,17'd63977,17'd65188,17'd65067,17'd65189,17'd65189,17'd63668,17'd10923,17'd14742,17'd14,17'd3905,17'd4089,17'd4089,17'd1416,17'd1415,17'd1415,17'd17,17'd1414,17'd2258,17'd52621,17'd10547,17'd12195,17'd34512,17'd34512,17'd3427,17'd3427,17'd2934,17'd3427,17'd3901,17'd3592,17'd5204,17'd5511,17'd5203,17'd5203,17'd3901,17'd2934,17'd11071,17'd12505,17'd16392,17'd15629,17'd15243,17'd65069,17'd61286,17'd44,17'd56671,17'd55568,17'd14872,17'd18151,17'd672,17'd65070,17'd2441,17'd2615,17'd2950,17'd62080,17'd2794,17'd64932,17'd2442,17'd2951,17'd998,17'd54880,17'd65190,17'd65191,17'd65192,17'd65193,17'd65194,17'd65195,17'd65196,17'd65197,17'd65198,17'd65199,17'd65200,17'd7098,17'd8070,17'd8073,17'd8379,17'd25803,17'd7101,17'd6779,17'd65201,17'd6318,17'd54262,17'd53305,17'd64416,17'd63135,17'd64943,17'd3952,17'd8066,17'd8066,17'd58644,17'd52471,17'd53302,17'd58396,17'd53370,17'd56343,17'd56343,17'd57382,17'd58647,17'd54532,17'd64821,17'd64419,17'd64283,17'd64283,17'd65202,17'd54893,17'd65203,17'd54433,17'd65204,17'd65205,17'd64553,17'd57639,17'd65206,17'd57277,17'd55282,17'd65207,17'd58282,17'd57921,17'd62474,17'd57515,17'd60663,17'd65208,17'd58657,17'd64557,17'd57512,17'd57512,17'd59275,17'd58771,17'd59145,17'd60542,17'd62230,17'd62734,17'd65209,17'd65210,17'd65211,17'd65212,17'd5690,17'd65213,17'd9444,17'd23157,17'd65214,17'd65215,17'd65216,17'd65094,17'd65217,17'd65096,17'd65097,17'd65218,17'd65219,17'd65100,17'd65220,17'd65221,17'd63719,17'd62901,17'd62758,17'd65222,17'd65105,17'd65223,17'd64965,17'd65106,17'd65107,17'd65108,17'd64028,17'd62382,17'd65224,17'd65225,17'd65226,17'd65227,17'd65228,17'd15423,17'd26751,17'd62262,17'd42948,17'd13763,17'd13363,17'd65229,17'd12863,17'd65230,17'd8566,17'd11810,17'd15180,17'd12117,17'd8881,17'd65231,17'd53476,17'd7957,17'd14143,17'd15446,17'd15577,17'd59841,17'd61232,17'd61232,17'd12731,17'd61617,17'd11536,17'd64312,17'd59841,17'd64978,17'd16452,17'd60232,17'd65232,17'd56171,17'd65233,17'd65234,17'd65235,17'd65236,17'd65237,17'd15198,17'd65238,17'd65239,17'd12124,17'd12733,17'd65240,17'd7809,17'd65241,17'd53258,17'd21375,17'd13900,17'd13899,17'd22664,17'd18211,17'd14275,17'd8444,17'd52960,17'd65242,17'd65243,17'd65244,17'd65245,17'd65246,17'd65247,17'd65248,17'd65249,17'd65250,17'd65251,17'd65251,17'd65252,17'd65253,17'd65254,17'd65255,17'd64603,17'd65256,17'd65257,17'd50729,17'd65258,17'd65259,17'd64601,17'd58462,17'd59207,17'd58329,17'd58462,17'd51993,17'd59206,17'd59206,17'd58584,17'd58584,17'd65004,17'd65004,17'd58463,17'd65004,17'd65004,17'd65004,17'd65004,17'd59205,17'd59205,17'd59206,17'd59206,17'd58706,17'd58706,17'd58706,17'd58951,17'd51074,17'd51074,17'd51074,17'd51074,17'd56285,17'd56285,17'd65006,17'd65006,17'd65260,17'd65261,17'd65261,17'd65262,17'd65262,17'd65263,17'd65264,17'd65265,17'd65266,17'd65267,17'd64879,17'd64879,17'd59085,17'd65258,17'd50646,17'd52162,17'd65268,17'd65269,17'd52967,17'd64605,17'd65270,17'd65271,17'd65272,17'd64882,17'd65273,17'd32682,17'd30896,17'd28139,17'd25445,17'd23055,17'd20790,17'd27540,17'd65274,17'd65275,17'd65276,17'd65025,17'd65277,17'd21561,17'd20345,17'd65278,17'd65154,17'd65279,17'd64756,17'd21259,17'd20794,17'd19949,17'd19440,17'd65280,17'd18364,17'd65281,17'd53137,17'd22218,17'd22392,17'd23620,17'd65034,17'd54593,17'd26111,17'd26327,17'd22587,17'd8608,17'd10359,17'd10197,17'd26449,17'd26449,17'd26827,17'd26827,17'd5480,17'd5150,17'd5005,17'd5005,17'd5009,17'd5165,17'd5170,17'd65282,17'd8473,17'd8156,17'd8157,17'd13409,17'd13283,17'd64625,17'd13285,17'd15995,17'd65283,17'd65284,17'd65285,17'd64902,17'd64767,17'd65286,17'd63789,17'd63788,17'd65287,17'd65288,17'd14172,17'd25091,17'd63495,17'd64370,17'd63495,17'd63495,17'd64769,17'd63494,17'd64089,17'd64227,17'd65289,17'd63789,17'd15998,17'd65290,17'd18508,17'd65291,17'd65292,17'd65293,17'd65294,17'd47569,17'd65295,17'd65296,17'd65297,17'd65298,17'd63649,17'd59241,17'd63802,17'd64238,17'd65299,17'd65300,17'd65301,17'd65302,17'd65303,17'd2224,17'd41770,17'd41158,17'd6081,17'd40411,17'd39179,17'd38858,17'd58626,17'd38579,17'd38333,17'd5356,17'd37957,17'd5028,17'd4867,17'd4730,17'd6581,17'd5183,17'd27949,17'd31251,17'd64916,17'd64916,17'd64917,17'd64917,17'd60030,17'd65180,17'd38460,17'd7878,17'd16623,17'd13420,17'd5028,17'd38202,17'd41481,17'd60399,17'd13056,17'd65304,17'd15862,17'd62848,17'd63106,17'd64387,17'd64387,17'd65181,17'd65181,17'd65181,17'd65182,17'd65305,17'd64109,17'd65306,17'd64653,17'd65055,17'd64388,17'd65307,17'd64790,17'd64791,17'd65308,17'd65058,17'd65059,17'd46594,17'd3056,17'd65184,17'd65060,17'd41620,17'd64913,17'd65062,17'd57482,17'd65309
},
'{
17'd5204,17'd5204,17'd5204,17'd5204,17'd15496,17'd15877,17'd15877,17'd61679,17'd3592,17'd3901,17'd65310,17'd65311,17'd65187,17'd64928,17'd65312,17'd63977,17'd65188,17'd65067,17'd63978,17'd63978,17'd65313,17'd63668,17'd65314,17'd14742,17'd17187,17'd1416,17'd1416,17'd1415,17'd17187,17'd17187,17'd16,17'd17,17'd1414,17'd2258,17'd52621,17'd12195,17'd34512,17'd34512,17'd3427,17'd3427,17'd3427,17'd3427,17'd3901,17'd3592,17'd5204,17'd5203,17'd15117,17'd15359,17'd15496,17'd3427,17'd2934,17'd10924,17'd11888,17'd15118,17'd15360,17'd63261,17'd43,17'd44,17'd818,17'd51,17'd14750,17'd2791,17'd670,17'd65070,17'd2125,17'd15631,17'd1709,17'd62212,17'd61289,17'd2618,17'd65315,17'd2619,17'd23659,17'd54880,17'd65316,17'd65317,17'd65318,17'd65319,17'd65320,17'd65321,17'd65322,17'd65323,17'd65324,17'd64270,17'd61174,17'd65325,17'd8070,17'd7422,17'd8379,17'd8378,17'd7757,17'd7422,17'd64809,17'd63135,17'd61835,17'd53166,17'd62093,17'd64815,17'd63681,17'd4126,17'd7252,17'd4611,17'd58267,17'd58641,17'd53018,17'd53081,17'd56572,17'd56343,17'd56343,17'd53370,17'd58519,17'd53757,17'd65080,17'd59789,17'd64682,17'd64283,17'd65202,17'd55185,17'd65203,17'd65326,17'd65327,17'd65328,17'd54799,17'd65329,17'd65330,17'd63278,17'd65331,17'd58152,17'd54990,17'd58652,17'd65332,17'd62878,17'd65333,17'd65334,17'd58890,17'd65335,17'd57391,17'd59523,17'd59280,17'd63550,17'd56453,17'd58771,17'd59024,17'd59279,17'd65336,17'd65337,17'd65338,17'd65339,17'd2657,17'd65340,17'd15783,17'd10290,17'd20596,17'd65341,17'd65342,17'd65343,17'd65344,17'd65345,17'd65097,17'd65098,17'd65346,17'd65346,17'd65220,17'd65100,17'd64166,17'd63433,17'd62622,17'd65347,17'd65348,17'd64573,17'd65349,17'd65106,17'd64170,17'd65107,17'd63871,17'd62509,17'd64968,17'd63037,17'd65350,17'd62765,17'd57680,17'd17225,17'd11951,17'd65351,17'd12410,17'd12419,17'd12857,17'd50423,17'd15052,17'd36630,17'd11530,17'd15178,17'd10174,17'd10174,17'd8881,17'd61099,17'd65352,17'd8428,17'd65353,17'd65354,17'd65355,17'd62636,17'd8590,17'd12731,17'd8590,17'd61232,17'd65356,17'd12269,17'd61617,17'd16452,17'd65120,17'd16573,17'd12124,17'd65357,17'd65358,17'd65359,17'd62516,17'd65360,17'd11409,17'd14820,17'd52653,17'd13774,17'd12125,17'd22833,17'd10350,17'd9755,17'd65361,17'd20622,17'd15823,17'd13900,17'd13899,17'd13899,17'd14275,17'd14275,17'd14276,17'd14016,17'd52884,17'd65362,17'd65363,17'd65364,17'd65365,17'd65366,17'd65367,17'd65368,17'd65369,17'd65370,17'd64462,17'd65371,17'd65372,17'd65373,17'd65266,17'd65374,17'd65375,17'd65012,17'd59722,17'd57456,17'd64061,17'd65008,17'd58951,17'd65376,17'd59861,17'd58462,17'd64468,17'd51993,17'd65377,17'd57564,17'd58584,17'd52502,17'd65378,17'd59083,17'd59206,17'd59206,17'd65004,17'd58584,17'd59206,17'd59206,17'd59206,17'd59206,17'd58706,17'd58706,17'd59454,17'd59454,17'd50730,17'd50730,17'd50730,17'd50730,17'd50563,17'd50563,17'd65379,17'd65379,17'd65379,17'd65380,17'd65380,17'd65381,17'd65381,17'd65382,17'd65383,17'd65384,17'd65385,17'd65386,17'd65387,17'd65388,17'd65258,17'd57708,17'd57708,17'd50646,17'd65389,17'd65390,17'd64743,17'd65391,17'd65392,17'd65271,17'd65393,17'd65394,17'd31364,17'd61117,17'd28737,17'd65395,17'd23058,17'd65396,17'd65397,17'd65398,17'd65399,17'd65400,17'd65401,17'd65402,17'd65403,17'd65404,17'd20794,17'd65405,17'd65406,17'd65407,17'd65031,17'd64757,17'd65408,17'd65409,17'd65410,17'd65411,17'd24634,17'd65412,17'd65413,17'd22565,17'd23621,17'd22931,17'd62681,17'd24943,17'd26215,17'd26448,17'd10196,17'd9503,17'd52521,17'd10197,17'd26449,17'd26449,17'd26827,17'd26827,17'd5480,17'd5150,17'd5005,17'd30637,17'd5165,17'd53794,17'd65414,17'd8474,17'd8305,17'd8157,17'd8634,17'd13282,17'd13284,17'd16375,17'd65415,17'd65416,17'd65417,17'd65418,17'd64505,17'd65419,17'd64767,17'd64630,17'd63640,17'd63495,17'd65288,17'd63495,17'd64768,17'd64768,17'd65420,17'd65420,17'd63495,17'd63495,17'd64769,17'd65041,17'd64227,17'd65289,17'd64369,17'd65421,17'd63942,17'd15998,17'd17414,17'd65422,17'd65423,17'd65424,17'd65425,17'd47380,17'd65426,17'd65427,17'd65428,17'd65429,17'd65430,17'd65431,17'd65432,17'd65433,17'd65434,17'd65435,17'd65436,17'd64785,17'd65437,17'd65438,17'd61281,17'd3562,17'd7849,17'd48811,17'd18512,17'd5354,17'd5180,17'd38579,17'd38333,17'd38201,17'd37957,17'd12636,17'd13933,17'd6258,17'd6416,17'd11061,17'd36905,17'd60625,17'd64916,17'd63652,17'd65179,17'd65439,17'd65180,17'd65440,17'd7878,17'd14858,17'd13176,17'd44019,17'd38334,17'd39033,17'd12176,17'd13056,17'd62445,17'd14735,17'd64788,17'd63372,17'd64387,17'd64919,17'd65054,17'd65054,17'd65054,17'd65054,17'd65182,17'd65305,17'd64110,17'd65306,17'd64921,17'd65055,17'd64921,17'd64653,17'd64922,17'd64923,17'd65441,17'd64924,17'd65059,17'd65442,17'd3056,17'd65443,17'd65444,17'd41620,17'd64913,17'd65445,17'd58367,17'd65309
},
'{
17'd5204,17'd5204,17'd5204,17'd4086,17'd5204,17'd5204,17'd15877,17'd61679,17'd15496,17'd3901,17'd6892,17'd65446,17'd65064,17'd64928,17'd65312,17'd64253,17'd65447,17'd65448,17'd64537,17'd65449,17'd64254,17'd63979,17'd14441,17'd63258,17'd65450,17'd2257,17'd2257,17'd1415,17'd1415,17'd17187,17'd1277,17'd17,17'd1414,17'd2597,17'd3429,17'd10547,17'd10670,17'd10670,17'd3251,17'd3251,17'd3251,17'd3251,17'd3428,17'd3592,17'd5204,17'd5511,17'd5203,17'd5203,17'd4891,17'd3592,17'd2934,17'd11071,17'd12505,17'd472,17'd14599,17'd59774,17'd65451,17'd44,17'd818,17'd301,17'd14750,17'd2791,17'd837,17'd65070,17'd2125,17'd16145,17'd1710,17'd65452,17'd54787,17'd836,17'd2792,17'd2619,17'd2951,17'd62080,17'd65453,17'd61168,17'd65454,17'd65455,17'd65456,17'd65457,17'd65458,17'd65459,17'd65460,17'd65461,17'd64133,17'd65462,17'd64813,17'd7422,17'd8377,17'd8379,17'd8379,17'd8074,17'd8070,17'd6937,17'd53375,17'd61964,17'd65463,17'd43470,17'd65464,17'd5083,17'd4464,17'd64944,17'd63996,17'd65465,17'd65466,17'd53018,17'd52851,17'd56686,17'd53232,17'd53232,17'd58519,17'd65467,17'd65468,17'd57126,17'd65469,17'd56233,17'd54992,17'd56020,17'd65470,17'd54532,17'd54434,17'd63845,17'd65471,17'd56234,17'd65472,17'd65473,17'd64282,17'd60539,17'd63141,17'd60656,17'd58772,17'd57275,17'd64686,17'd63548,17'd65474,17'd60177,17'd58887,17'd65475,17'd59017,17'd1459,17'd59517,17'd61441,17'd58768,17'd61449,17'd65476,17'd65477,17'd65478,17'd65479,17'd65480,17'd65481,17'd65482,17'd10125,17'd65483,17'd65484,17'd65485,17'd65486,17'd65487,17'd65488,17'd65489,17'd65098,17'd65346,17'd65346,17'd65490,17'd65100,17'd64700,17'd63569,17'd65491,17'd63170,17'd65492,17'd64963,17'd65493,17'd65106,17'd64170,17'd64170,17'd63871,17'd64028,17'd62258,17'd60573,17'd65494,17'd65495,17'd65496,17'd13242,17'd11652,17'd11263,17'd21203,17'd12113,17'd12999,17'd17598,17'd21986,17'd11276,17'd41655,17'd15296,17'd8880,17'd39660,17'd8725,17'd25678,17'd9746,17'd65497,17'd65498,17'd65499,17'd65500,17'd8432,17'd13143,17'd8590,17'd21062,17'd12731,17'd59841,17'd61232,17'd8590,17'd65501,17'd13655,17'd12596,17'd25009,17'd12125,17'd10868,17'd65502,17'd65503,17'd24053,17'd11972,17'd16925,17'd65504,17'd65505,17'd14398,17'd13260,17'd8750,17'd9359,17'd7980,17'd16090,17'd11413,17'd14276,17'd14016,17'd8131,17'd9059,17'd9059,17'd14016,17'd23536,17'd24056,17'd21681,17'd65506,17'd65507,17'd65508,17'd64861,17'd65509,17'd61490,17'd65132,17'd64724,17'd65510,17'd65511,17'd65512,17'd65513,17'd65514,17'd65515,17'd64878,17'd65516,17'd65375,17'd65256,17'd65375,17'd65008,17'd65517,17'd65262,17'd64601,17'd64474,17'd59861,17'd58462,17'd59861,17'd65376,17'd57564,17'd59206,17'd59083,17'd59083,17'd58706,17'd59206,17'd58584,17'd58584,17'd59206,17'd59083,17'd59083,17'd59083,17'd59083,17'd59083,17'd59454,17'd59454,17'd58824,17'd58824,17'd58824,17'd58824,17'd56507,17'd57455,17'd65518,17'd65518,17'd65518,17'd65519,17'd65519,17'd65520,17'd65521,17'd65522,17'd65523,17'd59078,17'd65524,17'd65386,17'd58461,17'd65003,17'd64326,17'd57708,17'd50734,17'd57325,17'd65525,17'd65390,17'd49786,17'd64743,17'd65526,17'd65527,17'd65528,17'd65529,17'd32515,17'd65530,17'd65531,17'd65532,17'd23231,17'd65533,17'd65534,17'd65535,17'd65399,17'd65536,17'd65537,17'd65538,17'd65539,17'd65540,17'd65408,17'd65541,17'd65154,17'd65542,17'd20345,17'd21563,17'd65543,17'd65544,17'd65545,17'd19322,17'd20373,17'd24297,17'd22390,17'd57220,17'd23620,17'd22756,17'd53503,17'd25081,17'd26584,17'd30330,17'd8608,17'd7165,17'd52521,17'd10197,17'd7164,17'd7008,17'd26827,17'd26827,17'd5150,17'd5150,17'd5005,17'd5004,17'd5165,17'd53794,17'd65282,17'd8474,17'd8157,17'd7331,17'd65546,17'd65547,17'd15994,17'd65415,17'd65548,17'd65549,17'd65550,17'd65551,17'd65552,17'd64766,17'd64629,17'd65553,17'd65042,17'd65288,17'd63495,17'd63495,17'd63495,17'd65554,17'd65420,17'd65420,17'd63495,17'd65555,17'd65555,17'd65041,17'd64227,17'd65289,17'd65421,17'd65040,17'd65556,17'd15347,17'd65557,17'd65558,17'd65559,17'd65560,17'd65561,17'd65562,17'd42781,17'd42645,17'd64659,17'd63971,17'd63661,17'd65428,17'd63515,17'd63515,17'd65436,17'd52454,17'd37953,17'd2538,17'd51015,17'd2725,17'd41479,17'd41480,17'd7849,17'd4056,17'd39179,17'd65563,17'd5495,17'd5026,17'd5356,17'd38201,17'd5028,17'd12914,17'd4730,17'd6094,17'd8187,17'd11882,17'd60030,17'd64917,17'd65564,17'd64917,17'd60030,17'd65439,17'd59125,17'd58865,17'd44850,17'd16855,17'd13420,17'd38580,17'd38860,17'd39182,17'd12635,17'd65565,17'd65304,17'd62575,17'd62699,17'd65566,17'd65567,17'd64919,17'd65054,17'd65054,17'd65568,17'd65569,17'd65305,17'd65570,17'd64110,17'd64241,17'd64921,17'd65055,17'd64921,17'd64653,17'd64922,17'd64923,17'd65571,17'd65572,17'd64925,17'd64658,17'd3056,17'd52099,17'd65573,17'd41620,17'd65574,17'd65445,17'd58367,17'd65575
},
'{
17'd5204,17'd5204,17'd4086,17'd4086,17'd4086,17'd5204,17'd15877,17'd15877,17'd15496,17'd3901,17'd65576,17'd65577,17'd65578,17'd65312,17'd63975,17'd65579,17'd65580,17'd65580,17'd65581,17'd65582,17'd65583,17'd11885,17'd6594,17'd64930,17'd65584,17'd2597,17'd2597,17'd2936,17'd1414,17'd17,17'd18,17'd3905,17'd17,17'd1414,17'd2258,17'd52621,17'd10802,17'd10670,17'd3251,17'd3251,17'd3251,17'd3251,17'd3428,17'd15496,17'd5204,17'd5203,17'd15117,17'd15117,17'd4426,17'd4243,17'd3427,17'd2935,17'd10924,17'd295,17'd15362,17'd59911,17'd65585,17'd61286,17'd58505,17'd302,17'd14991,17'd2791,17'd18151,17'd487,17'd2269,17'd16145,17'd996,17'd41628,17'd61554,17'd54787,17'd65586,17'd40103,17'd23659,17'd62080,17'd63265,17'd60522,17'd63122,17'd65587,17'd65588,17'd65589,17'd65590,17'd65591,17'd65592,17'd65593,17'd63274,17'd65594,17'd8072,17'd7756,17'd7756,17'd8071,17'd65595,17'd8847,17'd7422,17'd7421,17'd53376,17'd43602,17'd65596,17'd65597,17'd62874,17'd63134,17'd5408,17'd63842,17'd65598,17'd65599,17'd65465,17'd65466,17'd57769,17'd59142,17'd56686,17'd53232,17'd58519,17'd65600,17'd65601,17'd63845,17'd65602,17'd56021,17'd54992,17'd56021,17'd56344,17'd54171,17'd54093,17'd58272,17'd65603,17'd65604,17'd65469,17'd64682,17'd65605,17'd65606,17'd54702,17'd58152,17'd55783,17'd65607,17'd57275,17'd59396,17'd63548,17'd63695,17'd59144,17'd1460,17'd65608,17'd58154,17'd59517,17'd61441,17'd57512,17'd60428,17'd60057,17'd59282,17'd65609,17'd65610,17'd65611,17'd65612,17'd65613,17'd9992,17'd65483,17'd65614,17'd65615,17'd65486,17'd65487,17'd65616,17'd65489,17'd64569,17'd65100,17'd65346,17'd65490,17'd65617,17'd65099,17'd64439,17'd63720,17'd62758,17'd65618,17'd65619,17'd65223,17'd64965,17'd64170,17'd64170,17'd63871,17'd64028,17'd62509,17'd63174,17'd59966,17'd65620,17'd65621,17'd65622,17'd12712,17'd11389,17'd65623,17'd11957,17'd11957,17'd12262,17'd23338,17'd65624,17'd29333,17'd34958,17'd65625,17'd56731,17'd8572,17'd25679,17'd15060,17'd65626,17'd65627,17'd65628,17'd61232,17'd59841,17'd61617,17'd61232,17'd21062,17'd12870,17'd13530,17'd61232,17'd8432,17'd65629,17'd15310,17'd65630,17'd65631,17'd65632,17'd22834,17'd12272,17'd65633,17'd65634,17'd65357,17'd13656,17'd16216,17'd14398,17'd13260,17'd12126,17'd12275,17'd8132,17'd133,17'd133,17'd8132,17'd11289,17'd9059,17'd6529,17'd9059,17'd11289,17'd13901,17'd21375,17'd20628,17'd65635,17'd65636,17'd65637,17'd65638,17'd65639,17'd65640,17'd65641,17'd65642,17'd65643,17'd64591,17'd65644,17'd65645,17'd65646,17'd65647,17'd65383,17'd65648,17'd65010,17'd64740,17'd65649,17'd65375,17'd64600,17'd65650,17'd65651,17'd65262,17'd65008,17'd65378,17'd59205,17'd57564,17'd57564,17'd65377,17'd57564,17'd59205,17'd59205,17'd58706,17'd58706,17'd59083,17'd52502,17'd59083,17'd59083,17'd65378,17'd65378,17'd65378,17'd65378,17'd59454,17'd59454,17'd58824,17'd60480,17'd58822,17'd53192,17'd59453,17'd56751,17'd65652,17'd65652,17'd65652,17'd65653,17'd65520,17'd65654,17'd65655,17'd65656,17'd59199,17'd59448,17'd65657,17'd64869,17'd50645,17'd64871,17'd51233,17'd51233,17'd50734,17'd50734,17'd65141,17'd65658,17'd50561,17'd65659,17'd65526,17'd65660,17'd36564,17'd65661,17'd60723,17'd34887,17'd65662,17'd65663,17'd63343,17'd65664,17'd62945,17'd65665,17'd65666,17'd65667,17'd65668,17'd65669,17'd64891,17'd20483,17'd65670,17'd65671,17'd65672,17'd65028,17'd65673,17'd65156,17'd65409,17'd65674,17'd65675,17'd65676,17'd25982,17'd47847,17'd23617,17'd56530,17'd54860,17'd24141,17'd47848,17'd29426,17'd29427,17'd65677,17'd7164,17'd7327,17'd52521,17'd7164,17'd24480,17'd24480,17'd6547,17'd6547,17'd5150,17'd4843,17'd5004,17'd5004,17'd5165,17'd5170,17'd65282,17'd8305,17'd8157,17'd11433,17'd65678,17'd65679,17'd65680,17'd65548,17'd65681,17'd65682,17'd65284,17'd65683,17'd65419,17'd64369,17'd65684,17'd64090,17'd65288,17'd64509,17'd64768,17'd64769,17'd65685,17'd65686,17'd63640,17'd63639,17'd63495,17'd65555,17'd65555,17'd65041,17'd64227,17'd65687,17'd65421,17'd65688,17'd65040,17'd65689,17'd14857,17'd65690,17'd65691,17'd65692,17'd3697,17'd65693,17'd65694,17'd65695,17'd65696,17'd65697,17'd65698,17'd40857,17'd40857,17'd40559,17'd51935,17'd65699,17'd3057,17'd3059,17'd41903,17'd41623,17'd41905,17'd42043,17'd4055,17'd40411,17'd41160,17'd5354,17'd18142,17'd5026,17'd38201,17'd5027,17'd12636,17'd13420,17'd16492,17'd6094,17'd7705,17'd35487,17'd64917,17'd65564,17'd65564,17'd64917,17'd65439,17'd65180,17'd65440,17'd65700,17'd16855,17'd43596,17'd44019,17'd38860,17'd39182,17'd12635,17'd13932,17'd65565,17'd14735,17'd16381,17'd65701,17'd65702,17'd64919,17'd65054,17'd65054,17'd65054,17'd65569,17'd65569,17'd65570,17'd65703,17'd65306,17'd64241,17'd64921,17'd65055,17'd65055,17'd64653,17'd64922,17'd65704,17'd65705,17'd65706,17'd65707,17'd49810,17'd2892,17'd52099,17'd37817,17'd65708,17'd65574,17'd65709,17'd58367,17'd65575
},
'{
17'd5204,17'd4086,17'd4086,17'd13943,17'd13943,17'd4086,17'd3592,17'd15496,17'd15496,17'd3751,17'd65576,17'd65710,17'd65711,17'd64795,17'd65712,17'd65713,17'd65714,17'd65715,17'd65716,17'd65717,17'd65718,17'd8344,17'd10921,17'd9270,17'd64668,17'd9815,17'd2596,17'd9969,17'd1414,17'd17,17'd11,17'd20404,17'd17,17'd1414,17'd2597,17'd3429,17'd10669,17'd10802,17'd3251,17'd3251,17'd3101,17'd3251,17'd3428,17'd15358,17'd15877,17'd5511,17'd5203,17'd5203,17'd4425,17'd27713,17'd3427,17'd10802,17'd656,17'd471,17'd986,17'd15497,17'd59497,17'd477,17'd57000,17'd302,17'd14991,17'd63,17'd18391,17'd488,17'd2440,17'd16145,17'd484,17'd2789,17'd65719,17'd13306,17'd61950,17'd32732,17'd65720,17'd39038,17'd1288,17'd63673,17'd63525,17'd65721,17'd64803,17'd65722,17'd65723,17'd65724,17'd65592,17'd65725,17'd46032,17'd65726,17'd8380,17'd8378,17'd7916,17'd64273,17'd65727,17'd8380,17'd65728,17'd7261,17'd6937,17'd62874,17'd65729,17'd53236,17'd6150,17'd63136,17'd5249,17'd65730,17'd65598,17'd65599,17'd65731,17'd58641,17'd58761,17'd65732,17'd57910,17'd53370,17'd58519,17'd53810,17'd65600,17'd53951,17'd65733,17'd65734,17'd65735,17'd56021,17'd55900,17'd56446,17'd58272,17'd65736,17'd65737,17'd65738,17'd54346,17'd54888,17'd56574,17'd64144,17'd65739,17'd63545,17'd64556,17'd65740,17'd57396,17'd59517,17'd61441,17'd61441,17'd64148,17'd58660,17'd57784,17'd59281,17'd62232,17'd63146,17'd56810,17'd64004,17'd58154,17'd59016,17'd62473,17'd65741,17'd65742,17'd65743,17'd65744,17'd9849,17'd65483,17'd65745,17'd65746,17'd65747,17'd65748,17'd65749,17'd65750,17'd64701,17'd65100,17'd65346,17'd65751,17'd65752,17'd65753,17'd65754,17'd63433,17'd63721,17'd63306,17'd65755,17'd64844,17'd65756,17'd64170,17'd64170,17'd65349,17'd63871,17'd64028,17'd63438,17'd59688,17'd65757,17'd65758,17'd65759,17'd15172,17'd10974,17'd65760,17'd28938,17'd11805,17'd12262,17'd13646,17'd49748,17'd17480,17'd32124,17'd65761,17'd50215,17'd8573,17'd8733,17'd65762,17'd19647,17'd63738,17'd12431,17'd23348,17'd63450,17'd63450,17'd64847,17'd63736,17'd23527,17'd55833,17'd65501,17'd7801,17'd7967,17'd65763,17'd65764,17'd65632,17'd65765,17'd65766,17'd65767,17'd17978,17'd65768,17'd65769,17'd17023,17'd65770,17'd17024,17'd10037,17'd13776,17'd8132,17'd133,17'd542,17'd542,17'd1044,17'd3167,17'd5463,17'd3167,17'd5309,17'd11289,17'd13901,17'd20623,17'd65771,17'd65772,17'd65773,17'd51888,17'd65774,17'd65775,17'd65776,17'd65777,17'd65778,17'd65779,17'd64724,17'd65780,17'd65781,17'd65782,17'd65783,17'd59852,17'd65514,17'd64877,17'd64603,17'd65784,17'd65649,17'd64061,17'd65261,17'd24420,17'd65785,17'd65518,17'd52074,17'd52074,17'd65378,17'd59083,17'd59206,17'd59205,17'd59206,17'd59206,17'd58951,17'd58951,17'd59083,17'd59083,17'd59083,17'd65378,17'd65378,17'd65378,17'd58707,17'd58707,17'd58707,17'd58707,17'd60480,17'd58822,17'd53192,17'd58949,17'd56751,17'd58821,17'd65786,17'd65787,17'd65520,17'd65788,17'd65654,17'd65655,17'd65523,17'd65789,17'd64728,17'd65790,17'd65791,17'd65792,17'd58952,17'd61500,17'd51233,17'd51233,17'd57708,17'd57708,17'd65793,17'd65794,17'd65794,17'd49786,17'd65526,17'd65660,17'd35876,17'd65795,17'd60723,17'd65796,17'd36561,17'd65797,17'd63769,17'd64613,17'd65798,17'd63349,17'd65275,17'd65667,17'd65799,17'd65800,17'd21103,17'd65801,17'd65802,17'd65803,17'd65279,17'd19671,17'd65804,17'd19949,17'd65805,17'd65806,17'd20796,17'd17399,17'd24469,17'd47847,17'd23617,17'd65807,17'd65808,17'd24141,17'd53138,17'd11830,17'd10359,17'd10197,17'd7165,17'd7009,17'd6842,17'd6841,17'd24480,17'd24480,17'd6547,17'd6547,17'd5478,17'd5478,17'd5002,17'd25627,17'd5165,17'd5170,17'd8630,17'd8156,17'd7331,17'd11433,17'd65809,17'd65810,17'd65811,17'd65812,17'd65813,17'd65417,17'd65814,17'd65037,17'd65815,17'd64507,17'd63941,17'd65042,17'd15101,17'd64509,17'd63357,17'd64769,17'd65687,17'd65421,17'd63640,17'd63640,17'd63639,17'd65555,17'd65555,17'd65041,17'd65685,17'd65687,17'd65421,17'd65040,17'd65816,17'd15231,17'd18031,17'd65817,17'd65818,17'd65819,17'd65820,17'd6571,17'd65821,17'd48732,17'd65822,17'd65823,17'd3208,17'd3054,17'd65824,17'd65825,17'd50383,17'd2725,17'd46238,17'd65826,17'd65827,17'd8786,17'd3563,17'd6081,17'd48558,17'd40100,17'd39180,17'd4554,17'd18142,17'd4711,17'd5027,17'd11868,17'd12773,17'd12914,17'd5789,17'd8187,17'd11882,17'd36903,17'd65179,17'd65828,17'd64917,17'd65179,17'd65439,17'd59125,17'd58865,17'd44850,17'd16855,17'd13176,17'd41481,17'd38334,17'd44966,17'd13571,17'd65565,17'd65565,17'd62575,17'd65829,17'd65830,17'd65702,17'd64919,17'd65054,17'd65054,17'd65568,17'd65568,17'd65569,17'd65570,17'd65703,17'd64241,17'd65307,17'd65055,17'd65831,17'd65055,17'd63809,17'd65832,17'd64389,17'd14734,17'd65833,17'd62205,17'd49810,17'd65834,17'd65835,17'd41620,17'd65708,17'd65836,17'd65837,17'd58367,17'd61278
},
'{
17'd4086,17'd4086,17'd13943,17'd13943,17'd13943,17'd3901,17'd3901,17'd3901,17'd15496,17'd3751,17'd4088,17'd65576,17'd65838,17'd63976,17'd65839,17'd65840,17'd65841,17'd65716,17'd65842,17'd65843,17'd65844,17'd65845,17'd7886,17'd6591,17'd9967,17'd12929,17'd9815,17'd65450,17'd2936,17'd16,17'd10,17'd1128,17'd3905,17'd1416,17'd2257,17'd2258,17'd52621,17'd10802,17'd3251,17'd34512,17'd2935,17'd3101,17'd3428,17'd15358,17'd15877,17'd15359,17'd14744,17'd14744,17'd5646,17'd4891,17'd3428,17'd2934,17'd11071,17'd471,17'd473,17'd15362,17'd59497,17'd65451,17'd58505,17'd817,17'd21329,17'd22616,17'd2790,17'd1980,17'd41162,17'd16145,17'd14451,17'd2789,17'd65846,17'd38722,17'd38866,17'd32090,17'd2950,17'd998,17'd1428,17'd62212,17'd65847,17'd65848,17'd65849,17'd65456,17'd65850,17'd65851,17'd65852,17'd65853,17'd16291,17'd65854,17'd65855,17'd8382,17'd7916,17'd64273,17'd65856,17'd65727,17'd25659,17'd7757,17'd7421,17'd6632,17'd65857,17'd53236,17'd6149,17'd61301,17'd4921,17'd5248,17'd14894,17'd65599,17'd65599,17'd65858,17'd58392,17'd57769,17'd58027,17'd53163,17'd58519,17'd53810,17'd53685,17'd65467,17'd57505,17'd56344,17'd54431,17'd65602,17'd55900,17'd58649,17'd54700,17'd65736,17'd65736,17'd65859,17'd58649,17'd65602,17'd54701,17'd59516,17'd57641,17'd63545,17'd58652,17'd61702,17'd56458,17'd58160,17'd59517,17'd57512,17'd59018,17'd57022,17'd58887,17'd59524,17'd58771,17'd62232,17'd56810,17'd62726,17'd65860,17'd58885,17'd57915,17'd57021,17'd56809,17'd3959,17'd65861,17'd9582,17'd65862,17'd65863,17'd65864,17'd65747,17'd65865,17'd65866,17'd64838,17'd65221,17'd65220,17'd65346,17'd65867,17'd65868,17'd65490,17'd64701,17'd63569,17'd65103,17'd65347,17'd63033,17'd63034,17'd64964,17'd65349,17'd64170,17'd65869,17'd64170,17'd64028,17'd64968,17'd62139,17'd58922,17'd65870,17'd65871,17'd12236,17'd11257,17'd30368,17'd32590,17'd16198,17'd15186,17'd11807,17'd49748,17'd56952,17'd65872,17'd65873,17'd51701,17'd9047,17'd8733,17'd65874,17'd22652,17'd17132,17'd65875,17'd12869,17'd13895,17'd15064,17'd65876,17'd65877,17'd20758,17'd63742,17'd16082,17'd65878,17'd9627,17'd11818,17'd12597,17'd23010,17'd13898,17'd65879,17'd65880,17'd13380,17'd13897,17'd65881,17'd11003,17'd14944,17'd11007,17'd7812,17'd11289,17'd3025,17'd1197,17'd133,17'd542,17'd6198,17'd5309,17'd3167,17'd1044,17'd23194,17'd6198,17'd13777,17'd20622,17'd21680,17'd52655,17'd65882,17'd65883,17'd65884,17'd65885,17'd65886,17'd65887,17'd65888,17'd65889,17'd65890,17'd65891,17'd65892,17'd65893,17'd65894,17'd65895,17'd65896,17'd65264,17'd64474,17'd64475,17'd64475,17'd65375,17'd64203,17'd65785,17'd65897,17'd65651,17'd51473,17'd52815,17'd52074,17'd51473,17'd58707,17'd58707,17'd58707,17'd58707,17'd58824,17'd59454,17'd65378,17'd65378,17'd59083,17'd65378,17'd65378,17'd58707,17'd51473,17'd51473,17'd52074,17'd52074,17'd53192,17'd53192,17'd53192,17'd58949,17'd56751,17'd58950,17'd65787,17'd65898,17'd65521,17'd65522,17'd65655,17'd65656,17'd59078,17'd64728,17'd65899,17'd63464,17'd63330,17'd65900,17'd58210,17'd64193,17'd61500,17'd63897,17'd61500,17'd63897,17'd57325,17'd50561,17'd61630,17'd64743,17'd65392,17'd65901,17'd63208,17'd65902,17'd65903,17'd65904,17'd65905,17'd65906,17'd20945,17'd65907,17'd65908,17'd65909,17'd65667,17'd65910,17'd65911,17'd64359,17'd65912,17'd65913,17'd65914,17'd65915,17'd65279,17'd64891,17'd65912,17'd65916,17'd65917,17'd17994,17'd65918,17'd18012,17'd65919,17'd65920,17'd22753,17'd65807,17'd65921,17'd24141,17'd25221,17'd65922,17'd10359,17'd52521,17'd7009,17'd7009,17'd6842,17'd6841,17'd6211,17'd6547,17'd6547,17'd5149,17'd5478,17'd4844,17'd25627,17'd25627,17'd5165,17'd51930,17'd6394,17'd6561,17'd7503,17'd65923,17'd65924,17'd65925,17'd65926,17'd65681,17'd65927,17'd65928,17'd65929,17'd65930,17'd64506,17'd64507,17'd65931,17'd15230,17'd64509,17'd64509,17'd64769,17'd65555,17'd65687,17'd65421,17'd64090,17'd63640,17'd63639,17'd63639,17'd63639,17'd65165,17'd65687,17'd65421,17'd64369,17'd65040,17'd65932,17'd15231,17'd18031,17'd65933,17'd65818,17'd65934,17'd10070,17'd65935,17'd65936,17'd9788,17'd65937,17'd65938,17'd48809,17'd65939,17'd2886,17'd65940,17'd41904,17'd2888,17'd4222,17'd45785,17'd62072,17'd45067,17'd65941,17'd5493,17'd43742,17'd39789,17'd65942,17'd18383,17'd18142,17'd38458,17'd11868,17'd12636,17'd12773,17'd14060,17'd6094,17'd7537,17'd35487,17'd36905,17'd65179,17'd65828,17'd64917,17'd65943,17'd65439,17'd65944,17'd65945,17'd15104,17'd14177,17'd12913,17'd38580,17'd39182,17'd65946,17'd65947,17'd65947,17'd65948,17'd62575,17'd65949,17'd65950,17'd63963,17'd65054,17'd65054,17'd65568,17'd65568,17'd65568,17'd65305,17'd65570,17'd63965,17'd64241,17'd64921,17'd65831,17'd65831,17'd65055,17'd63809,17'd65832,17'd65951,17'd62854,17'd62332,17'd65952,17'd3559,17'd2891,17'd65835,17'd2369,17'd39787,17'd65953,17'd65837,17'd58367,17'd62196
},
'{
17'd15496,17'd3901,17'd4738,17'd13943,17'd3901,17'd3427,17'd3428,17'd15358,17'd3592,17'd3901,17'd4088,17'd3904,17'd65577,17'd64795,17'd65954,17'd65955,17'd65956,17'd65957,17'd65958,17'd65843,17'd65959,17'd65960,17'd9807,17'd7220,17'd63820,17'd12652,17'd63260,17'd14742,17'd65961,17'd1415,17'd18,17'd20404,17'd1128,17'd3905,17'd2257,17'd2258,17'd2422,17'd2935,17'd3101,17'd34512,17'd3101,17'd3101,17'd3251,17'd15358,17'd15877,17'd15359,17'd14744,17'd15117,17'd14744,17'd5203,17'd4086,17'd3901,17'd10924,17'd12196,17'd12504,17'd14989,17'd65962,17'd59497,17'd477,17'd818,17'd53,17'd65963,17'd481,17'd14603,17'd2439,17'd670,17'd2613,17'd1428,17'd3917,17'd65964,17'd34167,17'd1708,17'd2611,17'd2949,17'd1561,17'd65965,17'd64262,17'd65966,17'd65967,17'd65968,17'd65969,17'd65970,17'd65971,17'd65972,17'd65973,17'd32266,17'd65974,17'd9161,17'd8219,17'd7755,17'd9985,17'd65975,17'd65976,17'd6304,17'd7100,17'd39647,17'd40581,17'd65857,17'd65977,17'd5839,17'd62873,17'd65978,17'd65979,17'd58267,17'd65980,17'd13842,17'd58269,17'd47974,17'd52710,17'd56572,17'd57382,17'd57382,17'd53950,17'd53950,17'd65981,17'd65733,17'd65982,17'd65983,17'd56126,17'd58150,17'd58521,17'd58399,17'd65736,17'd65984,17'd58521,17'd58649,17'd54346,17'd65202,17'd56448,17'd65985,17'd57395,17'd55182,17'd58405,17'd65986,17'd58654,17'd58893,17'd57779,17'd58654,17'd57918,17'd59274,17'd62475,17'd60176,17'd58042,17'd59280,17'd64004,17'd57915,17'd64004,17'd58406,17'd65987,17'd65988,17'd64134,17'd65989,17'd65990,17'd65991,17'd65746,17'd65486,17'd65992,17'd65866,17'd65489,17'd65219,17'd65993,17'd65994,17'd65868,17'd65867,17'd65867,17'd65100,17'd63867,17'd63432,17'd65995,17'd65996,17'd65997,17'd64573,17'd65349,17'd65869,17'd65998,17'd65999,17'd64028,17'd64968,17'd63175,17'd60962,17'd60344,17'd66000,17'd12235,17'd66001,17'd66002,17'd66003,17'd28827,17'd43219,17'd13138,17'd66004,17'd16314,17'd66005,17'd66006,17'd23866,17'd57186,17'd19923,17'd17482,17'd66007,17'd66008,17'd54650,17'd24050,17'd17243,17'd16572,17'd63736,17'd23691,17'd66009,17'd11408,17'd16214,17'd66010,17'd66011,17'd62269,17'd10348,17'd11681,17'd63047,17'd25010,17'd11148,17'd53713,17'd53713,17'd53904,17'd66012,17'd22488,17'd10351,17'd66013,17'd542,17'd1481,17'd133,17'd133,17'd1045,17'd11413,17'd8132,17'd6198,17'd6198,17'd356,17'd16220,17'd3025,17'd16090,17'd23536,17'd24056,17'd21068,17'd66014,17'd66015,17'd66016,17'd66017,17'd66018,17'd66019,17'd66020,17'd65369,17'd66021,17'd66022,17'd66023,17'd66024,17'd66024,17'd66025,17'd58816,17'd66026,17'd64877,17'd65259,17'd66027,17'd65374,17'd66028,17'd62536,17'd66029,17'd24254,17'd66030,17'd65786,17'd65786,17'd65652,17'd65519,17'd66031,17'd66031,17'd65519,17'd65519,17'd65382,17'd65382,17'd65263,17'd65263,17'd66028,17'd65381,17'd65518,17'd65518,17'd65651,17'd65651,17'd65652,17'd65652,17'd65652,17'd66032,17'd65787,17'd65520,17'd65788,17'd65521,17'd65522,17'd66033,17'd65384,17'd65137,17'd65524,17'd63604,17'd63896,17'd63896,17'd63756,17'd66034,17'd61900,17'd66035,17'd66035,17'd61901,17'd66036,17'd63897,17'd66037,17'd66038,17'd66039,17'd53051,17'd66040,17'd66041,17'd23553,17'd44229,17'd35574,17'd36711,17'd66042,17'd66043,17'd19944,17'd65275,17'd66044,17'd66045,17'd66046,17'd66047,17'd66048,17'd21102,17'd66049,17'd66050,17'd66051,17'd66052,17'd66053,17'd22364,17'd20483,17'd65157,17'd66054,17'd66055,17'd17158,17'd19709,17'd66056,17'd47957,17'd22583,17'd53576,17'd22585,17'd25877,17'd11830,17'd26584,17'd10627,17'd52521,17'd7009,17'd7009,17'd6548,17'd5149,17'd6548,17'd5149,17'd5149,17'd52352,17'd4844,17'd5611,17'd5612,17'd5160,17'd37030,17'd5338,17'd6394,17'd7839,17'd65678,17'd66057,17'd66058,17'd66059,17'd65681,17'd66060,17'd66061,17'd65162,17'd65930,17'd66062,17'd66063,17'd66064,17'd65555,17'd64769,17'd64768,17'd63495,17'd63640,17'd64090,17'd64090,17'd64090,17'd63640,17'd63640,17'd63640,17'd63640,17'd65687,17'd65687,17'd63789,17'd63789,17'd63789,17'd15998,17'd14857,17'd18139,17'd65933,17'd66065,17'd66066,17'd65819,17'd66067,17'd66067,17'd66068,17'd65936,17'd66069,17'd66069,17'd8638,17'd4550,17'd4550,17'd47085,17'd46594,17'd4222,17'd45785,17'd8480,17'd48186,17'd5351,17'd10071,17'd41002,17'd39789,17'd10388,17'd18383,17'd10906,17'd5026,17'd38458,17'd11868,17'd12636,17'd14060,17'd6258,17'd6418,17'd7538,17'd35487,17'd60030,17'd64917,17'd64917,17'd65439,17'd65439,17'd65944,17'd66070,17'd65700,17'd15104,17'd13572,17'd12635,17'd44966,17'd66071,17'd13932,17'd65565,17'd65947,17'd15232,17'd62698,17'd65950,17'd65567,17'd64919,17'd66072,17'd66072,17'd65054,17'd65054,17'd66073,17'd63964,17'd63965,17'd64528,17'd63809,17'd66074,17'd66075,17'd66076,17'd66077,17'd63809,17'd63965,17'd66078,17'd13687,17'd66079,17'd48639,17'd3209,17'd2892,17'd46592,17'd46475,17'd2538,17'd66080,17'd66081,17'd1928,17'd58502
},
'{
17'd15496,17'd3592,17'd13943,17'd13943,17'd3901,17'd3427,17'd3427,17'd3428,17'd3592,17'd3901,17'd4245,17'd3904,17'd66082,17'd65312,17'd66083,17'd66084,17'd66085,17'd66086,17'd66087,17'd65957,17'd66088,17'd66089,17'd66089,17'd9130,17'd13576,17'd66090,17'd64668,17'd63259,17'd10266,17'd14442,17'd19,17'd11,17'd11,17'd3905,17'd1416,17'd2597,17'd2422,17'd2784,17'd3101,17'd3251,17'd3101,17'd3101,17'd3251,17'd15358,17'd15877,17'd15359,17'd14744,17'd66091,17'd7049,17'd15117,17'd6730,17'd4086,17'd12505,17'd11071,17'd12505,17'd58016,17'd14321,17'd15361,17'd65451,17'd44,17'd66092,17'd66093,17'd666,17'd303,17'd995,17'd669,17'd833,17'd1427,17'd33850,17'd33053,17'd3915,17'd3598,17'd66094,17'd38462,17'd2610,17'd13306,17'd61950,17'd66095,17'd66096,17'd66097,17'd66098,17'd66099,17'd66100,17'd66101,17'd66102,17'd66103,17'd30659,17'd42349,17'd8075,17'd8377,17'd8846,17'd66104,17'd65854,17'd66105,17'd65728,17'd66106,17'd47279,17'd6323,17'd6311,17'd7419,17'd62999,17'd63134,17'd4125,17'd63841,17'd65980,17'd14769,17'd14623,17'd48474,17'd47973,17'd57012,17'd53370,17'd54350,17'd53810,17'd55576,17'd54093,17'd65468,17'd65733,17'd56344,17'd56126,17'd56344,17'd64820,17'd66107,17'd65984,17'd65736,17'd58272,17'd58521,17'd58150,17'd54346,17'd65469,17'd55380,17'd66108,17'd56579,17'd62474,17'd62726,17'd62593,17'd58654,17'd62475,17'd61190,17'd59275,17'd59275,17'd66109,17'd57391,17'd58654,17'd59024,17'd56810,17'd59393,17'd59280,17'd56458,17'd66110,17'd66111,17'd66112,17'd66113,17'd18178,17'd66114,17'd65615,17'd66115,17'd64567,17'd65866,17'd65096,17'd66116,17'd65993,17'd65994,17'd65868,17'd65868,17'd65867,17'd65490,17'd65750,17'd66117,17'd66118,17'd62759,17'd65348,17'd64573,17'd64964,17'd65869,17'd65998,17'd65999,17'd66119,17'd63035,17'd66120,17'd63439,17'd58925,17'd64173,17'd12086,17'd53242,17'd51877,17'd38240,17'd10324,17'd29332,17'd13001,17'd15427,17'd17838,17'd24997,17'd66006,17'd17352,17'd24710,17'd21208,17'd18203,17'd53476,17'd66121,17'd64310,17'd55030,17'd63316,17'd61617,17'd62636,17'd66009,17'd8268,17'd11000,17'd12871,17'd64854,17'd66122,17'd10348,17'd23880,17'd23696,17'd11682,17'd17736,17'd13775,17'd15820,17'd66123,17'd63886,17'd15958,17'd14692,17'd8131,17'd718,17'd1480,17'd1481,17'd133,17'd133,17'd133,17'd15823,17'd11413,17'd3025,17'd1197,17'd4163,17'd66124,17'd1197,17'd133,17'd13777,17'd24056,17'd66125,17'd66126,17'd66127,17'd66128,17'd66129,17'd66130,17'd66131,17'd66132,17'd66133,17'd66134,17'd59447,17'd66135,17'd66023,17'd66136,17'd66025,17'd66137,17'd66138,17'd65264,17'd66139,17'd64601,17'd66140,17'd64877,17'd65381,17'd62535,17'd66141,17'd62536,17'd66142,17'd66142,17'd66142,17'd66142,17'd66030,17'd66030,17'd66030,17'd66030,17'd66032,17'd66032,17'd65652,17'd65652,17'd65786,17'd65786,17'd66143,17'd66143,17'd65651,17'd66143,17'd24254,17'd66030,17'd65787,17'd65653,17'd66144,17'd65521,17'd66145,17'd65655,17'd66146,17'd66147,17'd65137,17'd65524,17'd64999,17'd66148,17'd66149,17'd63756,17'd64189,17'd63753,17'd61900,17'd61900,17'd66034,17'd63607,17'd66036,17'd50734,17'd66150,17'd66151,17'd27373,17'd66152,17'd38993,17'd59459,17'd23554,17'd38282,17'd66153,17'd66154,17'd66155,17'd66156,17'd66157,17'd66158,17'd66159,17'd66160,17'd66161,17'd63224,17'd66162,17'd64895,17'd66163,17'd66164,17'd66165,17'd66052,17'd20076,17'd66166,17'd20950,17'd66167,17'd66168,17'd66169,17'd25217,17'd20687,17'd66170,17'd66171,17'd52992,17'd24301,17'd24942,17'd25081,17'd26584,17'd10359,17'd52521,17'd29292,17'd7166,17'd7166,17'd6549,17'd6548,17'd52352,17'd52352,17'd27569,17'd52352,17'd4844,17'd5611,17'd5158,17'd5160,17'd37030,17'd35760,17'd7670,17'd66172,17'd66173,17'd66174,17'd66175,17'd66176,17'd66177,17'd66178,17'd66179,17'd65551,17'd64902,17'd64766,17'd66064,17'd66180,17'd64769,17'd64769,17'd63495,17'd65420,17'd63789,17'd65553,17'd64090,17'd64090,17'd64090,17'd63640,17'd63640,17'd63640,17'd65421,17'd65421,17'd63789,17'd63789,17'd15998,17'd66181,17'd66182,17'd66183,17'd66184,17'd66185,17'd66186,17'd65819,17'd66187,17'd66187,17'd11186,17'd10070,17'd9788,17'd66069,17'd66188,17'd65938,17'd66189,17'd66190,17'd3865,17'd48639,17'd66191,17'd5772,17'd7680,17'd45656,17'd46596,17'd18629,17'd10790,17'd10790,17'd18383,17'd10906,17'd38458,17'd44742,17'd12483,17'd13420,17'd16492,17'd6418,17'd7538,17'd9124,17'd36905,17'd60030,17'd65179,17'd66192,17'd65439,17'd66193,17'd66194,17'd65945,17'd15104,17'd66195,17'd13689,17'd12635,17'd62331,17'd66071,17'd13932,17'd65565,17'd15103,17'd15999,17'd66196,17'd66197,17'd64919,17'd64919,17'd66072,17'd66072,17'd65054,17'd66072,17'd66073,17'd63964,17'd63658,17'd63657,17'd66198,17'd66074,17'd66199,17'd66076,17'd65831,17'd63809,17'd64109,17'd62973,17'd66200,17'd66201,17'd46594,17'd42194,17'd65834,17'd46475,17'd66202,17'd38713,17'd55880,17'd66081,17'd2069,17'd58376
},
'{
17'd15496,17'd3592,17'd13943,17'd3901,17'd3427,17'd3427,17'd3101,17'd3427,17'd3592,17'd3901,17'd4733,17'd4733,17'd66203,17'd64928,17'd65954,17'd66204,17'd66205,17'd66206,17'd66086,17'd66206,17'd66207,17'd66208,17'd66209,17'd66210,17'd7547,17'd66211,17'd9814,17'd63387,17'd66212,17'd65450,17'd18,17'd11,17'd11,17'd18,17'd1416,17'd1414,17'd2597,17'd3429,17'd2935,17'd3101,17'd14070,17'd14070,17'd3251,17'd3428,17'd15877,17'd15359,17'd7049,17'd66213,17'd66213,17'd14744,17'd5203,17'd15496,17'd10925,17'd11071,17'd12505,17'd12504,17'd14989,17'd14321,17'd59911,17'd477,17'd817,17'd664,17'd666,17'd482,17'd2438,17'd994,17'd1287,17'd1708,17'd33054,17'd53013,17'd66214,17'd4093,17'd66215,17'd13952,17'd4094,17'd1842,17'd66216,17'd66217,17'd64541,17'd66218,17'd66219,17'd65723,17'd66220,17'd66221,17'd66222,17'd18779,17'd21042,17'd9845,17'd66223,17'd8378,17'd25659,17'd9842,17'd66224,17'd65727,17'd8220,17'd39812,17'd46999,17'd45528,17'd42350,17'd7419,17'd6630,17'd60783,17'd4125,17'd4769,17'd63996,17'd14769,17'd13842,17'd14099,17'd56340,17'd58030,17'd53370,17'd58519,17'd58519,17'd55668,17'd54171,17'd65468,17'd66225,17'd64552,17'd56344,17'd66226,17'd58031,17'd58272,17'd57013,17'd48931,17'd48931,17'd56803,17'd58272,17'd66227,17'd65982,17'd64824,17'd56241,17'd56912,17'd64146,17'd59517,17'd57396,17'd62726,17'd58154,17'd66228,17'd57512,17'd59275,17'd56697,17'd65335,17'd60177,17'd56453,17'd63146,17'd57512,17'd59280,17'd65607,17'd61188,17'd66229,17'd5082,17'd66230,17'd14638,17'd66231,17'd66232,17'd66115,17'd64699,17'd66233,17'd65096,17'd65616,17'd65346,17'd65994,17'd65868,17'd66234,17'd66235,17'd66236,17'd64839,17'd66237,17'd66238,17'd61468,17'd62904,17'd63724,17'd64964,17'd65349,17'd65999,17'd64170,17'd66239,17'd63173,17'd66120,17'd64444,17'd66240,17'd66241,17'd16433,17'd26490,17'd66242,17'd66243,17'd10161,17'd10472,17'd13001,17'd10605,17'd26497,17'd18556,17'd66244,17'd33716,17'd8732,17'd19923,17'd8420,17'd66245,17'd54048,17'd20615,17'd18690,17'd66246,17'd13530,17'd8267,17'd16082,17'd66247,17'd13531,17'd14820,17'd23879,17'd66248,17'd11974,17'd63047,17'd66249,17'd9898,17'd10350,17'd66012,17'd66012,17'd64855,17'd16577,17'd66250,17'd16811,17'd717,17'd542,17'd1481,17'd1481,17'd1481,17'd133,17'd133,17'd1045,17'd1045,17'd1197,17'd1197,17'd66124,17'd356,17'd133,17'd133,17'd15823,17'd24056,17'd66251,17'd52732,17'd66252,17'd66253,17'd66254,17'd66255,17'd66256,17'd66257,17'd66258,17'd66259,17'd66260,17'd66261,17'd66022,17'd66135,17'd66135,17'd66023,17'd66262,17'd65896,17'd66263,17'd65140,17'd66139,17'd64878,17'd65265,17'd65787,17'd66264,17'd66265,17'd66266,17'd66266,17'd66266,17'd66266,17'd66267,17'd66267,17'd66267,17'd66268,17'd66142,17'd66142,17'd66030,17'd66142,17'd66142,17'd66142,17'd66142,17'd66030,17'd66030,17'd24254,17'd66268,17'd66032,17'd66269,17'd65654,17'd65522,17'd65383,17'd65254,17'd66270,17'd65523,17'd66271,17'd59448,17'd65790,17'd63464,17'd63463,17'd66272,17'd66273,17'd66273,17'd66274,17'd66275,17'd63605,17'd61900,17'd58210,17'd66276,17'd66277,17'd50155,17'd51650,17'd26904,17'd66152,17'd32031,17'd59458,17'd42749,17'd66278,17'd66279,17'd62030,17'd66280,17'd66281,17'd66282,17'd66283,17'd66284,17'd66285,17'd66286,17'd66287,17'd66288,17'd66289,17'd66290,17'd66291,17'd66292,17'd66293,17'd20483,17'd22194,17'd66294,17'd66295,17'd66055,17'd66296,17'd66297,17'd20687,17'd66298,17'd52903,17'd24299,17'd66299,17'd25360,17'd25221,17'd26826,17'd10627,17'd29292,17'd8913,17'd7328,17'd7166,17'd6549,17'd6549,17'd4843,17'd4843,17'd4843,17'd4843,17'd5002,17'd5329,17'd5160,17'd5160,17'd51930,17'd8473,17'd7839,17'd66300,17'd66057,17'd66301,17'd66302,17'd66303,17'd66304,17'd66305,17'd65162,17'd65037,17'd65419,17'd64766,17'd65289,17'd64227,17'd64769,17'd64769,17'd63495,17'd63640,17'd63789,17'd66306,17'd65553,17'd65553,17'd65553,17'd65553,17'd65421,17'd65421,17'd65688,17'd65688,17'd65040,17'd65040,17'd66307,17'd16491,17'd65557,17'd66183,17'd66308,17'd66309,17'd66310,17'd18979,17'd66068,17'd10788,17'd10070,17'd9788,17'd66311,17'd66312,17'd8946,17'd66313,17'd3865,17'd48733,17'd48733,17'd45785,17'd66314,17'd45656,17'd45786,17'd10071,17'd46354,17'd43462,17'd45186,17'd10790,17'd18383,17'd10906,17'd11867,17'd66315,17'd12773,17'd13177,17'd6891,17'd6890,17'd7705,17'd38460,17'd36905,17'd63652,17'd65943,17'd65943,17'd65439,17'd66316,17'd66070,17'd65700,17'd15104,17'd16855,17'd13572,17'd13056,17'd66071,17'd13932,17'd65565,17'd65947,17'd15103,17'd15483,17'd66196,17'd63963,17'd66317,17'd66317,17'd66318,17'd66319,17'd65054,17'd66072,17'd66073,17'd63964,17'd63658,17'd64528,17'd64653,17'd65055,17'd66320,17'd66320,17'd65055,17'd63657,17'd66321,17'd66322,17'd64924,17'd18864,17'd4222,17'd3059,17'd38713,17'd38855,17'd2726,17'd53672,17'd62334,17'd32722,17'd1928,17'd58502
},
'{
17'd3592,17'd3901,17'd13943,17'd13943,17'd3901,17'd2934,17'd3101,17'd3101,17'd3428,17'd3427,17'd4246,17'd4733,17'd66323,17'd65187,17'd66324,17'd66325,17'd66326,17'd66327,17'd66328,17'd66327,17'd66329,17'd66330,17'd66331,17'd66332,17'd7718,17'd63977,17'd66333,17'd14441,17'd63387,17'd65961,17'd17,17'd11,17'd11,17'd1128,17'd3905,17'd1416,17'd2596,17'd3752,17'd2422,17'd3252,17'd14070,17'd14070,17'd3101,17'd3427,17'd15496,17'd15359,17'd7049,17'd14745,17'd66213,17'd66091,17'd5203,17'd5511,17'd16501,17'd10924,17'd12196,17'd12505,17'd58016,17'd14989,17'd15497,17'd815,17'd1419,17'd820,17'd666,17'd827,17'd2788,17'd2612,17'd1141,17'd1842,17'd32730,17'd51861,17'd51861,17'd5057,17'd66334,17'd66335,17'd66336,17'd4094,17'd34168,17'd66337,17'd64403,17'd66338,17'd66339,17'd66340,17'd66341,17'd66342,17'd66343,17'd66344,17'd66345,17'd43467,17'd66346,17'd8382,17'd24841,17'd24841,17'd28669,17'd65727,17'd8379,17'd7423,17'd49202,17'd51256,17'd52030,17'd6936,17'd6936,17'd62998,17'd63134,17'd60290,17'd59011,17'd58267,17'd14769,17'd14623,17'd66347,17'd47865,17'd56343,17'd58519,17'd58519,17'd55576,17'd54171,17'd54172,17'd54706,17'd66348,17'd65733,17'd55775,17'd66227,17'd48932,17'd53950,17'd48931,17'd57013,17'd56900,17'd57013,17'd48932,17'd66349,17'd66350,17'd64419,17'd55283,17'd57277,17'd55281,17'd56131,17'd58160,17'd58891,17'd59280,17'd57393,17'd61190,17'd59400,17'd59145,17'd66351,17'd65334,17'd66352,17'd62232,17'd64148,17'd58277,17'd62102,17'd60538,17'd4462,17'd66104,17'd18306,17'd66353,17'd66354,17'd66115,17'd65095,17'd65346,17'd65345,17'd66355,17'd65994,17'd66356,17'd66234,17'd66357,17'd66234,17'd65751,17'd64959,17'd64164,17'd62622,17'd61602,17'd66358,17'd66359,17'd63573,17'd65349,17'd65869,17'd64170,17'd66239,17'd63872,17'd61741,17'd66360,17'd66361,17'd66362,17'd13632,17'd66363,17'd66364,17'd51196,17'd33253,17'd41194,17'd31130,17'd10476,17'd26497,17'd15681,17'd12725,17'd10340,17'd8887,17'd37734,17'd8420,17'd55523,17'd21366,17'd7626,17'd59565,17'd63450,17'd64312,17'd66365,17'd15954,17'd8433,17'd66366,17'd14942,17'd13532,17'd66367,17'd66368,17'd22659,17'd13260,17'd11976,17'd10036,17'd66369,17'd64315,17'd66370,17'd52731,17'd65361,17'd53638,17'd542,17'd133,17'd356,17'd1481,17'd133,17'd133,17'd133,17'd133,17'd1045,17'd1197,17'd1197,17'd66124,17'd1481,17'd133,17'd133,17'd16090,17'd24056,17'd66371,17'd21377,17'd66372,17'd66373,17'd66374,17'd66375,17'd66376,17'd66377,17'd66378,17'd66379,17'd66380,17'd65133,17'd65781,17'd66022,17'd66381,17'd66023,17'd66382,17'd65647,17'd65788,17'd65263,17'd66383,17'd65648,17'd65265,17'd65264,17'd65787,17'd66266,17'd66264,17'd66384,17'd66266,17'd66266,17'd66267,17'd66267,17'd66266,17'd66266,17'd62536,17'd62536,17'd62536,17'd62536,17'd62536,17'd62535,17'd24254,17'd24254,17'd62535,17'd66385,17'd65653,17'd65521,17'd65522,17'd65514,17'd66033,17'd65656,17'd66270,17'd65523,17'd59078,17'd66386,17'd65899,17'd66387,17'd66388,17'd66389,17'd66390,17'd66391,17'd66392,17'd66274,17'd66275,17'd63605,17'd66035,17'd65003,17'd64741,17'd66393,17'd66394,17'd28721,17'd31211,17'd31211,17'd66395,17'd26175,17'd66396,17'd66397,17'd66398,17'd66399,17'd66400,17'd66401,17'd66402,17'd66403,17'd66404,17'd66405,17'd66406,17'd66407,17'd66408,17'd66409,17'd66410,17'd66411,17'd66412,17'd65802,17'd20485,17'd20795,17'd65805,17'd66413,17'd18718,17'd66414,17'd16945,17'd66415,17'd66416,17'd66417,17'd66418,17'd24473,17'd11985,17'd11830,17'd10627,17'd52521,17'd8913,17'd7990,17'd7328,17'd7166,17'd5913,17'd6549,17'd4843,17'd4843,17'd4843,17'd4844,17'd5329,17'd5160,17'd5160,17'd37030,17'd34336,17'd8156,17'd66419,17'd66420,17'd66421,17'd66059,17'd66422,17'd66423,17'd66061,17'd66179,17'd65551,17'd65163,17'd65419,17'd64766,17'd64227,17'd64089,17'd64769,17'd64769,17'd65555,17'd63640,17'd63789,17'd65553,17'd65553,17'd65684,17'd65684,17'd65684,17'd64369,17'd65688,17'd65688,17'd65688,17'd65040,17'd65040,17'd14733,17'd66424,17'd17178,17'd18139,17'd65691,17'd66425,17'd66426,17'd66427,17'd66428,17'd66429,17'd66430,17'd66431,17'd66432,17'd66432,17'd66190,17'd48639,17'd48639,17'd45785,17'd66191,17'd66314,17'd45656,17'd10071,17'd46136,17'd46354,17'd43462,17'd43462,17'd10790,17'd10790,17'd10906,17'd39181,17'd50291,17'd62845,17'd66433,17'd13176,17'd14858,17'd7878,17'd38460,17'd64648,17'd60030,17'd63652,17'd65943,17'd65943,17'd66193,17'd65944,17'd65700,17'd15735,17'd16855,17'd14584,17'd13689,17'd13056,17'd66071,17'd13932,17'd65565,17'd66434,17'd15232,17'd15483,17'd62970,17'd66435,17'd66436,17'd66317,17'd66319,17'd66319,17'd65054,17'd66437,17'd66073,17'd64109,17'd63658,17'd63657,17'd64921,17'd65055,17'd66320,17'd66320,17'd64921,17'd63809,17'd63246,17'd62701,17'd66438,17'd9941,17'd46594,17'd46476,17'd2891,17'd42193,17'd2727,17'd41768,17'd55563,17'd61283,17'd58742,17'd58502
},
'{
17'd3901,17'd3751,17'd4738,17'd3901,17'd3427,17'd2934,17'd3101,17'd3101,17'd3427,17'd3427,17'd2935,17'd2593,17'd6264,17'd64927,17'd66439,17'd66325,17'd66326,17'd66440,17'd66441,17'd66442,17'd66443,17'd66444,17'd66445,17'd66446,17'd8817,17'd65581,17'd66447,17'd11607,17'd14441,17'd14069,17'd16,17'd10,17'd11,17'd1128,17'd3905,17'd17,17'd1414,17'd2597,17'd2258,17'd3429,17'd14070,17'd14070,17'd3101,17'd3427,17'd4892,17'd4426,17'd4734,17'd6263,17'd5959,17'd5645,17'd15359,17'd5511,17'd16011,17'd10924,17'd10924,17'd12505,17'd16392,17'd58016,17'd15362,17'd41,17'd1697,17'd1555,17'd825,17'd992,17'd45404,17'd2949,17'd1425,17'd1707,17'd4093,17'd51861,17'd32562,17'd5381,17'd51415,17'd5057,17'd66334,17'd4435,17'd31732,17'd66216,17'd66217,17'd66448,17'd66449,17'd66450,17'd66451,17'd66342,17'd66452,17'd66453,17'd66454,17'd66455,17'd9580,17'd8696,17'd8848,17'd25259,17'd24976,17'd8381,17'd8380,17'd8379,17'd7423,17'd64413,17'd6636,17'd6474,17'd6936,17'd62999,17'd66456,17'd62997,17'd4769,17'd63996,17'd9704,17'd13842,17'd14624,17'd56340,17'd57012,17'd56343,17'd55483,17'd66457,17'd54020,17'd66458,17'd63845,17'd54706,17'd66348,17'd54894,17'd55899,17'd55774,17'd55668,17'd53810,17'd56232,17'd56232,17'd55483,17'd56125,17'd53756,17'd66459,17'd66350,17'd54803,17'd55380,17'd66460,17'd66461,17'd63003,17'd62878,17'd66462,17'd60176,17'd58526,17'd59024,17'd56453,17'd66463,17'd66464,17'd63695,17'd61190,17'd57022,17'd61309,17'd65741,17'd66465,17'd66466,17'd66105,17'd41922,17'd66467,17'd64564,17'd66115,17'd66468,17'd66356,17'd65616,17'd66469,17'd66470,17'd66471,17'd66472,17'd66473,17'd66472,17'd65867,17'd65993,17'd64165,17'd65491,17'd66474,17'd66475,17'd65105,17'd65223,17'd65869,17'd65869,17'd65869,17'd65999,17'd63872,17'd65224,17'd66476,17'd61613,17'd66477,17'd13242,17'd55119,17'd66478,17'd31437,17'd10020,17'd41194,17'd17009,17'd10855,17'd15052,17'd15051,17'd10607,17'd36775,17'd25678,17'd59845,17'd33716,17'd55419,17'd61618,17'd63882,17'd66479,17'd63450,17'd66480,17'd66365,17'd66009,17'd66366,17'd22830,17'd23008,17'd14398,17'd17245,17'd13382,17'd66481,17'd22838,17'd12126,17'd22145,17'd24054,17'd14692,17'd66482,17'd20058,17'd10874,17'd7980,17'd133,17'd132,17'd128,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd1197,17'd1197,17'd4163,17'd1481,17'd1197,17'd1045,17'd16090,17'd21376,17'd66483,17'd66484,17'd65636,17'd66485,17'd66486,17'd66487,17'd23021,17'd66488,17'd66489,17'd66490,17'd66491,17'd66492,17'd66261,17'd66381,17'd66493,17'd66494,17'd66495,17'd66495,17'd66496,17'd65788,17'd65654,17'd66497,17'd65264,17'd66026,17'd65264,17'd65520,17'd66267,17'd66267,17'd66266,17'd66384,17'd66384,17'd66384,17'd66384,17'd66384,17'd66498,17'd66498,17'd66498,17'd66498,17'd62535,17'd24254,17'd66268,17'd66385,17'd66385,17'd65653,17'd65654,17'd66499,17'd65254,17'd66500,17'd60587,17'd66501,17'd65789,17'd66386,17'd65899,17'd59714,17'd61360,17'd61758,17'd66502,17'd66503,17'd66504,17'd66505,17'd66506,17'd62784,17'd63605,17'd63607,17'd50645,17'd56391,17'd63613,17'd66507,17'd34481,17'd24408,17'd59459,17'd65902,17'd66508,17'd66509,17'd66510,17'd66511,17'd66512,17'd31063,17'd66513,17'd19555,17'd64489,17'd66514,17'd66515,17'd66516,17'd66517,17'd66518,17'd66519,17'd66520,17'd66521,17'd66522,17'd66523,17'd65802,17'd66524,17'd20078,17'd66525,17'd66526,17'd19313,17'd19318,17'd16832,17'd66415,17'd66527,17'd66528,17'd24472,17'd24641,17'd22413,17'd11692,17'd10627,17'd52521,17'd8913,17'd7990,17'd7328,17'd6844,17'd5913,17'd5913,17'd4844,17'd4843,17'd5002,17'd5002,17'd25627,17'd5160,17'd5167,17'd51930,17'd8473,17'd6712,17'd66529,17'd66530,17'd66301,17'd66422,17'd66531,17'd66532,17'd66305,17'd65162,17'd64505,17'd65419,17'd66064,17'd66180,17'd64089,17'd66533,17'd64769,17'd64769,17'd65555,17'd63639,17'd64090,17'd65553,17'd65684,17'd66534,17'd66535,17'd64767,17'd64767,17'd64630,17'd64904,17'd64904,17'd66536,17'd66536,17'd66537,17'd66538,17'd17178,17'd66539,17'd66540,17'd66541,17'd66542,17'd66543,17'd66431,17'd66544,17'd66545,17'd66546,17'd49407,17'd3865,17'd48733,17'd48639,17'd48186,17'd5024,17'd45656,17'd10071,17'd10071,17'd46354,17'd46354,17'd43462,17'd10649,17'd10790,17'd10388,17'd10388,17'd39181,17'd11720,17'd50291,17'd12483,17'd66433,17'd48187,17'd6890,17'd7878,17'd38460,17'd59125,17'd65439,17'd66547,17'd65439,17'd65439,17'd65944,17'd65440,17'd65700,17'd16132,17'd16855,17'd14584,17'd62445,17'd64918,17'd13932,17'd65565,17'd66434,17'd15103,17'd15232,17'd16959,17'd63107,17'd66073,17'd66437,17'd66072,17'd66319,17'd66319,17'd65054,17'd66437,17'd65570,17'd65570,17'd63965,17'd63809,17'd65055,17'd65831,17'd66320,17'd66320,17'd64921,17'd66548,17'd63247,17'd66549,17'd66438,17'd9941,17'd64658,17'd66550,17'd66202,17'd42333,17'd2537,17'd53940,17'd54873,17'd61283,17'd58742,17'd62196
},
'{
17'd3901,17'd3751,17'd4738,17'd3901,17'd3427,17'd2934,17'd3101,17'd3101,17'd2934,17'd3427,17'd2935,17'd2935,17'd4733,17'd65063,17'd66551,17'd66552,17'd66326,17'd66553,17'd66554,17'd66555,17'd66556,17'd66557,17'd66558,17'd66559,17'd66560,17'd66561,17'd64120,17'd13433,17'd63520,17'd14867,17'd1415,17'd19,17'd11,17'd1128,17'd18,17'd3905,17'd1416,17'd2257,17'd2597,17'd2258,17'd3252,17'd3252,17'd2935,17'd2934,17'd4428,17'd4087,17'd4734,17'd6263,17'd5374,17'd5959,17'd14744,17'd15359,17'd16011,17'd10925,17'd10924,17'd10924,17'd11888,17'd16392,17'd1279,17'd15362,17'd39,17'd56111,17'd822,17'd824,17'd992,17'd17079,17'd17079,17'd1707,17'd4093,17'd4897,17'd5381,17'd5221,17'd4581,17'd5219,17'd5218,17'd4254,17'd32730,17'd33851,17'd66562,17'd66563,17'd65849,17'd64129,17'd66564,17'd66565,17'd66566,17'd66567,17'd66568,17'd66569,17'd11092,17'd9846,17'd8696,17'd8848,17'd25259,17'd9304,17'd28669,17'd65727,17'd8220,17'd8377,17'd6778,17'd6634,17'd6776,17'd6775,17'd6477,17'd61566,17'd4125,17'd59011,17'd8688,17'd14769,17'd14623,17'd47673,17'd48189,17'd57120,17'd55483,17'd57013,17'd58272,17'd55899,17'd56344,17'd55776,17'd66348,17'd66348,17'd65733,17'd58400,17'd55774,17'd53950,17'd56232,17'd56232,17'd49814,17'd48821,17'd53950,17'd54021,17'd66570,17'd65982,17'd56020,17'd57510,17'd66571,17'd66572,17'd66573,17'd62232,17'd66574,17'd57922,17'd66575,17'd62475,17'd63695,17'd66576,17'd66577,17'd57514,17'd58530,17'd59792,17'd66578,17'd64143,17'd63540,17'd63401,17'd66579,17'd33558,17'd66580,17'd66581,17'd66116,17'd66582,17'd66583,17'd66584,17'd66585,17'd66586,17'd66472,17'd66587,17'd66472,17'd66588,17'd65346,17'd66589,17'd66590,17'd65995,17'd66591,17'd66592,17'd66593,17'd66594,17'd65869,17'd65869,17'd65999,17'd66595,17'd66596,17'd66597,17'd60462,17'd58688,17'd17339,17'd54456,17'd66598,17'd66599,17'd9881,17'd40603,17'd40447,17'd10855,17'd10605,17'd66600,17'd48326,17'd66601,17'd8417,17'd24215,17'd33874,17'd16208,17'd14389,17'd10343,17'd18810,17'd66602,17'd66603,17'd66604,17'd16214,17'd56625,17'd23006,17'd66605,17'd11004,17'd66606,17'd10872,17'd22308,17'd22145,17'd18928,17'd11977,17'd13776,17'd13776,17'd11152,17'd10874,17'd15823,17'd1045,17'd132,17'd130,17'd129,17'd132,17'd133,17'd133,17'd133,17'd133,17'd133,17'd1197,17'd1197,17'd356,17'd1481,17'd3025,17'd1045,17'd16090,17'd23537,17'd66607,17'd66608,17'd66609,17'd66610,17'd66611,17'd66612,17'd53715,17'd66613,17'd66614,17'd66490,17'd66615,17'd66616,17'd66617,17'd66022,17'd66618,17'd66137,17'd66025,17'd66025,17'd66619,17'd66496,17'd65898,17'd65788,17'd65382,17'd66497,17'd65264,17'd65264,17'd66144,17'd65653,17'd66032,17'd66267,17'd66266,17'd66266,17'd66267,17'd66268,17'd24092,17'd66620,17'd66620,17'd66620,17'd66030,17'd65786,17'd65787,17'd65653,17'd65382,17'd65654,17'd66145,17'd66621,17'd66622,17'd64868,17'd60716,17'd60716,17'd61110,17'd59714,17'd66623,17'd66624,17'd61492,17'd66625,17'd66626,17'd63602,17'd66627,17'd66628,17'd66629,17'd66630,17'd58709,17'd59084,17'd56391,17'd57707,17'd33793,17'd26284,17'd66631,17'd24240,17'd59211,17'd66632,17'd66633,17'd66634,17'd66635,17'd66636,17'd66637,17'd30767,17'd66638,17'd66639,17'd66640,17'd66641,17'd66642,17'd66643,17'd66644,17'd66645,17'd66646,17'd66647,17'd66648,17'd66649,17'd66650,17'd66651,17'd20078,17'd66652,17'd66653,17'd66654,17'd18950,17'd19192,17'd25760,17'd66655,17'd66656,17'd24638,17'd22082,17'd25220,17'd11692,17'd11548,17'd52521,17'd30331,17'd7990,17'd7825,17'd6845,17'd6844,17'd5913,17'd5913,17'd4844,17'd4844,17'd5002,17'd25627,17'd5160,17'd36887,17'd5338,17'd34336,17'd8156,17'd7840,17'd66657,17'd65925,17'd66658,17'd66659,17'd66660,17'd66661,17'd66179,17'd65418,17'd64902,17'd64766,17'd66064,17'd64227,17'd66533,17'd66662,17'd64769,17'd64769,17'd65041,17'd65165,17'd65165,17'd64090,17'd66534,17'd64767,17'd66663,17'd66663,17'd64767,17'd64767,17'd64630,17'd64630,17'd66536,17'd66536,17'd65932,17'd66424,17'd14857,17'd66664,17'd18139,17'd66540,17'd66308,17'd66665,17'd66666,17'd66667,17'd66544,17'd66668,17'd66669,17'd66670,17'd8312,17'd9661,17'd66671,17'd66672,17'd66673,17'd46239,17'd10247,17'd10247,17'd66674,17'd66674,17'd45186,17'd10388,17'd10388,17'd10790,17'd11720,17'd50291,17'd12483,17'd44019,17'd13176,17'd16623,17'd44850,17'd66675,17'd65440,17'd59125,17'd65439,17'd66547,17'd65439,17'd66193,17'd65440,17'd66070,17'd15735,17'd16132,17'd62444,17'd62444,17'd62445,17'd62445,17'd13932,17'd66434,17'd15103,17'd15999,17'd16959,17'd62851,17'd63963,17'd66676,17'd66437,17'd65054,17'd66319,17'd66319,17'd66072,17'd66677,17'd65570,17'd64110,17'd63657,17'd64653,17'd65831,17'd66077,17'd66320,17'd65831,17'd64653,17'd63658,17'd66678,17'd66679,17'd11718,17'd66680,17'd49810,17'd66681,17'd66682,17'd51407,17'd2537,17'd53940,17'd54873,17'd61163,17'd66683,17'd62196
},
'{
17'd3427,17'd3751,17'd4738,17'd3901,17'd3427,17'd3101,17'd3101,17'd3101,17'd2593,17'd2934,17'd2935,17'd2935,17'd4733,17'd65446,17'd66684,17'd66685,17'd66326,17'd66553,17'd66686,17'd66686,17'd66687,17'd66688,17'd66689,17'd66690,17'd66691,17'd66692,17'd65839,17'd66693,17'd11607,17'd6274,17'd1414,17'd18,17'd11,17'd20,17'd11,17'd18,17'd17,17'd1416,17'd2257,17'd2257,17'd1831,17'd3252,17'd2935,17'd2934,17'd4428,17'd4087,17'd4735,17'd6263,17'd5509,17'd5374,17'd7049,17'd15359,17'd15877,17'd3427,17'd10924,17'd10924,17'd10924,17'd16501,17'd473,17'd660,17'd1700,17'd1699,17'd989,17'd991,17'd16967,17'd1139,17'd1285,17'd2268,17'd4093,17'd4897,17'd5381,17'd5221,17'd5382,17'd4742,17'd4742,17'd5218,17'd66694,17'd65964,17'd34347,17'd62213,17'd64672,17'd64265,17'd66695,17'd66696,17'd65971,17'd66697,17'd66698,17'd13216,17'd13729,17'd66699,17'd9443,17'd66346,17'd8695,17'd9305,17'd10114,17'd66105,17'd28669,17'd8847,17'd7755,17'd6937,17'd66700,17'd6316,17'd6478,17'd64140,17'd4463,17'd4291,17'd8688,17'd9704,17'd13842,17'd48474,17'd47864,17'd57632,17'd56232,17'd55483,17'd55576,17'd54171,17'd65470,17'd56344,17'd54705,17'd66701,17'd65733,17'd64820,17'd55774,17'd55668,17'd56125,17'd57636,17'd54886,17'd49814,17'd48931,17'd57125,17'd56125,17'd66702,17'd58150,17'd55284,17'd66703,17'd64422,17'd66704,17'd65335,17'd58893,17'd57134,17'd57784,17'd58526,17'd58893,17'd59274,17'd57274,17'd56808,17'd66705,17'd57784,17'd58891,17'd56911,17'd66706,17'd4768,17'd66707,17'd66708,17'd66709,17'd64436,17'd65616,17'd66710,17'd66711,17'd66712,17'd66713,17'd66714,17'd66715,17'd66716,17'd66717,17'd66588,17'd65346,17'd66589,17'd66590,17'd65995,17'd65222,17'd66718,17'd66719,17'd66720,17'd65869,17'd65869,17'd65998,17'd64028,17'd66721,17'd66722,17'd60461,17'd58563,17'd13236,17'd26140,17'd53027,17'd66723,17'd66724,17'd9737,17'd10162,17'd27002,17'd13886,17'd66600,17'd66725,17'd52952,17'd8249,17'd16072,17'd34036,17'd55616,17'd61353,17'd54829,17'd19160,17'd63586,17'd66726,17'd66009,17'd12732,17'd14942,17'd21217,17'd14539,17'd13145,17'd22488,17'd23014,17'd15702,17'd9359,17'd8444,17'd8444,17'd14016,17'd11152,17'd7980,17'd17363,17'd1045,17'd1045,17'd132,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd134,17'd1759,17'd128,17'd130,17'd1197,17'd133,17'd16090,17'd23537,17'd66727,17'd66125,17'd66728,17'd66729,17'd66730,17'd66731,17'd54297,17'd66732,17'd66733,17'd66734,17'd66735,17'd66736,17'd65251,17'd66737,17'd66738,17'd66493,17'd66739,17'd66740,17'd66741,17'd66742,17'd66742,17'd66743,17'd65788,17'd65788,17'd65521,17'd65654,17'd65264,17'd66497,17'd66144,17'd65653,17'd65787,17'd66032,17'd65787,17'd65787,17'd66744,17'd66745,17'd66745,17'd66746,17'd66032,17'd65787,17'd66269,17'd65788,17'd65514,17'd65254,17'd66622,17'd66747,17'd64868,17'd66748,17'd66749,17'd66749,17'd66750,17'd66751,17'd62275,17'd66752,17'd66625,17'd66753,17'd66754,17'd66755,17'd66756,17'd66628,17'd66757,17'd63605,17'd59084,17'd56391,17'd50648,17'd34459,17'd32353,17'd24410,17'd24241,17'd24736,17'd66758,17'd36852,17'd66759,17'd66760,17'd66761,17'd66762,17'd66763,17'd66764,17'd23766,17'd65669,17'd66641,17'd66765,17'd66766,17'd66767,17'd66768,17'd66769,17'd66770,17'd66771,17'd66772,17'd66773,17'd66774,17'd19672,17'd66775,17'd66776,17'd66777,17'd66778,17'd66779,17'd66780,17'd17526,17'd21300,17'd24471,17'd21923,17'd27813,17'd11985,17'd10882,17'd10198,17'd29292,17'd9219,17'd7661,17'd6846,17'd6845,17'd28532,17'd50670,17'd50670,17'd5611,17'd4844,17'd25627,17'd25627,17'd5335,17'd37434,17'd5338,17'd8474,17'd6712,17'd66781,17'd66782,17'd66783,17'd66422,17'd66531,17'd66784,17'd66785,17'd66786,17'd65285,17'd64368,17'd66064,17'd65289,17'd64089,17'd15997,17'd66787,17'd63357,17'd64769,17'd65041,17'd65165,17'd65165,17'd64090,17'd64629,17'd66663,17'd66788,17'd66321,17'd66321,17'd66321,17'd63376,17'd65286,17'd66789,17'd66790,17'd66791,17'd66791,17'd15231,17'd14582,17'd18267,17'd18268,17'd12770,17'd66792,17'd66793,17'd66794,17'd66795,17'd66795,17'd66795,17'd5771,17'd5771,17'd66796,17'd66797,17'd66798,17'd66798,17'd66799,17'd10649,17'd11047,17'd11188,17'd11188,17'd10790,17'd10790,17'd39482,17'd39790,17'd44742,17'd66800,17'd12483,17'd44019,17'd14177,17'd14858,17'd65700,17'd66675,17'd65944,17'd66193,17'd66801,17'd66801,17'd66802,17'd65944,17'd58865,17'd65700,17'd15104,17'd16855,17'd62444,17'd62445,17'd62445,17'd62445,17'd66803,17'd15103,17'd16381,17'd65949,17'd65701,17'd66197,17'd66317,17'd66804,17'd66437,17'd65054,17'd66318,17'd66318,17'd65569,17'd66677,17'd65703,17'd64110,17'd63657,17'd64921,17'd65831,17'd66077,17'd66077,17'd65831,17'd63809,17'd63378,17'd62701,17'd66200,17'd11718,17'd66805,17'd66806,17'd66550,17'd2890,17'd51015,17'd66807,17'd66080,17'd2079,17'd32556,17'd1927,17'd61278
},
'{
17'd3428,17'd3427,17'd3751,17'd3901,17'd3427,17'd3101,17'd2935,17'd3101,17'd2782,17'd3101,17'd3252,17'd3252,17'd4246,17'd65186,17'd64395,17'd66808,17'd66328,17'd66440,17'd66809,17'd66810,17'd66687,17'd66811,17'd66812,17'd66813,17'd66814,17'd66089,17'd65840,17'd66815,17'd6594,17'd6267,17'd9969,17'd1277,17'd10,17'd11,17'd19,17'd18,17'd17,17'd1416,17'd1414,17'd2257,17'd1831,17'd1831,17'd3252,17'd2934,17'd4428,17'd4244,17'd5646,17'd5197,17'd7048,17'd5374,17'd66213,17'd66816,17'd5511,17'd3901,17'd10924,17'd10802,17'd10924,17'd11609,17'd472,17'd473,17'd37,17'd1700,17'd21949,17'd990,17'd991,17'd16967,17'd1284,17'd66094,17'd66817,17'd51861,17'd5381,17'd5221,17'd66818,17'd5382,17'd4742,17'd13069,17'd66819,17'd66820,17'd34346,17'd66821,17'd66822,17'd66823,17'd66824,17'd66825,17'd66826,17'd66827,17'd66828,17'd13097,17'd13853,17'd11482,17'd9580,17'd66829,17'd24523,17'd9306,17'd10946,17'd10946,17'd29181,17'd28669,17'd8073,17'd7098,17'd51584,17'd42060,17'd6776,17'd6476,17'd6934,17'd4126,17'd4464,17'd9704,17'd13842,17'd14624,17'd47864,17'd48079,17'd56343,17'd48819,17'd55668,17'd66107,17'd64820,17'd56126,17'd66830,17'd65082,17'd57268,17'd54894,17'd64820,17'd58031,17'd48820,17'd57636,17'd54797,17'd48641,17'd56900,17'd57013,17'd57636,17'd56125,17'd54430,17'd66831,17'd66832,17'd66833,17'd56907,17'd62229,17'd58037,17'd60427,17'd66834,17'd59144,17'd58036,17'd57022,17'd59145,17'd58038,17'd66835,17'd65478,17'd57134,17'd55906,17'd66836,17'd5082,17'd66837,17'd66708,17'd66709,17'd66838,17'd65616,17'd66710,17'd66839,17'd66840,17'd66841,17'd66714,17'd66715,17'd66716,17'd66842,17'd66843,17'd66844,17'd64838,17'd63715,17'd66845,17'd66846,17'd65348,17'd63034,17'd66847,17'd66594,17'd65869,17'd65998,17'd66848,17'd66849,17'd66850,17'd60216,17'd60344,17'd13626,17'd53969,17'd53180,17'd66851,17'd66852,17'd9736,17'd48491,17'd27002,17'd13886,17'd66853,17'd66854,17'd40595,17'd12867,17'd53836,17'd9889,17'd19034,17'd61353,17'd25815,17'd66855,17'd11283,17'd66856,17'd8433,17'd56625,17'd66857,17'd66858,17'd18576,17'd12273,17'd9495,17'd11977,17'd12275,17'd7813,17'd8132,17'd14276,17'd14276,17'd8132,17'd542,17'd133,17'd133,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd134,17'd1759,17'd128,17'd130,17'd133,17'd133,17'd133,17'd13901,17'd65124,17'd24056,17'd66859,17'd66860,17'd66861,17'd66862,17'd66863,17'd66864,17'd66865,17'd66734,17'd66866,17'd66867,17'd66868,17'd66869,17'd66870,17'd66871,17'd66872,17'd66873,17'd66874,17'd66875,17'd66741,17'd66742,17'd66741,17'd66269,17'd65788,17'd65788,17'd66144,17'd66144,17'd66144,17'd66144,17'd66144,17'd65520,17'd65653,17'd65653,17'd66876,17'd66876,17'd66877,17'd66878,17'd65788,17'd65521,17'd65522,17'd66499,17'd66499,17'd60587,17'd60716,17'd66879,17'd66748,17'd66880,17'd66751,17'd66881,17'd66881,17'd66882,17'd66883,17'd66884,17'd66885,17'd66886,17'd66887,17'd66888,17'd66756,17'd60356,17'd66275,17'd66035,17'd66889,17'd50648,17'd33644,17'd32007,17'd29101,17'd28721,17'd23553,17'd33970,17'd30300,17'd43023,17'd38820,17'd66890,17'd25185,17'd31373,17'd61132,17'd62043,17'd66891,17'd63780,17'd66892,17'd66893,17'd66894,17'd66895,17'd66769,17'd66896,17'd66897,17'd66898,17'd66899,17'd66900,17'd66901,17'd19440,17'd66902,17'd66903,17'd66904,17'd66905,17'd9643,17'd66906,17'd16726,17'd27196,17'd27690,17'd21924,17'd27692,17'd29157,17'd66907,17'd29292,17'd30331,17'd7825,17'd6846,17'd6214,17'd6213,17'd28532,17'd50670,17'd50670,17'd5611,17'd5612,17'd25627,17'd30638,17'd28185,17'd53214,17'd52182,17'd9092,17'd30937,17'd66908,17'd66909,17'd66910,17'd66659,17'd66660,17'd66911,17'd66912,17'd66913,17'd66914,17'd64368,17'd65289,17'd64227,17'd66533,17'd66787,17'd63356,17'd63357,17'd64769,17'd65041,17'd65041,17'd65165,17'd64090,17'd64629,17'd66788,17'd66321,17'd66321,17'd63377,17'd63377,17'd63378,17'd63376,17'd66789,17'd66790,17'd65816,17'd65816,17'd66915,17'd17659,17'd66539,17'd66539,17'd18268,17'd66916,17'd66917,17'd66918,17'd11046,17'd66919,17'd66920,17'd66920,17'd66921,17'd66920,17'd11187,17'd66798,17'd66922,17'd66799,17'd66923,17'd66923,17'd11587,17'd11587,17'd10388,17'd10790,17'd39790,17'd11720,17'd44742,17'd60399,17'd44019,17'd44387,17'd16623,17'd44850,17'd66924,17'd66194,17'd66193,17'd66801,17'd66801,17'd66801,17'd66925,17'd66926,17'd65945,17'd62846,17'd15104,17'd66195,17'd65304,17'd62445,17'd65304,17'd65304,17'd66434,17'd15232,17'd65949,17'd66927,17'd65950,17'd63963,17'd66072,17'd66804,17'd66072,17'd65054,17'd66318,17'd66928,17'd66677,17'd65570,17'd64110,17'd66929,17'd64388,17'd65055,17'd66077,17'd66077,17'd66077,17'd66930,17'd64528,17'd63247,17'd66931,17'd66932,17'd18863,17'd9661,17'd66933,17'd66550,17'd3057,17'd66934,17'd2223,17'd66080,17'd2079,17'd56664,17'd66935,17'd61540
},
'{
17'd3427,17'd3427,17'd3751,17'd3751,17'd3427,17'd3101,17'd14070,17'd3252,17'd3101,17'd2784,17'd10535,17'd10535,17'd2784,17'd63255,17'd63816,17'd65840,17'd66086,17'd66936,17'd66686,17'd66810,17'd66937,17'd66938,17'd66939,17'd66940,17'd66558,17'd66941,17'd66552,17'd65713,17'd66942,17'd63520,17'd65584,17'd1415,17'd19,17'd979,17'd18,17'd19,17'd18,17'd4089,17'd17,17'd22965,17'd2257,17'd2597,17'd3252,17'd3101,17'd4245,17'd3903,17'd4426,17'd4888,17'd5509,17'd5509,17'd14745,17'd7049,17'd5511,17'd15358,17'd10670,17'd10669,17'd10669,17'd10924,17'd471,17'd295,17'd2428,17'd1838,17'd1134,17'd1134,17'd1135,17'd1138,17'd66943,17'd66094,17'd3757,17'd4254,17'd5381,17'd5383,17'd13579,17'd14192,17'd5805,17'd5219,17'd66944,17'd13070,17'd65964,17'd54608,17'd66945,17'd66946,17'd66947,17'd66948,17'd66949,17'd66950,17'd66951,17'd13330,17'd13479,17'd66952,17'd43467,17'd24015,17'd9580,17'd9580,17'd29181,17'd7411,17'd10118,17'd9577,17'd8381,17'd66953,17'd66954,17'd6777,17'd6474,17'd7094,17'd64943,17'd4126,17'd7751,17'd8371,17'd13842,17'd52849,17'd47673,17'd54343,17'd66955,17'd54613,17'd57013,17'd48932,17'd58400,17'd55775,17'd59515,17'd65735,17'd56021,17'd66956,17'd54706,17'd58400,17'd58149,17'd49199,17'd54797,17'd54886,17'd49814,17'd49303,17'd57124,17'd66957,17'd66958,17'd65737,17'd56020,17'd55902,17'd55489,17'd65332,17'd58037,17'd60796,17'd66959,17'd66960,17'd59144,17'd58530,17'd63148,17'd66961,17'd61711,17'd66962,17'd58887,17'd58772,17'd64280,17'd4921,17'd66963,17'd32577,17'd66964,17'd66965,17'd66966,17'd66967,17'd66586,17'd66713,17'd66716,17'd66968,17'd66969,17'd66970,17'd66717,17'd66971,17'd66844,17'd64838,17'd66972,17'd66973,17'd66974,17'd66975,17'd65105,17'd66593,17'd66594,17'd65869,17'd65998,17'd66976,17'd66977,17'd66978,17'd60701,17'd66979,17'd14243,17'd11648,17'd53240,17'd28679,17'd51116,17'd9731,17'd66980,17'd66981,17'd11132,17'd53631,17'd51119,17'd8720,17'd38748,17'd23519,17'd15188,17'd21508,17'd59568,17'd66982,17'd18924,17'd13143,17'd23529,17'd17244,17'd66983,17'd66984,17'd10755,17'd22488,17'd64716,17'd7812,17'd52140,17'd888,17'd888,17'd719,17'd6198,17'd66124,17'd1481,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd11541,17'd20623,17'd20465,17'd21376,17'd22313,17'd66985,17'd66986,17'd66987,17'd66988,17'd66989,17'd66990,17'd66991,17'd66992,17'd66993,17'd66994,17'd66995,17'd66868,17'd64462,17'd64592,17'd64187,17'd60474,17'd66621,17'd66874,17'd59852,17'd59852,17'd66875,17'd66743,17'd66741,17'd65788,17'd66269,17'd66269,17'd66269,17'd65788,17'd65788,17'd66269,17'd65898,17'd66996,17'd66997,17'd66138,17'd66145,17'd66499,17'd66998,17'd66621,17'd63895,17'd66747,17'd66999,17'd67000,17'd67001,17'd67002,17'd62522,17'd66881,17'd67003,17'd67004,17'd67005,17'd67006,17'd67007,17'd66887,17'd67008,17'd50558,17'd67009,17'd60717,17'd62784,17'd57833,17'd59085,17'd57707,17'd34106,17'd32007,17'd25320,17'd28484,17'd25435,17'd67010,17'd39141,17'd30149,17'd30447,17'd35995,17'd27263,17'd67011,17'd60739,17'd67012,17'd67013,17'd67014,17'd66766,17'd67015,17'd66894,17'd67016,17'd67017,17'd67018,17'd67019,17'd67020,17'd67021,17'd67022,17'd66648,17'd67023,17'd65674,17'd67024,17'd67025,17'd67026,17'd67027,17'd18357,17'd16112,17'd67028,17'd25480,17'd21451,17'd21924,17'd21142,17'd12741,17'd10198,17'd52521,17'd7990,17'd7825,17'd6213,17'd8931,17'd6552,17'd27930,17'd5612,17'd5612,17'd5158,17'd5331,17'd5158,17'd5159,17'd5614,17'd6708,17'd35760,17'd9092,17'd66419,17'd66657,17'd67029,17'd67030,17'd67031,17'd67032,17'd67033,17'd66912,17'd67034,17'd67035,17'd66064,17'd66064,17'd66180,17'd63940,17'd67036,17'd24660,17'd25232,17'd63940,17'd67037,17'd64089,17'd66180,17'd65289,17'd65688,17'd65286,17'd64109,17'd65570,17'd65570,17'd64109,17'd63244,17'd63108,17'd66078,17'd66078,17'd66322,17'd66322,17'd16255,17'd67038,17'd67039,17'd67039,17'd14059,17'd66932,17'd18628,17'd18382,17'd63111,17'd12316,17'd12316,17'd63111,17'd63111,17'd62071,17'd67040,17'd63659,17'd10905,17'd67041,17'd66923,17'd67042,17'd67043,17'd66674,17'd40716,17'd11188,17'd11720,17'd50186,17'd12176,17'd60399,17'd12913,17'd44387,17'd16623,17'd65700,17'd66194,17'd66926,17'd67044,17'd67045,17'd67044,17'd67046,17'd67047,17'd67048,17'd65700,17'd15735,17'd15104,17'd14584,17'd65304,17'd62445,17'd65565,17'd65565,17'd66434,17'd15348,17'd62699,17'd62849,17'd66197,17'd67049,17'd66437,17'd65569,17'd66072,17'd66072,17'd66072,17'd66072,17'd66677,17'd66677,17'd67050,17'd66929,17'd64921,17'd66320,17'd67051,17'd67051,17'd65831,17'd67052,17'd67053,17'd66322,17'd62976,17'd18382,17'd10387,17'd67054,17'd67055,17'd66550,17'd3057,17'd67056,17'd67057,17'd67058,17'd62335,17'd57358,17'd67059,17'd67060
},
'{
17'd3427,17'd3427,17'd3751,17'd3751,17'd2934,17'd3101,17'd14070,17'd3252,17'd3101,17'd2422,17'd10535,17'd17917,17'd2422,17'd63255,17'd67061,17'd67062,17'd66086,17'd66936,17'd66686,17'd66810,17'd66937,17'd66938,17'd66939,17'd67063,17'd67064,17'd66559,17'd66327,17'd65582,17'd13815,17'd6433,17'd63260,17'd2936,17'd16,17'd3748,17'd19,17'd19,17'd18,17'd3905,17'd16,17'd1416,17'd2257,17'd2257,17'd1831,17'd2935,17'd4245,17'd4088,17'd3902,17'd4734,17'd5509,17'd5509,17'd67065,17'd7049,17'd5511,17'd15496,17'd10925,17'd10669,17'd10669,17'd10802,17'd984,17'd811,17'd13578,17'd2428,17'd1838,17'd1281,17'd1281,17'd1137,17'd67066,17'd67067,17'd2434,17'd4255,17'd5381,17'd5807,17'd67068,17'd67069,17'd14192,17'd5805,17'd13069,17'd13438,17'd67070,17'd65965,17'd67071,17'd67072,17'd67073,17'd67074,17'd67075,17'd67076,17'd17695,17'd67077,17'd13217,17'd13608,17'd19899,17'd67078,17'd9989,17'd9989,17'd24198,17'd10432,17'd10696,17'd9578,17'd67079,17'd8071,17'd67080,17'd6637,17'd6639,17'd7754,17'd7097,17'd6933,17'd3952,17'd58393,17'd58394,17'd52849,17'd47673,17'd15900,17'd66955,17'd54613,17'd57013,17'd57504,17'd57772,17'd58150,17'd65734,17'd65735,17'd56021,17'd56020,17'd54993,17'd65733,17'd58272,17'd57504,17'd49199,17'd56569,17'd32260,17'd54797,17'd67081,17'd67082,17'd67082,17'd66958,17'd57773,17'd54895,17'd67083,17'd67084,17'd58042,17'd67085,17'd59935,17'd56459,17'd67086,17'd67086,17'd56459,17'd61063,17'd67087,17'd67088,17'd64287,17'd67089,17'd55285,17'd67090,17'd65976,17'd33706,17'd67091,17'd67092,17'd67093,17'd66967,17'd67094,17'd67095,17'd67096,17'd66968,17'd66969,17'd66970,17'd66717,17'd66843,17'd66236,17'd64838,17'd63713,17'd67097,17'd67098,17'd67099,17'd67100,17'd66593,17'd66594,17'd65869,17'd65998,17'd66239,17'd67101,17'd67102,17'd60088,17'd67103,17'd57054,17'd12239,17'd53384,17'd51955,17'd50947,17'd67104,17'd28341,17'd40603,17'd11400,17'd20610,17'd21205,17'd9346,17'd12725,17'd17850,17'd16802,17'd13377,17'd14389,17'd62007,17'd55321,17'd15954,17'd14396,17'd67105,17'd67106,17'd23358,17'd22838,17'd11977,17'd16811,17'd7813,17'd888,17'd889,17'd542,17'd719,17'd356,17'd4163,17'd1481,17'd1481,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd65123,17'd67107,17'd66859,17'd66985,17'd67108,17'd66730,17'd67109,17'd67110,17'd67111,17'd66490,17'd67112,17'd67113,17'd67114,17'd67115,17'd67116,17'd62397,17'd67117,17'd64186,17'd64049,17'd67118,17'd67119,17'd67120,17'd63895,17'd66874,17'd67121,17'd65896,17'd66743,17'd66743,17'd66741,17'd66269,17'd65788,17'd65521,17'd65521,17'd66138,17'd58816,17'd67122,17'd66621,17'd66500,17'd66622,17'd66747,17'd67120,17'd66999,17'd64594,17'd67001,17'd67002,17'd62522,17'd67123,17'd63328,17'd63195,17'd67124,17'd67125,17'd67126,17'd67127,17'd67128,17'd67129,17'd67009,17'd67130,17'd60475,17'd60356,17'd67131,17'd64730,17'd57707,17'd48987,17'd24895,17'd25178,17'd28850,17'd28484,17'd36716,17'd29547,17'd36135,17'd30893,17'd36411,17'd67132,17'd67133,17'd67134,17'd67135,17'd25206,17'd23422,17'd67136,17'd67137,17'd67138,17'd67139,17'd67140,17'd67141,17'd66771,17'd17877,17'd67142,17'd67143,17'd67022,17'd67144,17'd67145,17'd67146,17'd67147,17'd67148,17'd18719,17'd67149,17'd15591,17'd16478,17'd17894,17'd25480,17'd25765,17'd67150,17'd20992,17'd21143,17'd28904,17'd9219,17'd7167,17'd7991,17'd8931,17'd7667,17'd6552,17'd5761,17'd5158,17'd5158,17'd5158,17'd26218,17'd5159,17'd32243,17'd6390,17'd7178,17'd67151,17'd67152,17'd67153,17'd67154,17'd67155,17'd67156,17'd67157,17'd67158,17'd67159,17'd67160,17'd67161,17'd64226,17'd64227,17'd66064,17'd67037,17'd63940,17'd26956,17'd24660,17'd67162,17'd63940,17'd67037,17'd66180,17'd66180,17'd64369,17'd64507,17'd66788,17'd64527,17'd65305,17'd65570,17'd65570,17'd63808,17'd63808,17'd63510,17'd66078,17'd67163,17'd67163,17'd65705,17'd66679,17'd13687,17'd67164,17'd12912,17'd64924,17'd64924,17'd13175,17'd13175,17'd13570,17'd13570,17'd67165,17'd12771,17'd61941,17'd67166,17'd67167,17'd11586,17'd67168,17'd67043,17'd67043,17'd11047,17'd66674,17'd11188,17'd11587,17'd11720,17'd12318,17'd12176,17'd44019,17'd44387,17'd63960,17'd44850,17'd65945,17'd66194,17'd66926,17'd67044,17'd67045,17'd67044,17'd67046,17'd66926,17'd67169,17'd62846,17'd15862,17'd66195,17'd63653,17'd65304,17'd62445,17'd65947,17'd66434,17'd15103,17'd15483,17'd62849,17'd63107,17'd63963,17'd66073,17'd66677,17'd66677,17'd66072,17'd66072,17'd66072,17'd66437,17'd66677,17'd67170,17'd66929,17'd67171,17'd67172,17'd66320,17'd67051,17'd66077,17'd65055,17'd63809,17'd63376,17'd65705,17'd67173,17'd67174,17'd67175,17'd48639,17'd67176,17'd62704,17'd53516,17'd66934,17'd67177,17'd67178,17'd62335,17'd53434,17'd58987,17'd67060
},
'{
17'd3427,17'd3427,17'd3751,17'd2934,17'd3101,17'd3101,17'd3252,17'd2422,17'd3252,17'd1688,17'd2594,17'd17917,17'd10535,17'd2784,17'd63665,17'd65582,17'd67179,17'd66326,17'd66686,17'd66810,17'd67180,17'd67181,17'd67063,17'd67063,17'd66940,17'd67182,17'd66207,17'd67183,17'd64254,17'd64799,17'd10923,17'd9815,17'd15,17'd5051,17'd1276,17'd1277,17'd19,17'd18,17'd18,17'd3905,17'd1416,17'd2257,17'd1831,17'd3252,17'd2935,17'd3751,17'd4892,17'd5646,17'd6263,17'd5509,17'd5052,17'd4734,17'd15359,17'd15496,17'd10925,17'd11071,17'd10669,17'd10802,17'd10802,17'd984,17'd13303,17'd2261,17'd2121,17'd1557,17'd1282,17'd1135,17'd67066,17'd66943,17'd67184,17'd4255,17'd5381,17'd5383,17'd12200,17'd5974,17'd67069,17'd14192,17'd5382,17'd66944,17'd66820,17'd34346,17'd63121,17'd67185,17'd67186,17'd67187,17'd67188,17'd67189,17'd67190,17'd13847,17'd66455,17'd67191,17'd67192,17'd43346,17'd11092,17'd10949,17'd20436,17'd9705,17'd22635,17'd9705,17'd66113,17'd65595,17'd7916,17'd67080,17'd51100,17'd67193,17'd7258,17'd7089,17'd4126,17'd4292,17'd58882,17'd65858,17'd14624,17'd47673,17'd48079,17'd67194,17'd56232,17'd48931,17'd58272,17'd58400,17'd65734,17'd67195,17'd65735,17'd57014,17'd65735,17'd57268,17'd65981,17'd58272,17'd48820,17'd49199,17'd55373,17'd54797,17'd56801,17'd57386,17'd57385,17'd57013,17'd50094,17'd67196,17'd67197,17'd67198,17'd67199,17'd67200,17'd67201,17'd67202,17'd60793,17'd67203,17'd67204,17'd59399,17'd1321,17'd60060,17'd58661,17'd66575,17'd67205,17'd67206,17'd67207,17'd33864,17'd67208,17'd67092,17'd67209,17'd67210,17'd67094,17'd67095,17'd67211,17'd67212,17'd67213,17'd66970,17'd67214,17'd66843,17'd66236,17'd67215,17'd63712,17'd67216,17'd67098,17'd67217,17'd67218,17'd67219,17'd66594,17'd65869,17'd65869,17'd66239,17'd67101,17'd64574,17'd59689,17'd58685,17'd67220,17'd12701,17'd11253,17'd51784,17'd10453,17'd67221,17'd9730,17'd67222,17'd10330,17'd12721,17'd21205,17'd11809,17'd9744,17'd18203,17'd15192,17'd67223,17'd14388,17'd55420,17'd67224,17'd67225,17'd67226,17'd67227,17'd67228,17'd67229,17'd11977,17'd888,17'd888,17'd889,17'd542,17'd133,17'd133,17'd133,17'd133,17'd133,17'd1481,17'd1481,17'd133,17'd133,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd134,17'd131,17'd131,17'd67230,17'd67231,17'd66859,17'd21222,17'd67232,17'd66861,17'd67233,17'd67234,17'd67235,17'd67236,17'd67237,17'd67238,17'd67239,17'd67240,17'd67241,17'd67242,17'd67243,17'd67244,17'd67245,17'd67246,17'd67247,17'd66879,17'd64594,17'd64868,17'd60474,17'd66621,17'd66621,17'd66621,17'd66998,17'd66998,17'd66998,17'd66998,17'd60106,17'd66874,17'd63895,17'd63895,17'd67118,17'd66999,17'd64594,17'd64594,17'd66748,17'd67002,17'd66880,17'd67123,17'd66882,17'd67124,17'd63054,17'd67248,17'd67125,17'd67249,17'd50557,17'd67250,17'd67251,17'd67252,17'd67253,17'd67254,17'd60717,17'd66757,17'd67255,17'd59207,17'd67256,17'd50363,17'd30126,17'd28596,17'd25177,17'd28484,17'd40379,17'd59089,17'd30893,17'd67257,17'd30150,17'd67258,17'd67259,17'd67260,17'd67261,17'd67262,17'd67263,17'd22894,17'd67264,17'd67265,17'd67266,17'd67267,17'd67268,17'd67269,17'd67270,17'd67271,17'd67272,17'd67273,17'd67022,17'd67274,17'd67275,17'd67275,17'd66904,17'd67276,17'd67277,17'd10887,17'd66906,17'd17051,17'd17894,17'd24940,17'd21924,17'd21610,17'd21611,17'd12884,17'd67278,17'd7990,17'd6703,17'd6214,17'd7667,17'd8932,17'd9523,17'd26218,17'd26218,17'd26218,17'd30638,17'd28185,17'd28185,17'd6554,17'd6708,17'd7011,17'd8631,17'd67152,17'd67279,17'd67280,17'd67281,17'd67282,17'd67032,17'd67283,17'd67160,17'd67284,17'd64505,17'd63940,17'd64227,17'd66180,17'd67037,17'd67285,17'd67036,17'd24660,17'd67036,17'd64226,17'd67286,17'd66180,17'd65815,17'd67287,17'd65039,17'd63377,17'd65570,17'd66677,17'd66677,17'd66677,17'd66676,17'd66073,17'd63375,17'd62971,17'd65441,17'd65441,17'd17179,17'd67288,17'd67289,17'd67290,17'd67290,17'd62576,17'd14583,17'd62447,17'd62447,17'd67291,17'd67291,17'd13688,17'd13688,17'd67292,17'd12634,17'd18511,17'd12016,17'd18511,17'd63659,17'd67041,17'd10247,17'd11047,17'd11587,17'd67293,17'd50756,17'd12318,17'd60399,17'd12913,17'd43596,17'd16132,17'd65700,17'd66194,17'd67047,17'd67047,17'd67044,17'd67044,17'd67044,17'd66926,17'd67294,17'd62846,17'd15735,17'd15862,17'd66195,17'd65304,17'd65304,17'd65565,17'd66434,17'd15103,17'd15232,17'd16959,17'd65950,17'd63243,17'd64919,17'd66437,17'd65570,17'd65570,17'd66072,17'd66072,17'd66072,17'd66437,17'd65703,17'd67170,17'd66929,17'd67171,17'd67295,17'd67296,17'd67051,17'd66077,17'd64653,17'd63658,17'd66790,17'd62702,17'd67297,17'd10387,17'd7511,17'd3865,17'd67176,17'd62704,17'd2542,17'd67298,17'd67299,17'd67300,17'd67301,17'd53434,17'd59616,17'd59121
},
'{
17'd3427,17'd3427,17'd3751,17'd3751,17'd2934,17'd2935,17'd3252,17'd2422,17'd3252,17'd1689,17'd4247,17'd15745,17'd17917,17'd2935,17'd67302,17'd65581,17'd67179,17'd66328,17'd66686,17'd66810,17'd67303,17'd67181,17'd66940,17'd67304,17'd66812,17'd66940,17'd66330,17'd65957,17'd67305,17'd67306,17'd63668,17'd63257,17'd14742,17'd67307,17'd67308,17'd1277,17'd979,17'd18,17'd3905,17'd18,17'd1416,17'd1414,17'd1688,17'd2422,17'd2935,17'd2593,17'd4428,17'd4891,17'd6263,17'd5509,17'd5052,17'd4888,17'd15359,17'd5204,17'd11888,17'd10924,17'd10669,17'd10669,17'd10802,17'd10802,17'd656,17'd2939,17'd1972,17'd1972,17'd16966,17'd1281,17'd67066,17'd67066,17'd14194,17'd3913,17'd5381,17'd5807,17'd5974,17'd5974,17'd67068,17'd67069,17'd13579,17'd13579,17'd5057,17'd33850,17'd54608,17'd67309,17'd63392,17'd67310,17'd67311,17'd67312,17'd67313,17'd16988,17'd67314,17'd67315,17'd19761,17'd67192,17'd11766,17'd66699,17'd10698,17'd20435,17'd67316,17'd9705,17'd24522,17'd65855,17'd8380,17'd8377,17'd7099,17'd7258,17'd7096,17'd7089,17'd6933,17'd4126,17'd59265,17'd58517,17'd58269,17'd16031,17'd48078,17'd57632,17'd56343,17'd56232,17'd53950,17'd48932,17'd58150,17'd54346,17'd65735,17'd67317,17'd67318,17'd55185,17'd54894,17'd54172,17'd48932,17'd48931,17'd53080,17'd49814,17'd56801,17'd56801,17'd57266,17'd57636,17'd34179,17'd55897,17'd58518,17'd67319,17'd57015,17'd56132,17'd61190,17'd59020,17'd67320,17'd67321,17'd67322,17'd60180,17'd67323,17'd55681,17'd67324,17'd59524,17'd58152,17'd66706,17'd67325,17'd67326,17'd67327,17'd67328,17'd67329,17'd67330,17'd67331,17'd67210,17'd67332,17'd67333,17'd67334,17'd67335,17'd67336,17'd67337,17'd67338,17'd67339,17'd67340,17'd67341,17'd67342,17'd67343,17'd67100,17'd67219,17'd66594,17'd67344,17'd65869,17'd67345,17'd67346,17'd67347,17'd62003,17'd58068,17'd11497,17'd16429,17'd67348,17'd67349,17'd32912,17'd50606,17'd67350,17'd47596,17'd17719,17'd10478,17'd13886,17'd16070,17'd8570,17'd25290,17'd11534,17'd67223,17'd22301,17'd67351,17'd67352,17'd23879,17'd67353,17'd67354,17'd10619,17'd67355,17'd7813,17'd889,17'd542,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd133,17'd1481,17'd1481,17'd133,17'd133,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd131,17'd131,17'd20466,17'd67356,17'd67357,17'd67358,17'd67359,17'd67360,17'd67361,17'd67362,17'd67363,17'd67364,17'd67365,17'd67366,17'd67367,17'd67368,17'd67369,17'd67370,17'd67371,17'd67372,17'd67373,17'd67374,17'd67374,17'd67247,17'd67002,17'd66750,17'd66749,17'd66879,17'd67000,17'd66999,17'd67120,17'd66747,17'd66747,17'd66747,17'd66747,17'd66747,17'd67375,17'd67376,17'd67247,17'd67001,17'd67002,17'd67377,17'd62522,17'd67123,17'd66881,17'd63195,17'd67378,17'd67379,17'd67380,17'd67381,17'd67382,17'd67383,17'd67384,17'd67251,17'd67383,17'd67253,17'd67385,17'd62399,17'd62784,17'd66034,17'd64468,17'd58582,17'd50363,17'd29688,17'd24897,17'd28719,17'd25709,17'd27765,17'd40379,17'd60362,17'd67386,17'd37133,17'd34763,17'd25039,17'd67387,17'd67388,17'd67389,17'd67390,17'd67391,17'd67392,17'd67393,17'd67394,17'd67395,17'd67396,17'd67397,17'd67398,17'd67399,17'd67400,17'd67401,17'd67402,17'd67403,17'd67404,17'd67405,17'd67406,17'd67276,17'd67407,17'd11019,17'd10768,17'd66906,17'd17055,17'd25876,17'd67408,17'd67409,17'd67410,17'd67411,17'd20993,17'd9068,17'd7169,17'd6214,17'd8931,17'd8779,17'd7999,17'd6553,17'd6389,17'd26218,17'd28185,17'd30638,17'd31717,17'd6554,17'd32073,17'd7177,17'd67412,17'd8935,17'd67413,17'd67414,17'd67415,17'd67416,17'd67031,17'd67417,17'd67418,17'd67419,17'd67420,17'd64628,17'd67037,17'd64089,17'd67037,17'd67037,17'd66533,17'd67162,17'd67162,17'd67285,17'd64226,17'd64368,17'd66063,17'd65164,17'd67421,17'd67422,17'd63377,17'd65703,17'd67423,17'd66677,17'd67423,17'd66676,17'd64651,17'd62971,17'd67424,17'd67425,17'd67425,17'd67426,17'd67426,17'd15618,17'd67427,17'd67427,17'd15618,17'd15483,17'd15999,17'd15103,17'd66434,17'd67428,17'd67429,17'd67430,17'd67430,17'd18033,17'd18140,17'd18511,17'd18511,17'd67168,17'd67041,17'd67041,17'd67043,17'd67293,17'd67431,17'd50756,17'd44966,17'd44019,17'd63959,17'd16132,17'd15735,17'd66070,17'd66926,17'd67432,17'd67047,17'd67044,17'd67044,17'd67044,17'd67433,17'd67434,17'd15862,17'd62574,17'd62575,17'd63653,17'd65565,17'd65565,17'd65565,17'd15103,17'd15103,17'd15483,17'd67435,17'd63107,17'd63655,17'd66072,17'd66804,17'd65570,17'd65305,17'd66072,17'd66072,17'd66072,17'd66437,17'd65703,17'd67050,17'd67436,17'd67295,17'd67437,17'd67438,17'd67439,17'd66077,17'd63809,17'd67440,17'd66322,17'd62855,17'd62452,17'd66795,17'd4862,17'd65442,17'd67441,17'd62704,17'd51182,17'd37818,17'd53290,17'd53515,17'd67442,17'd67443,17'd59121,17'd59121
},
'{
17'd3427,17'd3427,17'd3751,17'd2934,17'd3101,17'd2935,17'd2422,17'd2422,17'd2422,17'd1689,17'd1127,17'd15745,17'd17917,17'd14070,17'd67444,17'd67445,17'd65844,17'd66327,17'd67446,17'd66810,17'd67303,17'd66937,17'd67447,17'd67448,17'd67449,17'd67063,17'd66559,17'd67450,17'd12191,17'd13064,17'd64798,17'd67451,17'd63386,17'd67452,17'd67453,17'd4884,17'd19,17'd19,17'd26127,17'd3905,17'd1416,17'd1416,17'd1414,17'd3429,17'd2784,17'd2784,17'd2934,17'd4244,17'd5197,17'd10397,17'd5052,17'd4888,17'd15359,17'd5511,17'd3592,17'd2934,17'd10669,17'd10669,17'd10669,17'd10802,17'd656,17'd3103,17'd1973,17'd2122,17'd2600,17'd1557,17'd14449,17'd1284,17'd2268,17'd3913,17'd5220,17'd5659,17'd5975,17'd67454,17'd67455,17'd5974,17'd12200,17'd5807,17'd5381,17'd66214,17'd3440,17'd67456,17'd67457,17'd67458,17'd67459,17'd67460,17'd67461,17'd46994,17'd67462,17'd18785,17'd67463,17'd67192,17'd11482,17'd67464,17'd11235,17'd10698,17'd10120,17'd9843,17'd9578,17'd67465,17'd65855,17'd8847,17'd8073,17'd8070,17'd7258,17'd7258,17'd67466,17'd6934,17'd4124,17'd59512,17'd65858,17'd58269,17'd66347,17'd48079,17'd48080,17'd55373,17'd56232,17'd53950,17'd58400,17'd55775,17'd56021,17'd57014,17'd54799,17'd57014,17'd57126,17'd65733,17'd65981,17'd66107,17'd57504,17'd56125,17'd49814,17'd55373,17'd32260,17'd32260,17'd34178,17'd34178,17'd50094,17'd54020,17'd63542,17'd56027,17'd55486,17'd67467,17'd67468,17'd67469,17'd63282,17'd58531,17'd67470,17'd67471,17'd60792,17'd61449,17'd67472,17'd60167,17'd67473,17'd67474,17'd67475,17'd67476,17'd67329,17'd67477,17'd67478,17'd67479,17'd67480,17'd67333,17'd67334,17'd66970,17'd67214,17'd67481,17'd67482,17'd67483,17'd67340,17'd67341,17'd67484,17'd67485,17'd67218,17'd67219,17'd66594,17'd67344,17'd65869,17'd67345,17'd67486,17'd67487,17'd67488,17'd13491,17'd67489,17'd11646,17'd15165,17'd29319,17'd30826,17'd50690,17'd67490,17'd47689,17'd9740,17'd20756,17'd14518,17'd26759,17'd67491,17'd25680,17'd9485,17'd38903,17'd56167,17'd67492,17'd18094,17'd66368,17'd67493,17'd67494,17'd8131,17'd717,17'd133,17'd1197,17'd133,17'd133,17'd133,17'd132,17'd131,17'd131,17'd132,17'd132,17'd133,17'd133,17'd1481,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd134,17'd132,17'd131,17'd11541,17'd132,17'd132,17'd134,17'd20625,17'd67495,17'd67496,17'd67497,17'd67498,17'd67499,17'd67500,17'd67501,17'd67502,17'd67503,17'd67504,17'd67505,17'd67506,17'd67507,17'd67508,17'd67509,17'd67510,17'd67511,17'd63751,17'd67372,17'd67512,17'd67513,17'd67123,17'd67514,17'd63752,17'd62275,17'd66751,17'd66880,17'd67515,17'd67516,17'd67001,17'd67515,17'd67002,17'd67377,17'd67377,17'd67517,17'd67123,17'd66881,17'd63328,17'd67518,17'd67005,17'd67519,17'd67125,17'd67249,17'd50557,17'd67250,17'd67384,17'd67520,17'd67521,17'd67383,17'd67251,17'd67522,17'd67254,17'd62525,17'd66630,17'd57833,17'd59085,17'd67256,17'd63762,17'd34621,17'd24744,17'd25029,17'd25438,17'd28369,17'd25567,17'd25436,17'd38820,17'd28014,17'd67523,17'd67524,17'd67525,17'd67526,17'd67527,17'd67528,17'd23767,17'd67529,17'd63352,17'd67530,17'd67140,17'd67531,17'd67532,17'd67533,17'd67534,17'd67535,17'd67536,17'd67537,17'd67402,17'd67538,17'd67539,17'd67540,17'd67541,17'd67407,17'd10366,17'd18357,17'd16473,17'd66906,17'd16729,17'd26110,17'd21451,17'd21452,17'd27693,17'd12444,17'd10499,17'd8290,17'd6847,17'd6215,17'd7667,17'd7999,17'd7999,17'd8303,17'd26708,17'd31717,17'd6554,17'd50282,17'd53214,17'd6853,17'd7178,17'd6557,17'd7836,17'd67152,17'd67542,17'd67543,17'd67544,17'd67545,17'd67546,17'd67547,17'd67548,17'd67549,17'd67550,17'd64226,17'd67551,17'd67037,17'd67286,17'd67037,17'd66533,17'd25232,17'd25232,17'd67552,17'd64628,17'd65038,17'd67287,17'd67422,17'd66321,17'd67422,17'd63658,17'd67170,17'd67553,17'd66677,17'd66677,17'd66676,17'd63655,17'd62970,17'd67554,17'd67555,17'd67555,17'd66803,17'd15103,17'd15348,17'd15348,17'd15348,17'd15232,17'd15232,17'd15103,17'd66434,17'd66803,17'd65948,17'd65948,17'd66071,17'd66071,17'd65946,17'd13055,17'd12482,17'd67293,17'd67556,17'd11047,17'd67043,17'd67043,17'd67431,17'd50756,17'd44966,17'd44966,17'd44019,17'd62444,17'd15735,17'd66924,17'd66194,17'd67047,17'd67045,17'd67044,17'd67044,17'd67044,17'd67433,17'd67433,17'd67169,17'd62574,17'd62444,17'd63653,17'd63653,17'd65565,17'd65565,17'd67291,17'd67557,17'd67557,17'd16959,17'd62850,17'd63243,17'd64651,17'd66437,17'd66677,17'd65305,17'd65305,17'd66072,17'd66072,17'd66072,17'd66437,17'd65703,17'd67050,17'd64789,17'd66320,17'd67438,17'd67558,17'd67559,17'd67560,17'd63657,17'd63376,17'd65705,17'd12481,17'd11046,17'd67561,17'd46698,17'd2889,17'd67441,17'd53744,17'd53291,17'd53147,17'd67562,17'd67563,17'd67564,17'd67565,17'd61541,17'd58861
},
'{
17'd3427,17'd3427,17'd3751,17'd3751,17'd2934,17'd2935,17'd2422,17'd3250,17'd2422,17'd1967,17'd1127,17'd2595,17'd2594,17'd14070,17'd63385,17'd67566,17'd67567,17'd66327,17'd67446,17'd67568,17'd67569,17'd66937,17'd67570,17'd67448,17'd67571,17'd67572,17'd67573,17'd66089,17'd8344,17'd67574,17'd67575,17'd67576,17'd11736,17'd6274,17'd67577,17'd14319,17'd1277,17'd19,17'd20404,17'd20404,17'd3905,17'd17,17'd1414,17'd2597,17'd2422,17'd2784,17'd2593,17'd4428,17'd4890,17'd5198,17'd5052,17'd6263,17'd7049,17'd5203,17'd5204,17'd3901,17'd11071,17'd10669,17'd10669,17'd10669,17'd656,17'd656,17'd2260,17'd2122,17'd2600,17'd2121,17'd1556,17'd14449,17'd2123,17'd3912,17'd5214,17'd5808,17'd6109,17'd67454,17'd67454,17'd67454,17'd12786,17'd12786,17'd5383,17'd12338,17'd3758,17'd67578,17'd66822,17'd67579,17'd67580,17'd67581,17'd67582,17'd67583,17'd67584,17'd67585,17'd67586,17'd14487,17'd12368,17'd12367,17'd11766,17'd12068,17'd20436,17'd9843,17'd9987,17'd24522,17'd24522,17'd9441,17'd8847,17'd8072,17'd8375,17'd7097,17'd67587,17'd67587,17'd4463,17'd59265,17'd58393,17'd65858,17'd66347,17'd47864,17'd47971,17'd48080,17'd56343,17'd55483,17'd58272,17'd58649,17'd55900,17'd56020,17'd64419,17'd54701,17'd64824,17'd54705,17'd54894,17'd65981,17'd58272,17'd48931,17'd55483,17'd56343,17'd32100,17'd32100,17'd54797,17'd54797,17'd56569,17'd49303,17'd67588,17'd55185,17'd55674,17'd67589,17'd67590,17'd60178,17'd67591,17'd61062,17'd55494,17'd63410,17'd67592,17'd63148,17'd67593,17'd54707,17'd61565,17'd67594,17'd67595,17'd67596,17'd67329,17'd67597,17'd67598,17'd67096,17'd67599,17'd67600,17'd67334,17'd67335,17'd67601,17'd67337,17'd66971,17'd67483,17'd67602,17'd62376,17'd67484,17'd67603,17'd67604,17'd67219,17'd66594,17'd67344,17'd65869,17'd67345,17'd67605,17'd66977,17'd67606,17'd13621,17'd67607,17'd14510,17'd15165,17'd29059,17'd67608,17'd67609,17'd9725,17'd67610,17'd17011,17'd15688,17'd10606,17'd14928,17'd28584,17'd52223,17'd13768,17'd67611,17'd8427,17'd67612,17'd10753,17'd67613,17'd16578,17'd22312,17'd542,17'd542,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd133,17'd1481,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd134,17'd132,17'd132,17'd131,17'd21376,17'd51716,17'd67614,17'd21071,17'd67615,17'd51809,17'd67616,17'd67617,17'd67618,17'd67619,17'd67620,17'd67621,17'd67370,17'd67508,17'd67622,17'd67622,17'd67623,17'd67624,17'd67625,17'd63601,17'd67626,17'd67627,17'd63328,17'd63054,17'd67628,17'd66886,17'd66885,17'd66884,17'd66753,17'd63195,17'd63328,17'd63328,17'd63054,17'd63054,17'd63054,17'd62926,17'd67628,17'd67379,17'd67126,17'd67249,17'd67128,17'd67128,17'd67384,17'd67629,17'd67629,17'd67629,17'd67629,17'd67629,17'd67383,17'd67630,17'd67631,17'd67632,17'd66275,17'd63899,17'd59582,17'd67633,17'd57076,17'd48987,17'd30126,17'd24896,17'd28254,17'd27882,17'd27765,17'd27882,17'd34127,17'd30598,17'd37260,17'd61003,17'd67634,17'd59881,17'd44840,17'd67635,17'd67636,17'd67637,17'd62952,17'd66643,17'd67638,17'd67639,17'd67640,17'd67641,17'd67642,17'd17504,17'd67643,17'd67644,17'd67645,17'd67646,17'd67647,17'd67648,17'd67649,17'd67650,17'd12607,17'd67651,17'd67652,17'd17393,17'd66906,17'd17055,17'd25480,17'd67408,17'd67653,17'd20531,17'd20689,17'd67654,17'd7827,17'd6550,17'd7667,17'd7667,17'd7999,17'd8000,17'd8303,17'd26708,17'd6554,17'd53214,17'd52182,17'd35760,17'd7178,17'd7177,17'd8001,17'd7836,17'd67655,17'd67656,17'd67657,17'd67658,17'd67659,17'd67660,17'd67661,17'd67662,17'd67663,17'd67664,17'd67286,17'd67551,17'd67037,17'd67286,17'd67037,17'd64089,17'd67665,17'd25232,17'd67552,17'd65552,17'd65815,17'd67421,17'd64109,17'd64109,17'd66321,17'd63658,17'd67666,17'd67667,17'd66677,17'd66677,17'd66073,17'd66435,17'd65950,17'd66927,17'd15999,17'd67668,17'd66803,17'd66434,17'd15103,17'd15232,17'd15103,17'd66434,17'd66803,17'd66803,17'd66803,17'd66803,17'd66803,17'd66803,17'd13932,17'd13932,17'd13571,17'd13571,17'd12482,17'd11442,17'd67556,17'd11327,17'd67043,17'd11442,17'd12318,17'd67669,17'd12635,17'd64918,17'd63959,17'd62574,17'd67670,17'd66070,17'd66926,17'd67047,17'd67044,17'd67044,17'd67044,17'd67044,17'd67433,17'd63104,17'd15862,17'd64649,17'd62445,17'd63653,17'd65947,17'd65565,17'd13688,17'd67557,17'd67557,17'd67426,17'd62850,17'd62971,17'd63655,17'd65305,17'd66677,17'd66677,17'd65305,17'd65305,17'd66072,17'd66072,17'd66437,17'd67671,17'd64529,17'd65306,17'd65055,17'd67296,17'd67672,17'd67673,17'd67674,17'd67675,17'd63377,17'd66678,17'd62702,17'd67676,17'd67677,17'd46882,17'd65939,17'd42195,17'd62704,17'd61674,17'd51016,17'd40407,17'd67678,17'd67679,17'd67680,17'd56329,17'd58861,17'd67681
},
'{
17'd3427,17'd3427,17'd3751,17'd2934,17'd3101,17'd2935,17'd2422,17'd1831,17'd1688,17'd14,17'd466,17'd2595,17'd4247,17'd3252,17'd63813,17'd67682,17'd67683,17'd67684,17'd67685,17'd67686,17'd67687,17'd67688,17'd67689,17'd67448,17'd67690,17'd67690,17'd67691,17'd67692,17'd8513,17'd11885,17'd64255,17'd64124,17'd67693,17'd67694,17'd8042,17'd67695,17'd1277,17'd979,17'd11,17'd20404,17'd3905,17'd17,17'd1414,17'd2597,17'd3752,17'd3429,17'd2935,17'd3751,17'd5201,17'd5053,17'd5052,17'd5052,17'd7049,17'd15359,17'd5204,17'd3592,17'd2593,17'd2593,17'd10669,17'd10669,17'd1130,17'd1130,17'd3103,17'd2262,17'd3103,17'd1973,17'd20405,17'd17919,17'd2267,17'd2948,17'd5214,17'd5660,17'd12337,17'd11737,17'd11890,17'd11737,17'd5976,17'd5975,17'd5384,17'd67696,17'd30348,17'd29615,17'd67697,17'd67698,17'd67699,17'd67700,17'd63831,17'd67701,17'd63837,17'd67702,17'd67703,17'd67704,17'd13481,17'd67705,17'd66952,17'd11766,17'd42348,17'd65974,17'd9843,17'd9843,17'd9705,17'd9578,17'd28669,17'd8847,17'd8070,17'd7421,17'd6637,17'd64140,17'd4463,17'd4124,17'd58393,17'd48190,17'd58266,17'd66347,17'd47973,17'd47971,17'd48080,17'd48821,17'd53810,17'd54172,17'd55776,17'd54893,17'd54803,17'd54799,17'd65081,17'd66830,17'd55775,17'd58400,17'd54172,17'd58272,17'd55576,17'd55483,17'd57123,17'd67194,17'd67706,17'd56342,17'd56342,17'd67707,17'd57385,17'd67708,17'd67709,17'd55674,17'd58276,17'd60176,17'd58279,17'd61195,17'd67710,17'd59941,17'd67711,17'd60424,17'd55090,17'd65203,17'd5687,17'd67712,17'd67595,17'd67713,17'd67329,17'd67330,17'd66968,17'd67211,17'd67599,17'd67714,17'd67334,17'd66970,17'd67715,17'd67481,17'd67482,17'd67483,17'd67716,17'd62376,17'd67484,17'd67717,17'd67718,17'd67219,17'd66720,17'd67719,17'd66594,17'd67344,17'd67720,17'd67721,17'd67606,17'd12690,17'd67722,17'd55811,17'd15416,17'd67723,17'd67724,17'd35368,17'd67725,17'd67726,17'd16554,17'd18196,17'd10325,17'd10856,17'd67727,17'd67728,17'd67729,17'd16444,17'd8427,17'd67730,17'd67731,17'd67732,17'd13777,17'd11541,17'd20762,17'd20762,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd1481,17'd1481,17'd130,17'd130,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd131,17'd131,17'd132,17'd134,17'd130,17'd132,17'd20622,17'd66251,17'd51716,17'd67733,17'd67734,17'd67735,17'd67736,17'd67737,17'd67738,17'd67739,17'd67740,17'd67741,17'd67742,17'd67743,17'd50641,17'd67744,17'd67745,17'd67746,17'd67747,17'd67748,17'd67748,17'd67749,17'd67749,17'd67750,17'd67751,17'd67752,17'd67380,17'd67753,17'd67753,17'd67381,17'd67380,17'd67754,17'd67380,17'd67755,17'd67756,17'd50557,17'd50557,17'd50557,17'd67250,17'd67629,17'd67629,17'd67629,17'd67520,17'd67520,17'd67520,17'd67520,17'd67629,17'd67251,17'd67757,17'd67009,17'd66628,17'd66274,17'd64466,17'd58329,17'd67256,17'd62656,17'd38978,17'd30126,17'd24744,17'd24898,17'd25178,17'd27511,17'd27882,17'd28717,17'd31367,17'd30904,17'd67758,17'd35731,17'd67759,17'd67760,17'd60607,17'd67761,17'd67762,17'd67763,17'd22197,17'd67764,17'd67765,17'd67639,17'd67766,17'd67767,17'd67768,17'd17381,17'd67769,17'd67770,17'd67771,17'd67772,17'd67773,17'd67774,17'd67775,17'd67776,17'd67777,17'd19587,17'd14710,17'd14710,17'd16112,17'd67778,17'd25480,17'd21451,17'd21141,17'd67779,17'd11159,17'd10361,17'd7170,17'd6847,17'd6215,17'd7667,17'd7999,17'd8629,17'd8154,17'd6390,17'd6853,17'd6853,17'd35760,17'd6224,17'd7011,17'd6557,17'd6854,17'd7837,17'd67780,17'd67781,17'd67782,17'd67783,17'd67784,17'd67785,17'd67786,17'd67549,17'd67787,17'd67788,17'd66180,17'd67551,17'd67037,17'd67286,17'd67037,17'd64089,17'd67789,17'd67790,17'd64628,17'd65552,17'd67791,17'd67792,17'd67050,17'd67170,17'd67793,17'd64110,17'd67667,17'd67794,17'd66677,17'd66677,17'd66072,17'd64919,17'd65702,17'd66197,17'd65830,17'd62699,17'd16381,17'd16381,17'd62575,17'd14735,17'd14735,17'd14735,17'd65947,17'd14176,17'd14176,17'd65947,17'd65947,17'd65947,17'd63653,17'd63653,17'd13571,17'd65946,17'd67795,17'd67796,17'd67293,17'd67431,17'd67431,17'd67293,17'd12318,17'd65946,17'd13056,17'd62445,17'd62444,17'd15735,17'd66070,17'd66194,17'd66193,17'd66193,17'd67044,17'd67046,17'd67797,17'd67797,17'd67433,17'd62847,17'd15862,17'd67798,17'd62445,17'd63653,17'd65947,17'd65565,17'd62447,17'd15618,17'd15618,17'd65571,17'd62851,17'd63375,17'd66073,17'd65703,17'd66677,17'd67799,17'd65305,17'd65305,17'd66073,17'd66073,17'd64530,17'd67671,17'd64529,17'd64241,17'd65831,17'd67439,17'd67672,17'd67674,17'd67560,17'd67800,17'd63246,17'd67801,17'd67802,17'd11187,17'd5771,17'd4551,17'd65940,17'd2723,17'd62704,17'd61674,17'd67803,17'd67804,17'd67805,17'd67564,17'd67806,17'd2230,17'd56109,17'd67807
},
'{
17'd3427,17'd3427,17'd3751,17'd2934,17'd3101,17'd2935,17'd2422,17'd1831,17'd1688,17'd14,17'd466,17'd2595,17'd4247,17'd3252,17'd67808,17'd67809,17'd67183,17'd67810,17'd66555,17'd67568,17'd67687,17'd67688,17'd67811,17'd67812,17'd67813,17'd67813,17'd67814,17'd66559,17'd9674,17'd67815,17'd67816,17'd11885,17'd65189,17'd67817,17'd8194,17'd14187,17'd9422,17'd5969,17'd3748,17'd20404,17'd3905,17'd3905,17'd1416,17'd2257,17'd2597,17'd3752,17'd2422,17'd2934,17'd4087,17'd4734,17'd52928,17'd52928,17'd7049,17'd14744,17'd5203,17'd4086,17'd2934,17'd2593,17'd10669,17'd10669,17'd1130,17'd1130,17'd3103,17'd2262,17'd45516,17'd3103,17'd47968,17'd20405,17'd1558,17'd2948,17'd4741,17'd5808,17'd12337,17'd6279,17'd11345,17'd11737,17'd5976,17'd5976,17'd5975,17'd12657,17'd25903,17'd30949,17'd67818,17'd67819,17'd67820,17'd67821,17'd67822,17'd63832,17'd67823,17'd67824,17'd67825,17'd19139,17'd13610,17'd67826,17'd13481,17'd66952,17'd10698,17'd43467,17'd9845,17'd9843,17'd9705,17'd24522,17'd9441,17'd6138,17'd8073,17'd42795,17'd67587,17'd7095,17'd67466,17'd4463,17'd3954,17'd58644,17'd67827,17'd66347,17'd47973,17'd48299,17'd47972,17'd56343,17'd57013,17'd66107,17'd65733,17'd65082,17'd64000,17'd59789,17'd65081,17'd67828,17'd65735,17'd65734,17'd56901,17'd54614,17'd48932,17'd55576,17'd53810,17'd57123,17'd67829,17'd67830,17'd67707,17'd67830,17'd67831,17'd57385,17'd56901,17'd58151,17'd56581,17'd57278,17'd59274,17'd60180,17'd67832,17'd67833,17'd56460,17'd59796,17'd57273,17'd67834,17'd5082,17'd67835,17'd67836,17'd67837,17'd67329,17'd67838,17'd67600,17'd67839,17'd67840,17'd67841,17'd67334,17'd66970,17'd67601,17'd67337,17'd67338,17'd67842,17'd67716,17'd67843,17'd67484,17'd67603,17'd67604,17'd67844,17'd66720,17'd67719,17'd67845,17'd67845,17'd67345,17'd67846,17'd67847,17'd15161,17'd67848,17'd11108,17'd67849,17'd67850,17'd30213,17'd35368,17'd67851,17'd9608,17'd18194,17'd15048,17'd26034,17'd9341,17'd67852,17'd67853,17'd67854,17'd26040,17'd14266,17'd67855,17'd67856,17'd67857,17'd17363,17'd134,17'd141,17'd67858,17'd130,17'd132,17'd130,17'd130,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd1481,17'd1481,17'd130,17'd130,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd130,17'd130,17'd130,17'd130,17'd132,17'd134,17'd11541,17'd131,17'd132,17'd134,17'd128,17'd132,17'd133,17'd21375,17'd67859,17'd67860,17'd67861,17'd67862,17'd67863,17'd67864,17'd67737,17'd67865,17'd67866,17'd67867,17'd67868,17'd67869,17'd67870,17'd67870,17'd67871,17'd67872,17'd67873,17'd67873,17'd67874,17'd67875,17'd67876,17'd67877,17'd67877,17'd67248,17'd67878,17'd67879,17'd67880,17'd67755,17'd67881,17'd67882,17'd67882,17'd67882,17'd50557,17'd67883,17'd67883,17'd67883,17'd67884,17'd67885,17'd67885,17'd67886,17'd67886,17'd67886,17'd67521,17'd67520,17'd67629,17'd67630,17'd67887,17'd60356,17'd66274,17'd67888,17'd67889,17'd65138,17'd62797,17'd38978,17'd29688,17'd28718,17'd28595,17'd27637,17'd29103,17'd25438,17'd33484,17'd25568,17'd31521,17'd67890,17'd67891,17'd26071,17'd67892,17'd67893,17'd67635,17'd67894,17'd67895,17'd67896,17'd66517,17'd67897,17'd67898,17'd67899,17'd67900,17'd67272,17'd67901,17'd67902,17'd67769,17'd67903,17'd67904,17'd67271,17'd18478,17'd67905,17'd67906,17'd9074,17'd67907,17'd15846,17'd14561,17'd14846,17'd15211,17'd16474,17'd25480,17'd25480,17'd14295,17'd17268,17'd67908,17'd9068,17'd6847,17'd6216,17'd7176,17'd7999,17'd8629,17'd9090,17'd6220,17'd6219,17'd6853,17'd6223,17'd35760,17'd7011,17'd6558,17'd6709,17'd6854,17'd67909,17'd67910,17'd67911,17'd67912,17'd67913,17'd67914,17'd67915,17'd67916,17'd67549,17'd67664,17'd67917,17'd66180,17'd67551,17'd63940,17'd64226,17'd67037,17'd64089,17'd67789,17'd64902,17'd64902,17'd67918,17'd67919,17'd63658,17'd67920,17'd67921,17'd64110,17'd67050,17'd67667,17'd67922,17'd67923,17'd66677,17'd66072,17'd64919,17'd64919,17'd67924,17'd66197,17'd65830,17'd65701,17'd62699,17'd62698,17'd67925,17'd67926,17'd67925,17'd67927,17'd67928,17'd67929,17'd67929,17'd67927,17'd67927,17'd65947,17'd65565,17'd65946,17'd67795,17'd62199,17'd67795,17'd12175,17'd12175,17'd12175,17'd67930,17'd65946,17'd66071,17'd62445,17'd67925,17'd62574,17'd63961,17'd66070,17'd66926,17'd67044,17'd67044,17'd67046,17'd63105,17'd67797,17'd67797,17'd67433,17'd17180,17'd62574,17'd62445,17'd64918,17'd65947,17'd65947,17'd65565,17'd62447,17'd67426,17'd17179,17'd65441,17'd63375,17'd63244,17'd65570,17'd65703,17'd67423,17'd65569,17'd65569,17'd65305,17'd66073,17'd66676,17'd67671,17'd64112,17'd64922,17'd65307,17'd67296,17'd67931,17'd67672,17'd67674,17'd66075,17'd67932,17'd63109,17'd66549,17'd65572,17'd67933,17'd5771,17'd46698,17'd67934,17'd67935,17'd53870,17'd61674,17'd61161,17'd21942,17'd53515,17'd60033,17'd67936,17'd56109,17'd2383,17'd67937
},
'{
17'd3901,17'd3901,17'd2934,17'd2934,17'd2935,17'd3252,17'd2258,17'd2258,17'd1415,17'd1414,17'd1414,17'd1415,17'd1688,17'd10535,17'd2592,17'd67444,17'd65581,17'd67938,17'd67939,17'd66809,17'd67940,17'd67941,17'd67447,17'd67942,17'd67943,17'd67944,17'd67945,17'd67573,17'd67946,17'd9265,17'd65717,17'd67815,17'd64254,17'd65067,17'd9683,17'd8669,17'd14319,17'd12,17'd808,17'd1128,17'd1128,17'd3905,17'd17,17'd1414,17'd2597,17'd2597,17'd2258,17'd2935,17'd3751,17'd5511,17'd52778,17'd67947,17'd14744,17'd15117,17'd6730,17'd4086,17'd10925,17'd10802,17'd52621,17'd3429,17'd32,17'd32,17'd656,17'd656,17'd3253,17'd2262,17'd1973,17'd1702,17'd1702,17'd2431,17'd25902,17'd4741,17'd12786,17'd5977,17'd6111,17'd6111,17'd11345,17'd6279,17'd11737,17'd5975,17'd4898,17'd30811,17'd67948,17'd67949,17'd67950,17'd67951,17'd67952,17'd67953,17'd67954,17'd67955,17'd67956,17'd67957,17'd21655,17'd67826,17'd67958,17'd12820,17'd67959,17'd13098,17'd12068,17'd10121,17'd9843,17'd9578,17'd29181,17'd65975,17'd9985,17'd8072,17'd8070,17'd7421,17'd7095,17'd7090,17'd3950,17'd59265,17'd65858,17'd14624,17'd47974,17'd47973,17'd52932,17'd56343,17'd56232,17'd53810,17'd58272,17'd54172,17'd65733,17'd54993,17'd56021,17'd54701,17'd54615,17'd65469,17'd56804,17'd65603,17'd58272,17'd67960,17'd67960,17'd53880,17'd57265,17'd55374,17'd67830,17'd56342,17'd34177,17'd67961,17'd57636,17'd54021,17'd54705,17'd56351,17'd57516,17'd58893,17'd57778,17'd67962,17'd60426,17'd60052,17'd55580,17'd67963,17'd62223,17'd67964,17'd67965,17'd67966,17'd67093,17'd67967,17'd67968,17'd67969,17'd67970,17'd67971,17'd67972,17'd67601,17'd67973,17'd67974,17'd67975,17'd67976,17'd67340,17'd63302,17'd67484,17'd67977,17'd67978,17'd67979,17'd67980,17'd67845,17'd67981,17'd67845,17'd67982,17'd67983,17'd67984,17'd15034,17'd11373,17'd15284,17'd67985,17'd67986,17'd31757,17'd9330,17'd67987,17'd50411,17'd9337,17'd9479,17'd33722,17'd27856,17'd15430,17'd67988,17'd16918,17'd10610,17'd13378,17'd67989,17'd67990,17'd67991,17'd7980,17'd132,17'd130,17'd130,17'd130,17'd128,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd20623,17'd67992,17'd67993,17'd67994,17'd67995,17'd67996,17'd67997,17'd67998,17'd67999,17'd68000,17'd68001,17'd68002,17'd68003,17'd68004,17'd68005,17'd68006,17'd68007,17'd68008,17'd68009,17'd68009,17'd68006,17'd68010,17'd68011,17'd68011,17'd68012,17'd68013,17'd68014,17'd68014,17'd68015,17'd68015,17'd68016,17'd68016,17'd68017,17'd68017,17'd68018,17'd68019,17'd68020,17'd68020,17'd68021,17'd68022,17'd68023,17'd68024,17'd68025,17'd68026,17'd67251,17'd50558,17'd68027,17'd68028,17'd68029,17'd58464,17'd65377,17'd58823,17'd57839,17'd33317,17'd30446,17'd68030,17'd37387,17'd25318,17'd25320,17'd28254,17'd24411,17'd24898,17'd33968,17'd31057,17'd68031,17'd22700,17'd68032,17'd60863,17'd68033,17'd24621,17'd68034,17'd68035,17'd68036,17'd68037,17'd68038,17'd68039,17'd68040,17'd68041,17'd68042,17'd68043,17'd68044,17'd68045,17'd68041,17'd67271,17'd68046,17'd67541,17'd68047,17'd11425,17'd16472,17'd12604,17'd14710,17'd16238,17'd15212,17'd25617,17'd68048,17'd24940,17'd16601,17'd11160,17'd9220,17'd8146,17'd6550,17'd7176,17'd6704,17'd6553,17'd8154,17'd7668,17'd7668,17'd7177,17'd6393,17'd6393,17'd67151,17'd11039,17'd6854,17'd7013,17'd6855,17'd68049,17'd68050,17'd68051,17'd68052,17'd68053,17'd68054,17'd68055,17'd67662,17'd67420,17'd65930,17'd67286,17'd68056,17'd64368,17'd67286,17'd63940,17'd67790,17'd67790,17'd68057,17'd66062,17'd68058,17'd67919,17'd67932,17'd65306,17'd67170,17'd67050,17'd67050,17'd67553,17'd67923,17'd68059,17'd68059,17'd68060,17'd66318,17'd66319,17'd68061,17'd64387,17'd64387,17'd63962,17'd63106,17'd62848,17'd65949,17'd62698,17'd15999,17'd15232,17'd65829,17'd68062,17'd17785,17'd17785,17'd17785,17'd67927,17'd13571,17'd13055,17'd67930,17'd67930,17'd67930,17'd67930,17'd67669,17'd65946,17'd12772,17'd12772,17'd13056,17'd65304,17'd62444,17'd64649,17'd15735,17'd63104,17'd67047,17'd67046,17'd67046,17'd64386,17'd64526,17'd64386,17'd67433,17'd63371,17'd17180,17'd16381,17'd64918,17'd65946,17'd12772,17'd68063,17'd67291,17'd14434,17'd67557,17'd67426,17'd62971,17'd68064,17'd68065,17'd64527,17'd65703,17'd64529,17'd65570,17'd66072,17'd66072,17'd65054,17'd65305,17'd65703,17'd64654,17'd63657,17'd64388,17'd67295,17'd67296,17'd67438,17'd67931,17'd67296,17'd63809,17'd66321,17'd68066,17'd66679,17'd68067,17'd68068,17'd8011,17'd4051,17'd68069,17'd68070,17'd53291,17'd41312,17'd68071,17'd67058,17'd63650,17'd60149,17'd68072,17'd68073,17'd68074,17'd1085
},
'{
17'd3901,17'd3901,17'd2934,17'd2934,17'd2935,17'd2784,17'd3429,17'd2258,17'd1414,17'd1414,17'd2596,17'd2936,17'd1688,17'd10535,17'd3250,17'd68075,17'd64396,17'd65844,17'd66554,17'd66809,17'd67940,17'd68076,17'd68077,17'd68078,17'd68079,17'd68080,17'd68081,17'd67304,17'd66691,17'd65960,17'd66087,17'd68082,17'd65583,17'd64122,17'd64799,17'd8194,17'd68083,17'd1,17'd3748,17'd11,17'd1128,17'd18,17'd17,17'd1416,17'd1414,17'd2597,17'd2258,17'd52621,17'd2593,17'd15496,17'd53228,17'd52778,17'd7049,17'd14744,17'd5203,17'd4086,17'd10925,17'd10802,17'd52621,17'd3429,17'd32,17'd32,17'd33,17'd33,17'd3253,17'd3253,17'd2785,17'd1973,17'd1702,17'd1974,17'd25902,17'd5805,17'd12786,17'd12337,17'd6111,17'd6112,17'd11345,17'd6279,17'd11737,17'd5975,17'd12787,17'd4093,17'd34513,17'd68084,17'd68085,17'd68086,17'd63395,17'd68087,17'd68088,17'd68089,17'd68090,17'd68091,17'd67704,17'd13610,17'd67958,17'd68092,17'd68093,17'd68094,17'd11235,17'd10566,17'd10121,17'd9579,17'd9578,17'd29181,17'd68095,17'd9985,17'd8073,17'd8070,17'd7097,17'd6934,17'd7090,17'd52625,17'd58517,17'd58269,17'd48300,17'd68096,17'd59012,17'd57012,17'd56343,17'd55483,17'd53950,17'd58272,17'd54172,17'd56446,17'd55185,17'd60171,17'd64682,17'd68097,17'd67195,17'd56804,17'd56446,17'd57773,17'd66349,17'd54020,17'd53810,17'd57123,17'd54797,17'd56342,17'd34177,17'd34937,17'd49814,17'd55483,17'd54171,17'd56021,17'd68098,17'd58653,17'd62232,17'd58888,17'd59647,17'd62105,17'd59016,17'd64143,17'd68099,17'd68100,17'd67965,17'd67966,17'd67093,17'd67967,17'd68101,17'd68102,17'd68103,17'd67971,17'd68104,17'd67601,17'd67973,17'd68105,17'd68106,17'd68107,17'd68108,17'd63302,17'd62132,17'd68109,17'd68110,17'd68111,17'd68112,17'd67845,17'd67981,17'd67845,17'd68113,17'd67983,17'd68114,17'd68115,17'd68116,17'd68117,17'd68118,17'd68119,17'd68120,17'd9330,17'd68121,17'd68122,17'd24039,17'd10334,17'd24998,17'd9344,17'd16318,17'd28963,17'd12726,17'd58078,17'd13378,17'd68123,17'd68124,17'd10757,17'd7980,17'd131,17'd132,17'd131,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd134,17'd20623,17'd65635,17'd21682,17'd51822,17'd68125,17'd68126,17'd68127,17'd68128,17'd68129,17'd68130,17'd67869,17'd68131,17'd68132,17'd68006,17'd68133,17'd68134,17'd68135,17'd68136,17'd68137,17'd68138,17'd68016,17'd67883,17'd67883,17'd68139,17'd68140,17'd68141,17'd68141,17'd68140,17'd68140,17'd68142,17'd68142,17'd68143,17'd68020,17'd68020,17'd68144,17'd68145,17'd68146,17'd68146,17'd68147,17'd68148,17'd68025,17'd68149,17'd67252,17'd50558,17'd60356,17'd58330,17'd62022,17'd64730,17'd58583,17'd51307,17'd56285,17'd56966,17'd32659,17'd68030,17'd68150,17'd68151,17'd31521,17'd28254,17'd28254,17'd23559,17'd31512,17'd25711,17'd30607,17'd68152,17'd31059,17'd68153,17'd68154,17'd68155,17'd68156,17'd68157,17'd66643,17'd68158,17'd68159,17'd68160,17'd68161,17'd68162,17'd67904,17'd68163,17'd68164,17'd68165,17'd68166,17'd67536,17'd68167,17'd67276,17'd68168,17'd68169,17'd18720,17'd9767,17'd15329,17'd14846,17'd17511,17'd15213,17'd68170,17'd66655,17'd25876,17'd14417,17'd11423,17'd68171,17'd6849,17'd68172,17'd7176,17'd7999,17'd8303,17'd7499,17'd8780,17'd10380,17'd10238,17'd6558,17'd6557,17'd57866,17'd11039,17'd7012,17'd68173,17'd7013,17'd68174,17'd68175,17'd68176,17'd68177,17'd68178,17'd68179,17'd68180,17'd67419,17'd65683,17'd65930,17'd67286,17'd68056,17'd67286,17'd64226,17'd63940,17'd67552,17'd67790,17'd68057,17'd66062,17'd67791,17'd68181,17'd63657,17'd65306,17'd67170,17'd67050,17'd67921,17'd67922,17'd68059,17'd68059,17'd68182,17'd68182,17'd66318,17'd66319,17'd66319,17'd68061,17'd64387,17'd63807,17'd63106,17'd63372,17'd66927,17'd66196,17'd15483,17'd15483,17'd65829,17'd16381,17'd17785,17'd67927,17'd65947,17'd65565,17'd13055,17'd18033,17'd18033,17'd18033,17'd18033,17'd13055,17'd12772,17'd12772,17'd12772,17'd12772,17'd65304,17'd65304,17'd62574,17'd15862,17'd62847,17'd67433,17'd67044,17'd67044,17'd63105,17'd64386,17'd64386,17'd63106,17'd68183,17'd65949,17'd16381,17'd67927,17'd62331,17'd65946,17'd13055,17'd68063,17'd67291,17'd14583,17'd67426,17'd62700,17'd68184,17'd68185,17'd68186,17'd67793,17'd65703,17'd65703,17'd66676,17'd66073,17'd66072,17'd66072,17'd65570,17'd63965,17'd63657,17'd64111,17'd67172,17'd66320,17'd68187,17'd68187,17'd67296,17'd65055,17'd64528,17'd65286,17'd62701,17'd66200,17'd68188,17'd68068,17'd9529,17'd4051,17'd68189,17'd3211,17'd55165,17'd40407,17'd61162,17'd63958,17'd66081,17'd60033,17'd56552,17'd60146,17'd68190,17'd25894
},
'{
17'd3901,17'd3901,17'd2934,17'd2934,17'd2935,17'd2422,17'd2258,17'd2258,17'd1414,17'd1414,17'd1414,17'd1415,17'd1688,17'd10535,17'd1831,17'd68191,17'd65312,17'd67683,17'd66554,17'd66329,17'd68192,17'd68076,17'd68193,17'd68194,17'd68195,17'd68080,17'd68196,17'd68197,17'd68198,17'd68199,17'd66086,17'd68200,17'd8043,17'd64397,17'd63821,17'd8341,17'd67452,17'd1412,17'd979,17'd10,17'd11,17'd1128,17'd3905,17'd1416,17'd1414,17'd2257,17'd2258,17'd3429,17'd2784,17'd3901,17'd52704,17'd66816,17'd7049,17'd14744,17'd5203,17'd5204,17'd11888,17'd10670,17'd52621,17'd52621,17'd982,17'd2259,17'd32,17'd32,17'd16866,17'd3253,17'd2263,17'd2785,17'd19874,17'd1974,17'd25902,17'd5805,17'd5808,17'd5977,17'd30948,17'd6112,17'd10672,17'd11345,17'd11737,17'd67454,17'd12200,17'd5057,17'd68201,17'd68202,17'd68203,17'd68204,17'd62347,17'd68087,17'd68205,17'd64415,17'd67466,17'd67824,17'd68206,17'd11236,17'd68207,17'd68208,17'd13336,17'd13608,17'd12366,17'd10948,17'd9988,17'd9705,17'd9705,17'd10118,17'd30059,17'd68095,17'd63834,17'd64813,17'd8376,17'd43069,17'd7090,17'd3784,17'd59512,17'd58517,17'd58759,17'd52933,17'd64817,17'd58027,17'd57120,17'd56232,17'd55483,17'd48931,17'd58272,17'd54172,17'd54894,17'd54804,17'd65735,17'd68209,17'd67317,17'd57014,17'd57126,17'd65733,17'd64820,17'd48932,17'd57504,17'd49303,17'd54797,17'd54797,17'd54797,17'd49814,17'd49814,17'd55483,17'd48931,17'd65733,17'd60170,17'd56694,17'd56239,17'd58524,17'd59933,17'd58036,17'd55580,17'd64145,17'd68210,17'd68211,17'd68212,17'd68213,17'd67093,17'd67096,17'd68214,17'd67970,17'd68215,17'd68216,17'd68217,17'd68104,17'd67334,17'd68105,17'd68106,17'd67976,17'd67340,17'd67843,17'd68218,17'd68219,17'd68220,17'd68221,17'd66847,17'd67845,17'd66594,17'd67845,17'd68113,17'd67983,17'd68222,17'd68223,17'd56722,17'd54641,17'd68224,17'd30825,17'd68225,17'd68226,17'd68227,17'd68228,17'd9193,17'd15807,17'd19279,17'd9346,17'd24039,17'd28963,17'd54046,17'd24864,17'd13378,17'd68123,17'd68229,17'd68230,17'd68231,17'd131,17'd135,17'd135,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd21834,17'd51624,17'd68232,17'd68233,17'd68234,17'd68235,17'd68236,17'd67364,17'd68237,17'd68238,17'd68239,17'd68240,17'd68241,17'd68138,17'd68242,17'd68243,17'd68244,17'd68245,17'd68246,17'd68021,17'd68020,17'd68247,17'd68248,17'd68249,17'd68249,17'd68249,17'd68250,17'd68251,17'd68021,17'd68145,17'd68146,17'd68252,17'd68253,17'd68253,17'd68254,17'd68254,17'd68255,17'd68256,17'd68257,17'd68149,17'd67253,17'd67130,17'd66506,17'd64189,17'd65003,17'd64870,17'd58207,17'd50464,17'd62797,17'd53405,17'd30431,17'd28601,17'd27763,17'd28596,17'd31521,17'd68258,17'd28596,17'd25029,17'd24898,17'd33666,17'd68259,17'd60603,17'd68260,17'd68261,17'd68262,17'd68263,17'd68264,17'd68265,17'd68266,17'd68267,17'd68268,17'd68269,17'd68270,17'd68271,17'd67770,17'd68166,17'd68272,17'd68273,17'd68274,17'd68275,17'd17633,17'd68276,17'd68277,17'd9377,17'd68278,17'd18720,17'd9767,17'd14415,17'd14293,17'd68279,17'd15715,17'd68280,17'd25478,17'd68281,17'd16600,17'd11551,17'd8292,17'd6386,17'd6850,17'd6705,17'd6553,17'd8154,17'd7668,17'd27815,17'd10516,17'd9934,17'd6557,17'd8471,17'd11039,17'd10517,17'd29299,17'd29163,17'd68282,17'd68283,17'd68284,17'd68285,17'd68286,17'd68287,17'd68179,17'd68288,17'd67549,17'd68289,17'd67286,17'd64368,17'd67286,17'd67286,17'd64628,17'd67790,17'd67790,17'd67790,17'd66062,17'd65815,17'd68290,17'd68291,17'd64654,17'd64529,17'd67423,17'd68292,17'd68293,17'd67922,17'd68059,17'd68182,17'd68182,17'd68182,17'd66318,17'd66319,17'd66319,17'd66319,17'd64387,17'd63807,17'd66197,17'd65950,17'd65701,17'd65701,17'd16959,17'd16959,17'd15232,17'd15232,17'd15232,17'd66434,17'd65565,17'd13932,17'd66071,17'd66071,17'd13932,17'd13932,17'd65565,17'd65947,17'd65947,17'd65565,17'd65304,17'd62445,17'd14584,17'd14584,17'd15862,17'd68294,17'd67433,17'd67797,17'd64386,17'd64386,17'd63105,17'd63105,17'd68295,17'd68295,17'd68296,17'd65829,17'd63653,17'd65565,17'd62331,17'd67430,17'd13055,17'd68063,17'd67291,17'd67557,17'd17179,17'd62853,17'd68064,17'd68065,17'd68297,17'd64110,17'd65703,17'd65570,17'd66073,17'd66073,17'd66072,17'd66437,17'd65570,17'd65703,17'd64110,17'd63657,17'd66075,17'd67674,17'd68298,17'd68187,17'd66320,17'd63657,17'd68299,17'd66790,17'd14976,17'd66438,17'd68300,17'd67175,17'd8480,17'd68301,17'd68302,17'd3061,17'd39027,17'd56324,17'd61282,17'd52770,17'd53145,17'd35904,17'd58002,17'd58494,17'd68303,17'd51582
},
'{
17'd3901,17'd3901,17'd2934,17'd2934,17'd2935,17'd2422,17'd2258,17'd2258,17'd2257,17'd2257,17'd1414,17'd1415,17'd1689,17'd1831,17'd1831,17'd2592,17'd65187,17'd67062,17'd68304,17'd66686,17'd68192,17'd67569,17'd68305,17'd68306,17'd68307,17'd68308,17'd68309,17'd68310,17'd68311,17'd68312,17'd68304,17'd68313,17'd8515,17'd67305,17'd63979,17'd8983,17'd63521,17'd4884,17'd19,17'd10,17'd11,17'd1128,17'd3905,17'd17,17'd1416,17'd1414,17'd2597,17'd3429,17'd2592,17'd2934,17'd15877,17'd53228,17'd66816,17'd14744,17'd5203,17'd5204,17'd16501,17'd10925,17'd10802,17'd52621,17'd982,17'd982,17'd292,17'd292,17'd16866,17'd16866,17'd2602,17'd2263,17'd1974,17'd1975,17'd25902,17'd5805,17'd5808,17'd12337,17'd6280,17'd6112,17'd10672,17'd10672,17'd11345,17'd11737,17'd67454,17'd68314,17'd13189,17'd68315,17'd68316,17'd68317,17'd62588,17'd68318,17'd68319,17'd68320,17'd68321,17'd67080,17'd65744,17'd41497,17'd11482,17'd68322,17'd13336,17'd13479,17'd13729,17'd11917,17'd11092,17'd10566,17'd9844,17'd10119,17'd10118,17'd29181,17'd66105,17'd63834,17'd8073,17'd8376,17'd7258,17'd7090,17'd4123,17'd52782,17'd52471,17'd52471,17'd53018,17'd53081,17'd53163,17'd56343,17'd55483,17'd55483,17'd53810,17'd66107,17'd65981,17'd54706,17'd55900,17'd57014,17'd68323,17'd64823,17'd64419,17'd55185,17'd68324,17'd65738,17'd54251,17'd68325,17'd48641,17'd55373,17'd55373,17'd55374,17'd56232,17'd56232,17'd55483,17'd66107,17'd64552,17'd68326,17'd55489,17'd56909,17'd57915,17'd63279,17'd68327,17'd56351,17'd68328,17'd68329,17'd68330,17'd68331,17'd68332,17'd67096,17'd67714,17'd68333,17'd68334,17'd68216,17'd68217,17'd68335,17'd67334,17'd68336,17'd68337,17'd68338,17'd68339,17'd68340,17'd68218,17'd68341,17'd68110,17'd68342,17'd68343,17'd67845,17'd66594,17'd67845,17'd68113,17'd67983,17'd68222,17'd15033,17'd68344,17'd68345,17'd68346,17'd68347,17'd68348,17'd9463,17'd68349,17'd68228,17'd16318,17'd14674,17'd19279,17'd9346,17'd11529,17'd68350,17'd22133,17'd24716,17'd24552,17'd68123,17'd68351,17'd9358,17'd68231,17'd131,17'd135,17'd135,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd134,17'd131,17'd21375,17'd68352,17'd68353,17'd68354,17'd68355,17'd68356,17'd68357,17'd68358,17'd50891,17'd68359,17'd68360,17'd68361,17'd68362,17'd68363,17'd68242,17'd68364,17'd68365,17'd68366,17'd68367,17'd68368,17'd68369,17'd68369,17'd68370,17'd68371,17'd68372,17'd68372,17'd68373,17'd68374,17'd68375,17'd68375,17'd68376,17'd68377,17'd68378,17'd68379,17'd68380,17'd68381,17'd68382,17'd68383,17'd61891,17'd67385,17'd60475,17'd62784,17'd67131,17'd50728,17'd56391,17'd50650,17'd50464,17'd57205,17'd53405,17'd29534,17'd24743,17'd34622,17'd28595,17'd25029,17'd31521,17'd68151,17'd24896,17'd24896,17'd24417,17'd68384,17'd68385,17'd68386,17'd68387,17'd66637,17'd68388,17'd68389,17'd68390,17'd68391,17'd68035,17'd68392,17'd68393,17'd67533,17'd68394,17'd67903,17'd68166,17'd68395,17'd68273,17'd68396,17'd68397,17'd68398,17'd17748,17'd18479,17'd68168,17'd68399,17'd68278,17'd18720,17'd9767,17'd15328,17'd14845,17'd19843,17'd15842,17'd68400,17'd68401,17'd16479,17'd15086,17'd9221,17'd7663,17'd11849,17'd6850,17'd8000,17'd6707,17'd8154,17'd8780,17'd10515,17'd10778,17'd10380,17'd10517,17'd10779,17'd8001,17'd7012,17'd29026,17'd68402,17'd29300,17'd68403,17'd68404,17'd68285,17'd68405,17'd68406,17'd68407,17'd68408,17'd68409,17'd65163,17'd64902,17'd66180,17'd67286,17'd67286,17'd64628,17'd67790,17'd67790,17'd68057,17'd65038,17'd65815,17'd68290,17'd64528,17'd64529,17'd64529,17'd67423,17'd68292,17'd68293,17'd67922,17'd68059,17'd68059,17'd68182,17'd68182,17'd66318,17'd66319,17'd66319,17'd68061,17'd63807,17'd63807,17'd66197,17'd65950,17'd65830,17'd65701,17'd16959,17'd16959,17'd15232,17'd15232,17'd15232,17'd66434,17'd13932,17'd66071,17'd13932,17'd13932,17'd65565,17'd65565,17'd65947,17'd65947,17'd65947,17'd63653,17'd63653,17'd63653,17'd68410,17'd15862,17'd17180,17'd68183,17'd68411,17'd67797,17'd63105,17'd63105,17'd64386,17'd63372,17'd68183,17'd65701,17'd68412,17'd16381,17'd65565,17'd66071,17'd68413,17'd67430,17'd68063,17'd67291,17'd14434,17'd15618,17'd62853,17'd62974,17'd63108,17'd64527,17'd64110,17'd64110,17'd65570,17'd65305,17'd66073,17'd66073,17'd66437,17'd66437,17'd65703,17'd65306,17'd63657,17'd64388,17'd66076,17'd68414,17'd68298,17'd67439,17'd65055,17'd68415,17'd65286,17'd68416,17'd62702,17'd66438,17'd66079,17'd68417,17'd5772,17'd3381,17'd68418,17'd52613,17'd2546,17'd52275,17'd2379,17'd68419,17'd52840,17'd68420,17'd56327,17'd68421,17'd18632,17'd36907
},
'{
17'd3901,17'd3901,17'd3427,17'd2934,17'd2935,17'd2422,17'd2258,17'd2258,17'd2257,17'd2257,17'd1127,17'd14,17'd1689,17'd1831,17'd1831,17'd2784,17'd65311,17'd68422,17'd66692,17'd66686,17'd68192,17'd67569,17'd67303,17'd66813,17'd68423,17'd68424,17'd68309,17'd68425,17'd68426,17'd68427,17'd66207,17'd66692,17'd8512,17'd12191,17'd13576,17'd10403,17'd6102,17'd14319,17'd18,17'd10,17'd20,17'd11,17'd1128,17'd3905,17'd17,17'd1414,17'd2597,17'd3752,17'd2592,17'd2593,17'd3592,17'd52704,17'd66816,17'd15359,17'd6730,17'd5204,17'd3592,17'd3427,17'd10802,17'd10669,17'd982,17'd982,17'd982,17'd469,17'd2940,17'd2940,17'd2943,17'd2602,17'd2265,17'd2946,17'd4894,17'd5055,17'd12507,17'd27445,17'd27592,17'd10672,17'd7730,17'd7730,17'd11345,17'd11345,17'd11737,17'd5974,17'd66336,17'd68428,17'd68429,17'd68430,17'd65194,17'd64408,17'd68431,17'd68432,17'd66456,17'd46489,17'd68433,17'd68434,17'd10122,17'd13481,17'd13337,17'd13336,17'd13337,17'd13479,17'd66952,17'd11235,17'd10947,17'd9844,17'd9705,17'd10118,17'd29181,17'd68435,17'd68436,17'd8073,17'd8691,17'd68437,17'd4124,17'd52625,17'd68438,17'd68438,17'd53082,17'd64817,17'd58027,17'd56686,17'd53080,17'd56232,17'd56232,17'd53950,17'd66107,17'd67588,17'd54172,17'd54347,17'd54529,17'd68439,17'd68440,17'd55280,17'd68441,17'd68442,17'd68443,17'd68444,17'd48819,17'd53080,17'd57123,17'd57265,17'd57385,17'd57636,17'd49303,17'd56125,17'd54021,17'd65082,17'd56235,17'd55782,17'd58159,17'd58402,17'd68445,17'd54799,17'd3943,17'd68446,17'd68330,17'd68447,17'd68448,17'd68449,17'd67841,17'd68333,17'd68334,17'd68450,17'd68451,17'd68335,17'd67213,17'd68452,17'd67975,17'd67976,17'd67340,17'd68340,17'd68453,17'd68454,17'd68455,17'd68342,17'd68343,17'd68113,17'd68456,17'd67982,17'd67845,17'd68457,17'd68458,17'd68459,17'd68460,17'd16191,17'd68346,17'd68461,17'd68462,17'd68463,17'd68464,17'd68465,17'd26626,17'd14674,17'd16549,17'd9344,17'd9044,17'd57818,17'd54378,17'd14938,17'd10482,17'd67855,17'd68466,17'd52139,17'd68231,17'd131,17'd132,17'd135,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd720,17'd130,17'd132,17'd134,17'd133,17'd20623,17'd68467,17'd68468,17'd68469,17'd68470,17'd68471,17'd68472,17'd68473,17'd68474,17'd68475,17'd68476,17'd50724,17'd68008,17'd68243,17'd68365,17'd68477,17'd68365,17'd68478,17'd68479,17'd68372,17'd68480,17'd68481,17'd68481,17'd68482,17'd68483,17'd50456,17'd68484,17'd50456,17'd50456,17'd50456,17'd68378,17'd68378,17'd68380,17'd68382,17'd68257,17'd68149,17'd67252,17'd67254,17'd67632,17'd66630,17'd67131,17'd58461,17'd59582,17'd50650,17'd50648,17'd62797,17'd56966,17'd29375,17'd23917,17'd28601,17'd29240,17'd24896,17'd24897,17'd24898,17'd24898,17'd24745,17'd24252,17'd29100,17'd68485,17'd68486,17'd68487,17'd68488,17'd68489,17'd68490,17'd68491,17'd68492,17'd68493,17'd68494,17'd68495,17'd68496,17'd68497,17'd68498,17'd68499,17'd68500,17'd68501,17'd68502,17'd68503,17'd68504,17'd68505,17'd17628,17'd68506,17'd9509,17'd9378,17'd12608,17'd11694,17'd16472,17'd14846,17'd68507,17'd68508,17'd17773,17'd68400,17'd68509,17'd14295,17'd14161,17'd8292,17'd6849,17'd11849,17'd10512,17'd8000,17'd6707,17'd9090,17'd28184,17'd10515,17'd68510,17'd10778,17'd10779,17'd12625,17'd10517,17'd68511,17'd68512,17'd68513,17'd68514,17'd68403,17'd68404,17'd67912,17'd68515,17'd68406,17'd68055,17'd68516,17'd67787,17'd64628,17'd67286,17'd66180,17'd64902,17'd64628,17'd64628,17'd67790,17'd68057,17'd66062,17'd65815,17'd67421,17'd63377,17'd64654,17'd64529,17'd68292,17'd67923,17'd68517,17'd68059,17'd68059,17'd68059,17'd68059,17'd68518,17'd68519,17'd66318,17'd66319,17'd68520,17'd68521,17'd63807,17'd63807,17'd66197,17'd65950,17'd65701,17'd62699,17'd16959,17'd15483,17'd16381,17'd16381,17'd15232,17'd15103,17'd66803,17'd66803,17'd65947,17'd65947,17'd63653,17'd63653,17'd14735,17'd14735,17'd14735,17'd15862,17'd17180,17'd17180,17'd68294,17'd17180,17'd67169,17'd67797,17'd68411,17'd63105,17'd63241,17'd63241,17'd63106,17'd63372,17'd62848,17'd62699,17'd65829,17'd15103,17'd13932,17'd62331,17'd68413,17'd13419,17'd67291,17'd14434,17'd68522,17'd62448,17'd65441,17'd66078,17'd63244,17'd64109,17'd64110,17'd64110,17'd65570,17'd65305,17'd66073,17'd66073,17'd66437,17'd66804,17'd64529,17'd67050,17'd65306,17'd64921,17'd67674,17'd67672,17'd67673,17'd67674,17'd66075,17'd67792,17'd66790,17'd67038,17'd62855,17'd18628,17'd68523,17'd68417,17'd5772,17'd3562,17'd54875,17'd2894,17'd51852,17'd52191,17'd68524,17'd2386,17'd2553,17'd56666,17'd68525,17'd29036,17'd790,17'd20001
},
'{
17'd3592,17'd3901,17'd3427,17'd2934,17'd2935,17'd3252,17'd2258,17'd2258,17'd2257,17'd2257,17'd1127,17'd14,17'd1967,17'd1688,17'd1831,17'd2784,17'd65186,17'd63976,17'd67179,17'd66554,17'd68192,17'd67303,17'd67569,17'd68526,17'd68527,17'd68528,17'd68529,17'd67944,17'd68530,17'd68311,17'd68531,17'd68304,17'd9675,17'd8344,17'd67574,17'd67306,17'd8194,17'd63669,17'd19,17'd10,17'd21,17'd20,17'd1128,17'd18,17'd17,17'd1416,17'd1414,17'd2597,17'd2422,17'd2935,17'd3427,17'd15877,17'd52704,17'd5203,17'd6730,17'd6730,17'd4086,17'd3901,17'd10924,17'd10669,17'd982,17'd982,17'd469,17'd469,17'd2940,17'd2940,17'd2943,17'd2943,17'd2264,17'd2946,17'd4739,17'd5055,17'd13067,17'd12931,17'd6279,17'd10672,17'd7392,17'd7392,17'd7562,17'd11345,17'd11211,17'd6109,17'd68532,17'd68533,17'd68534,17'd68535,17'd68536,17'd68537,17'd65852,17'd68538,17'd68539,17'd51676,17'd49202,17'd68540,17'd68541,17'd11237,17'd13729,17'd13336,17'd13336,17'd13336,17'd13608,17'd12366,17'd11235,17'd10947,17'd10121,17'd9705,17'd10118,17'd29181,17'd66104,17'd9985,17'd8692,17'd8375,17'd4463,17'd52625,17'd59390,17'd59264,17'd53082,17'd68542,17'd53081,17'd56572,17'd48821,17'd48821,17'd56232,17'd56125,17'd55576,17'd66107,17'd65981,17'd66225,17'd68543,17'd68544,17'd57637,17'd68545,17'd68546,17'd68547,17'd66831,17'd54430,17'd66702,17'd57504,17'd57013,17'd56900,17'd57385,17'd57124,17'd49199,17'd49610,17'd55576,17'd64820,17'd68548,17'd54991,17'd56352,17'd58152,17'd68549,17'd68550,17'd3620,17'd68551,17'd68552,17'd68553,17'd68554,17'd68555,17'd68556,17'd68557,17'd68334,17'd68450,17'd68451,17'd68558,17'd68336,17'd68559,17'd68560,17'd68561,17'd68562,17'd68563,17'd68564,17'd68565,17'd68566,17'd68567,17'd67844,17'd68113,17'd67982,17'd67982,17'd67982,17'd68568,17'd14499,17'd68569,17'd56482,17'd52123,17'd68570,17'd68571,17'd68572,17'd68573,17'd68122,17'd68574,17'd26626,17'd17716,17'd16065,17'd15187,17'd9044,17'd35797,17'd11279,17'd14938,17'd10748,17'd68575,17'd68576,17'd68577,17'd7813,17'd133,17'd132,17'd135,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd128,17'd130,17'd132,17'd134,17'd356,17'd133,17'd20625,17'd21682,17'd68578,17'd68579,17'd68580,17'd68581,17'd68582,17'd68583,17'd68584,17'd68585,17'd68586,17'd68587,17'd68588,17'd68589,17'd68590,17'd68482,17'd68482,17'd68591,17'd68591,17'd68482,17'd68482,17'd68591,17'd68591,17'd68483,17'd68592,17'd68592,17'd50456,17'd68593,17'd68377,17'd68380,17'd68255,17'd68025,17'd67521,17'd67251,17'd67129,17'd66756,17'd66506,17'd66274,17'd67131,17'd58461,17'd65139,17'd68594,17'd67256,17'd51735,17'd62655,17'd30424,17'd23731,17'd29100,17'd34884,17'd23561,17'd24417,17'd28718,17'd28718,17'd24742,17'd30431,17'd24086,17'd29242,17'd68595,17'd68596,17'd68597,17'd68598,17'd68599,17'd68600,17'd68601,17'd68602,17'd68603,17'd68604,17'd68605,17'd68606,17'd68607,17'd68608,17'd68609,17'd68610,17'd68611,17'd68612,17'd68613,17'd68614,17'd68615,17'd68616,17'd68617,17'd9645,17'd10888,17'd68618,17'd16717,17'd16472,17'd17393,17'd68619,17'd68508,17'd19569,17'd68620,17'd25876,17'd20531,17'd9639,17'd7172,17'd7010,17'd11849,17'd68621,17'd8000,17'd9090,17'd9657,17'd27815,17'd28183,17'd68622,17'd68510,17'd68623,17'd68624,17'd68625,17'd68626,17'd68627,17'd68628,17'd68513,17'd68629,17'd67911,17'd67912,17'd68630,17'd68054,17'd68288,17'd68409,17'd65163,17'd68631,17'd64902,17'd67286,17'd64628,17'd64628,17'd64628,17'd68057,17'd66062,17'd64766,17'd65815,17'd67421,17'd63377,17'd65703,17'd68292,17'd67423,17'd67923,17'd67923,17'd68059,17'd68182,17'd68059,17'd68059,17'd68518,17'd68519,17'd66318,17'd66319,17'd68520,17'd68521,17'd63807,17'd63807,17'd65950,17'd62849,17'd65701,17'd62699,17'd15483,17'd15483,17'd16381,17'd16381,17'd15232,17'd15232,17'd15103,17'd15103,17'd17785,17'd17785,17'd17660,17'd62575,17'd62575,17'd14735,17'd15862,17'd17180,17'd68294,17'd68294,17'd68294,17'd62848,17'd67433,17'd67797,17'd64386,17'd63105,17'd63241,17'd62969,17'd63106,17'd62849,17'd62699,17'd15483,17'd15232,17'd66434,17'd13932,17'd68413,17'd67430,17'd13419,17'd14434,17'd67557,17'd15618,17'd65571,17'd62973,17'd63376,17'd64527,17'd63965,17'd64110,17'd64110,17'd65570,17'd65305,17'd66073,17'd66676,17'd66437,17'd65703,17'd67050,17'd65306,17'd64921,17'd66320,17'd67672,17'd68632,17'd68633,17'd66076,17'd67800,17'd66663,17'd68416,17'd68634,17'd12481,17'd62452,17'd66680,17'd5625,17'd7849,17'd51856,17'd41314,17'd2894,17'd2899,17'd52191,17'd58995,17'd2735,17'd68635,17'd68636,17'd68637,17'd1238,17'd281,17'd620
},
'{
17'd3592,17'd3592,17'd3427,17'd2934,17'd3101,17'd3252,17'd1831,17'd1831,17'd2257,17'd1414,17'd1127,17'd14,17'd1967,17'd1689,17'd1688,17'd2422,17'd66323,17'd64928,17'd67183,17'd68638,17'd66329,17'd68639,17'd68192,17'd66937,17'd66812,17'd68640,17'd68641,17'd68642,17'd68643,17'd68197,17'd68644,17'd66207,17'd65959,17'd9265,17'd68645,17'd13064,17'd6269,17'd6274,17'd1277,17'd10,17'd21,17'd20,17'd1128,17'd1128,17'd3905,17'd17,17'd1414,17'd2597,17'd1831,17'd2422,17'd2593,17'd15496,17'd5511,17'd5511,17'd6730,17'd5204,17'd3592,17'd3427,17'd10802,17'd10669,17'd3429,17'd2258,17'd1129,17'd1129,17'd291,17'd291,17'd2940,17'd2940,17'd2601,17'd2604,17'd4739,17'd5210,17'd13067,17'd12931,17'd27445,17'd11345,17'd7392,17'd7392,17'd7730,17'd10672,17'd11211,17'd68646,17'd66818,17'd68647,17'd68648,17'd68649,17'd68650,17'd68651,17'd68652,17'd68653,17'd68654,17'd68655,17'd53086,17'd68656,17'd8384,17'd68541,17'd68657,17'd13479,17'd68658,17'd13219,17'd68093,17'd13608,17'd11482,17'd10948,17'd68659,17'd68660,17'd9705,17'd10118,17'd10115,17'd68095,17'd6304,17'd5251,17'd44521,17'd4124,17'd4128,17'd4293,17'd68438,17'd53019,17'd58395,17'd52851,17'd57012,17'd49200,17'd48641,17'd49199,17'd48931,17'd58399,17'd54700,17'd68661,17'd54706,17'd54705,17'd64682,17'd68545,17'd68662,17'd65329,17'd56234,17'd68663,17'd54252,17'd55774,17'd58399,17'd65736,17'd65736,17'd57013,17'd57504,17'd55668,17'd48932,17'd58649,17'd68664,17'd68665,17'd58522,17'd56905,17'd65081,17'd68666,17'd52471,17'd68667,17'd68552,17'd68668,17'd68669,17'd68670,17'd68216,17'd68671,17'd68672,17'd68450,17'd68451,17'd68558,17'd68336,17'd68559,17'd68673,17'd68561,17'd68562,17'd68674,17'd68675,17'd68676,17'd68566,17'd68567,17'd67844,17'd68113,17'd68677,17'd67982,17'd67345,17'd68568,17'd68678,17'd13864,17'd68679,17'd10581,17'd27728,17'd68680,17'd68681,17'd68573,17'd68228,17'd68682,17'd15430,17'd24361,17'd15569,17'd18080,17'd8720,17'd35930,17'd54378,17'd14938,17'd10997,17'd68683,17'd68684,17'd11288,17'd8131,17'd133,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd138,17'd130,17'd21375,17'd21835,17'd21224,17'd51896,17'd68685,17'd68686,17'd68687,17'd68688,17'd68689,17'd68690,17'd67741,17'd68691,17'd68240,17'd68692,17'd68368,17'd68376,17'd50456,17'd68693,17'd68694,17'd68694,17'd68695,17'd68695,17'd68375,17'd68696,17'd68380,17'd68380,17'd68254,17'd68147,17'd68148,17'd68025,17'd67521,17'd67383,17'd67129,17'd68697,17'd68698,17'd68699,17'd68700,17'd67888,17'd59581,17'd58329,17'd68701,17'd57196,17'd64202,17'd65006,17'd58459,17'd24087,17'd30879,17'd28722,17'd29100,17'd24090,17'd24901,17'd24901,17'd30879,17'd23732,17'd35877,17'd50988,17'd31836,17'd68702,17'd68703,17'd68704,17'd68705,17'd68706,17'd68389,17'd68707,17'd68708,17'd68709,17'd68710,17'd68711,17'd68497,17'd68712,17'd68713,17'd68714,17'd68715,17'd17157,17'd68716,17'd68717,17'd68718,17'd68719,17'd68720,17'd68721,17'd9770,17'd9071,17'd11694,17'd68722,17'd11017,17'd17393,17'd19586,17'd68723,17'd19682,17'd68620,17'd17894,17'd14296,17'd8610,17'd7174,17'd11848,17'd68621,17'd10236,17'd10236,17'd9090,17'd9657,17'd27815,17'd28057,17'd68622,17'd68724,17'd68725,17'd68726,17'd68727,17'd68728,17'd68729,17'd68730,17'd68731,17'd68284,17'd68732,17'd68733,17'd68734,17'd68735,17'd67662,17'd67787,17'd65163,17'd64902,17'd64368,17'd67286,17'd64628,17'd64628,17'd64628,17'd68057,17'd66062,17'd68736,17'd65164,17'd67422,17'd63377,17'd65703,17'd68292,17'd67923,17'd68059,17'd68059,17'd68059,17'd68182,17'd68518,17'd68518,17'd68518,17'd68519,17'd66318,17'd66319,17'd68520,17'd68520,17'd63106,17'd63106,17'd63106,17'd63372,17'd62699,17'd62699,17'd16959,17'd16959,17'd65949,17'd65949,17'd62698,17'd62698,17'd65829,17'd65829,17'd65829,17'd65829,17'd17180,17'd17180,17'd17180,17'd64788,17'd63961,17'd63961,17'd62847,17'd62847,17'd62847,17'd67433,17'd67797,17'd64386,17'd63241,17'd63241,17'd63372,17'd63372,17'd68183,17'd65701,17'd68412,17'd15348,17'd67927,17'd13688,17'd13419,17'd67430,17'd68737,17'd67289,17'd62449,17'd65705,17'd17179,17'd65441,17'd63510,17'd67440,17'd63965,17'd63965,17'd64110,17'd67793,17'd65570,17'd65305,17'd65570,17'd65703,17'd65703,17'd65703,17'd67050,17'd64241,17'd65055,17'd67558,17'd67672,17'd67672,17'd68738,17'd68739,17'd68740,17'd68741,17'd68742,17'd67173,17'd11865,17'd68743,17'd5625,17'd46595,17'd7849,17'd41000,17'd55362,17'd68744,17'd68745,17'd68746,17'd58995,17'd2235,17'd68747,17'd38457,17'd68748,17'd455,17'd589,17'd68749
},
'{
17'd3592,17'd3592,17'd3901,17'd3427,17'd3101,17'd2935,17'd2422,17'd1831,17'd2257,17'd1414,17'd1127,17'd14,17'd1967,17'd1689,17'd1688,17'd2422,17'd6584,17'd68750,17'd68751,17'd68752,17'd66686,17'd68753,17'd68076,17'd67941,17'd66813,17'd67571,17'd68641,17'd68642,17'd68754,17'd68310,17'd66690,17'd67940,17'd66088,17'd65959,17'd68755,17'd67574,17'd10922,17'd9552,17'd3749,17'd979,17'd10,17'd20,17'd11,17'd1128,17'd18,17'd17,17'd1414,17'd2257,17'd1688,17'd1688,17'd2784,17'd3428,17'd15877,17'd5511,17'd5203,17'd5511,17'd3592,17'd3901,17'd10924,17'd10669,17'd3429,17'd2258,17'd1129,17'd1129,17'd291,17'd291,17'd2941,17'd2940,17'd2601,17'd2601,17'd3105,17'd5210,17'd5657,17'd12507,17'd6110,17'd11345,17'd7392,17'd7392,17'd7392,17'd7730,17'd11211,17'd68756,17'd12037,17'd12338,17'd3440,17'd68757,17'd68758,17'd68759,17'd68760,17'd68761,17'd68762,17'd68763,17'd47094,17'd39647,17'd64810,17'd8384,17'd18666,17'd68657,17'd13217,17'd13219,17'd68764,17'd68093,17'd12366,17'd66699,17'd10949,17'd9988,17'd9705,17'd24198,17'd30059,17'd68435,17'd9303,17'd5088,17'd5687,17'd4125,17'd3955,17'd3632,17'd3632,17'd53019,17'd64817,17'd52851,17'd58030,17'd49200,17'd50191,17'd56125,17'd48931,17'd58272,17'd54700,17'd55484,17'd65981,17'd54894,17'd56020,17'd68097,17'd65739,17'd65331,17'd68765,17'd68766,17'd65202,17'd55900,17'd58649,17'd54614,17'd58521,17'd66107,17'd58272,17'd55774,17'd57772,17'd58150,17'd65471,17'd55185,17'd60170,17'd54617,17'd54895,17'd54434,17'd65466,17'd68667,17'd68767,17'd68668,17'd68669,17'd68670,17'd68450,17'd68671,17'd68672,17'd68450,17'd68451,17'd68558,17'd68336,17'd68559,17'd68673,17'd68561,17'd68768,17'd68769,17'd61211,17'd68676,17'd68770,17'd68771,17'd68772,17'd68773,17'd68774,17'd68775,17'd67345,17'd68568,17'd68678,17'd13741,17'd16783,17'd21198,17'd68776,17'd68777,17'd68778,17'd68779,17'd68465,17'd29325,17'd16441,17'd23859,17'd17716,17'd53547,17'd9041,17'd8575,17'd54378,17'd14938,17'd7625,17'd68780,17'd68781,17'd17360,17'd53402,17'd1045,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd130,17'd136,17'd128,17'd133,17'd68352,17'd22149,17'd68782,17'd68783,17'd68784,17'd68785,17'd68786,17'd68787,17'd68788,17'd68789,17'd68790,17'd68791,17'd67509,17'd68792,17'd68793,17'd68023,17'd68254,17'd68252,17'd68794,17'd68794,17'd68368,17'd68146,17'd68023,17'd68148,17'd68148,17'd68025,17'd68795,17'd67520,17'd67629,17'd67251,17'd67009,17'd66756,17'd68698,17'd68699,17'd68796,17'd63896,17'd68797,17'd64468,17'd68701,17'd51307,17'd52887,17'd65006,17'd68798,17'd29527,17'd31033,17'd30879,17'd30879,17'd29100,17'd30879,17'd44116,17'd45164,17'd23734,17'd35865,17'd46115,17'd46669,17'd40529,17'd68799,17'd68800,17'd68801,17'd68802,17'd68803,17'd68155,17'd68804,17'd68805,17'd68806,17'd68807,17'd68808,17'd68809,17'd68810,17'd68811,17'd68812,17'd68813,17'd68814,17'd68815,17'd68816,17'd17157,17'd16589,17'd68817,17'd9771,17'd11992,17'd11832,17'd8763,17'd68818,17'd11693,17'd17393,17'd68819,17'd68820,17'd25865,17'd68821,17'd16947,17'd14297,17'd10501,17'd7665,17'd68822,17'd68823,17'd11036,17'd9931,17'd9090,17'd10513,17'd27933,17'd68824,17'd68825,17'd68825,17'd68725,17'd68726,17'd68725,17'd68826,17'd68827,17'd68730,17'd68828,17'd68829,17'd68830,17'd68733,17'd68831,17'd68832,17'd67549,17'd67787,17'd68631,17'd64628,17'd64902,17'd67286,17'd64628,17'd64628,17'd64902,17'd66062,17'd64766,17'd68736,17'd67287,17'd67422,17'd63377,17'd65703,17'd68292,17'd67923,17'd67923,17'd68059,17'd68059,17'd68182,17'd68519,17'd68519,17'd68519,17'd68519,17'd66928,17'd66318,17'd68833,17'd68520,17'd63106,17'd63106,17'd63372,17'd63372,17'd62699,17'd62699,17'd16959,17'd68834,17'd62699,17'd65949,17'd62698,17'd65949,17'd68412,17'd68412,17'd65829,17'd65829,17'd68294,17'd68294,17'd63371,17'd63371,17'd62847,17'd62847,17'd62847,17'd63961,17'd63961,17'd67797,17'd64526,17'd63105,17'd63241,17'd63372,17'd63106,17'd63106,17'd65701,17'd65701,17'd16854,17'd15232,17'd67291,17'd13419,17'd13419,17'd13419,17'd68835,17'd62854,17'd14976,17'd68836,17'd62853,17'd62973,17'd63376,17'd67440,17'd63965,17'd63965,17'd67793,17'd67793,17'd65305,17'd65570,17'd65570,17'd65703,17'd65703,17'd67170,17'd65306,17'd64388,17'd66076,17'd67672,17'd68837,17'd67672,17'd68838,17'd68839,17'd65039,17'd68840,17'd68841,17'd12912,17'd62452,17'd63249,17'd5625,17'd46595,17'd7849,17'd68842,17'd58373,17'd41157,17'd51494,17'd68843,17'd2235,17'd68844,17'd52919,17'd68845,17'd1090,17'd68846,17'd1543,17'd68847
},
'{
17'd4086,17'd3901,17'd3901,17'd3427,17'd2935,17'd3252,17'd10535,17'd1831,17'd4247,17'd4247,17'd1127,17'd14,17'd14,17'd1127,17'd1688,17'd2422,17'd2784,17'd63385,17'd68848,17'd68849,17'd67939,17'd66329,17'd67940,17'd68192,17'd66690,17'd67814,17'd68850,17'd68851,17'd68641,17'd68852,17'd67304,17'd68192,17'd66207,17'd67450,17'd68853,17'd12191,17'd6593,17'd9419,17'd63117,17'd0,17'd10,17'd1128,17'd25,17'd11,17'd18,17'd1277,17'd2257,17'd2257,17'd4247,17'd1831,17'd2422,17'd2935,17'd3901,17'd15877,17'd5204,17'd13943,17'd15496,17'd3428,17'd10802,17'd52621,17'd2258,17'd2597,17'd2257,17'd2257,17'd290,17'd290,17'd3256,17'd3256,17'd2940,17'd3104,17'd3104,17'd4250,17'd5657,17'd5656,17'd27445,17'd11345,17'd7730,17'd7392,17'd7228,17'd7730,17'd68854,17'd11345,17'd11739,17'd12657,17'd65964,17'd68855,17'd68649,17'd68856,17'd64805,17'd68857,17'd68858,17'd68859,17'd68860,17'd39348,17'd66106,17'd39646,17'd28670,17'd18666,17'd68861,17'd68862,17'd68863,17'd68863,17'd68093,17'd12366,17'd10948,17'd10947,17'd10566,17'd21489,17'd30059,17'd30059,17'd68435,17'd49201,17'd63401,17'd5687,17'd4291,17'd59265,17'd52782,17'd52933,17'd64817,17'd58395,17'd58030,17'd52850,17'd48821,17'd56125,17'd57504,17'd48932,17'd58521,17'd58521,17'd54798,17'd54700,17'd65733,17'd55185,17'd59516,17'd60539,17'd68864,17'd68865,17'd65739,17'd55280,17'd64825,17'd68664,17'd56446,17'd64820,17'd64820,17'd55899,17'd68866,17'd65471,17'd68867,17'd64419,17'd68868,17'd60169,17'd54895,17'd54348,17'd68869,17'd68870,17'd68871,17'd68872,17'd68669,17'd67971,17'd68873,17'd68874,17'd68672,17'd68875,17'd68876,17'd68877,17'd68878,17'd68879,17'd68880,17'd68561,17'd68881,17'd61866,17'd68882,17'd68676,17'd68770,17'd68567,17'd68883,17'd68774,17'd68677,17'd68775,17'd67345,17'd68568,17'd68678,17'd68884,17'd54186,17'd52387,17'd68885,17'd68886,17'd68887,17'd68888,17'd9333,17'd8719,17'd8721,17'd15684,17'd24361,17'd24361,17'd9041,17'd24862,17'd16333,17'd10747,17'd7625,17'd68889,17'd68890,17'd68891,17'd7813,17'd11541,17'd132,17'd132,17'd11541,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd130,17'd130,17'd11541,17'd20916,17'd68892,17'd68893,17'd68894,17'd68895,17'd35014,17'd34457,17'd68896,17'd51913,17'd68897,17'd68898,17'd68899,17'd68900,17'd68901,17'd68902,17'd67630,17'd68026,17'd67884,17'd68142,17'd68143,17'd68020,17'd68144,17'd68903,17'd68019,17'd67884,17'd67250,17'd67756,17'd67126,17'd67007,17'd68902,17'd66627,17'd68904,17'd66506,17'd66273,17'd63756,17'd64466,17'd59581,17'd59582,17'd68594,17'd50819,17'd50563,17'd68905,17'd68906,17'd24087,17'd23731,17'd23731,17'd24415,17'd24249,17'd24249,17'd23209,17'd62796,17'd38806,17'd33158,17'd44591,17'd23926,17'd51167,17'd44485,17'd68907,17'd68908,17'd68909,17'd68490,17'd68910,17'd68911,17'd68912,17'd68913,17'd68914,17'd68915,17'd68916,17'd68917,17'd68918,17'd68919,17'd68920,17'd68921,17'd68922,17'd68923,17'd17157,17'd16590,17'd13027,17'd9076,17'd18001,17'd8763,17'd8763,17'd9641,17'd9642,17'd10767,17'd68924,17'd16595,17'd68925,17'd25477,17'd14294,17'd11551,17'd7172,17'd10235,17'd68926,17'd68927,17'd9932,17'd9932,17'd9394,17'd7499,17'd68928,17'd68929,17'd68930,17'd68931,17'd68932,17'd68933,17'd68934,17'd68935,17'd68936,17'd68937,17'd68938,17'd68939,17'd68940,17'd68941,17'd68942,17'd68832,17'd67549,17'd67664,17'd64628,17'd68057,17'd65419,17'd64902,17'd64628,17'd65930,17'd65552,17'd65419,17'd65038,17'd67287,17'd68943,17'd67422,17'd63658,17'd65703,17'd67423,17'd67923,17'd67923,17'd68060,17'd67923,17'd67923,17'd68519,17'd68519,17'd68519,17'd68944,17'd68944,17'd68944,17'd68945,17'd68833,17'd68521,17'd68521,17'd63106,17'd63372,17'd62849,17'd66927,17'd62699,17'd62699,17'd62848,17'd62848,17'd62848,17'd63371,17'd63371,17'd62848,17'd62848,17'd62848,17'd62848,17'd68183,17'd67433,17'd67433,17'd63241,17'd68946,17'd63241,17'd63241,17'd64386,17'd63105,17'd63241,17'd63105,17'd63106,17'd63372,17'd63106,17'd66197,17'd62699,17'd62699,17'd15348,17'd66434,17'd13688,17'd13419,17'd13175,17'd67802,17'd67290,17'd14976,17'd65705,17'd66322,17'd63248,17'd66789,17'd63376,17'd64528,17'd64654,17'd63965,17'd64109,17'd64527,17'd64527,17'd64109,17'd65703,17'd64529,17'd67050,17'd67050,17'd64241,17'd65055,17'd67558,17'd68632,17'd68947,17'd67672,17'd68948,17'd68949,17'd68950,17'd68951,17'd68952,17'd68953,17'd67174,17'd62703,17'd46595,17'd61672,17'd42043,17'd68954,17'd60628,17'd56428,17'd40097,17'd23474,17'd68955,17'd68956,17'd68957,17'd68958,17'd442,17'd68959,17'd15872,17'd68960
},
'{
17'd4086,17'd13943,17'd13943,17'd3901,17'd2934,17'd2935,17'd14070,17'd1831,17'd1688,17'd4247,17'd1127,17'd14,17'd14,17'd14,17'd1688,17'd1831,17'd3252,17'd68191,17'd63977,17'd68755,17'd68304,17'd66686,17'd68961,17'd68961,17'd68962,17'd67063,17'd68850,17'd68963,17'd68963,17'd68754,17'd67572,17'd66937,17'd66329,17'd68964,17'd68965,17'd67815,17'd6894,17'd6734,17'd14867,17'd1830,17'd979,17'd11,17'd20,17'd1128,17'd19,17'd19,17'd17,17'd1414,17'd4247,17'd4247,17'd1831,17'd3252,17'd3427,17'd15496,17'd15496,17'd4086,17'd3592,17'd3901,17'd10924,17'd10669,17'd3429,17'd2258,17'd2257,17'd1414,17'd290,17'd290,17'd3254,17'd3256,17'd2940,17'd2941,17'd3104,17'd3104,17'd5657,17'd5657,17'd12931,17'd6279,17'd7730,17'd7392,17'd7228,17'd7228,17'd7391,17'd11345,17'd6443,17'd5522,17'd66214,17'd34006,17'd67456,17'd68966,17'd68967,17'd68968,17'd32103,17'd67956,17'd7424,17'd39055,17'd49203,17'd52628,17'd7102,17'd40269,17'd19267,17'd68969,17'd68970,17'd68863,17'd68971,17'd68093,17'd21970,17'd11235,17'd10566,17'd10120,17'd24198,17'd30059,17'd68435,17'd10114,17'd5089,17'd5688,17'd4610,17'd4291,17'd59512,17'd52782,17'd52933,17'd58395,17'd59012,17'd58030,17'd56343,17'd55483,17'd53950,17'd64820,17'd56446,17'd58649,17'd65737,17'd65859,17'd53951,17'd54253,17'd54618,17'd59516,17'd60539,17'd68445,17'd68972,17'd63545,17'd56028,17'd55093,17'd54893,17'd54993,17'd58150,17'd54252,17'd54987,17'd56233,17'd54799,17'd64283,17'd60538,17'd60654,17'd54432,17'd68973,17'd68974,17'd68975,17'd68976,17'd68872,17'd68669,17'd67971,17'd68977,17'd68874,17'd68978,17'd68979,17'd68876,17'd68980,17'd68559,17'd68981,17'd68982,17'd68983,17'd68881,17'd61465,17'd68984,17'd68985,17'd68986,17'd68987,17'd68988,17'd68989,17'd68774,17'd68775,17'd68990,17'd68991,17'd68678,17'd68884,17'd68992,17'd10139,17'd68993,17'd68994,17'd68995,17'd68996,17'd68997,17'd8722,17'd9348,17'd9040,17'd9039,17'd17123,17'd9195,17'd24545,17'd16690,17'd14938,17'd21511,17'd17976,17'd68890,17'd63047,17'd53258,17'd131,17'd132,17'd132,17'd11541,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd11541,17'd52245,17'd21681,17'd68998,17'd68999,17'd69000,17'd51562,17'd22338,17'd21848,17'd22008,17'd69001,17'd40221,17'd69002,17'd64733,17'd69003,17'd50459,17'd66392,17'd66756,17'd67006,17'd69004,17'd68792,17'd69005,17'd67884,17'd67886,17'd67886,17'd67520,17'd67383,17'd67630,17'd67757,17'd67254,17'd60980,17'd67632,17'd66757,17'd66275,17'd61900,17'd57833,17'd50728,17'd64730,17'd51553,17'd67256,17'd57839,17'd58459,17'd24091,17'd23382,17'd30879,17'd30879,17'd24090,17'd24090,17'd23731,17'd24086,17'd26396,17'd69006,17'd22501,17'd22331,17'd36289,17'd37408,17'd69007,17'd69008,17'd45498,17'd69009,17'd69010,17'd69011,17'd69012,17'd69013,17'd69014,17'd69015,17'd68269,17'd69016,17'd69017,17'd68917,17'd68918,17'd68919,17'd69018,17'd69019,17'd68922,17'd69020,17'd16471,17'd69021,17'd69022,17'd11993,17'd8615,17'd8763,17'd12137,17'd9641,17'd8917,17'd17641,17'd69023,17'd69024,17'd69025,17'd69026,17'd14159,17'd69027,17'd7663,17'd11848,17'd69028,17'd68927,17'd9932,17'd9394,17'd8780,17'd29740,17'd68928,17'd68824,17'd69029,17'd68931,17'd68932,17'd69030,17'd69031,17'd68935,17'd68936,17'd69032,17'd69033,17'd69034,17'd68940,17'd68941,17'd69035,17'd67661,17'd69036,17'd67664,17'd64628,17'd64628,17'd64902,17'd64902,17'd64902,17'd69037,17'd65552,17'd65419,17'd65815,17'd67287,17'd69038,17'd66321,17'd64109,17'd63965,17'd64529,17'd68292,17'd67423,17'd67923,17'd67923,17'd67923,17'd68519,17'd68519,17'd68519,17'd68944,17'd68944,17'd68944,17'd68945,17'd68833,17'd68520,17'd68520,17'd63962,17'd63106,17'd63372,17'd62849,17'd62699,17'd62699,17'd62848,17'd62848,17'd62848,17'd62848,17'd68183,17'd68183,17'd68183,17'd68183,17'd68183,17'd68183,17'd63104,17'd63104,17'd68946,17'd68946,17'd63241,17'd63105,17'd64386,17'd63105,17'd63241,17'd64386,17'd63106,17'd63106,17'd65950,17'd66197,17'd65830,17'd16959,17'd15232,17'd62447,17'd13688,17'd13419,17'd13175,17'd67289,17'd67288,17'd65705,17'd68836,17'd66678,17'd66789,17'd65286,17'd66321,17'd66548,17'd64654,17'd63965,17'd64109,17'd64527,17'd64527,17'd64109,17'd65703,17'd64529,17'd67050,17'd65306,17'd64388,17'd66320,17'd67672,17'd68632,17'd68947,17'd69039,17'd69040,17'd69041,17'd69042,17'd69043,17'd68634,17'd12481,17'd69044,17'd18864,17'd69045,17'd69046,17'd4393,17'd69047,17'd60628,17'd19360,17'd39028,17'd56886,17'd19099,17'd40098,17'd61543,17'd1959,17'd20008,17'd68959,17'd69048,17'd648
},
'{
17'd6730,17'd4086,17'd13943,17'd3592,17'd2934,17'd3101,17'd14070,17'd1831,17'd1688,17'd1688,17'd1127,17'd14,17'd14,17'd14,17'd4247,17'd1831,17'd10535,17'd2592,17'd69049,17'd69050,17'd69051,17'd69052,17'd66686,17'd67446,17'd67941,17'd66940,17'd68640,17'd69053,17'd69054,17'd68080,17'd69055,17'd66940,17'd67568,17'd66207,17'd65959,17'd69056,17'd68645,17'd6593,17'd63520,17'd14742,17'd5969,17'd10,17'd2598,17'd20,17'd11,17'd18,17'd16,17'd1416,17'd4247,17'd4247,17'd1688,17'd2422,17'd3101,17'd3428,17'd15496,17'd3592,17'd3592,17'd3901,17'd2934,17'd2935,17'd52621,17'd2258,17'd2257,17'd1414,17'd290,17'd290,17'd1129,17'd1129,17'd2941,17'd2941,17'd3104,17'd3104,17'd5658,17'd5657,17'd5804,17'd6746,17'd10408,17'd10409,17'd7228,17'd7228,17'd7392,17'd10672,17'd10548,17'd5662,17'd5381,17'd33054,17'd69057,17'd69058,17'd69059,17'd69060,17'd66102,17'd69061,17'd65595,17'd69062,17'd52377,17'd51773,17'd69063,17'd69064,17'd69065,17'd67586,17'd13331,17'd69066,17'd68863,17'd69067,17'd68094,17'd69068,17'd12961,17'd20435,17'd24198,17'd10118,17'd10116,17'd10114,17'd6139,17'd5089,17'd4925,17'd4928,17'd4291,17'd59512,17'd58760,17'd69069,17'd59012,17'd57263,17'd57120,17'd57123,17'd53810,17'd54093,17'd58400,17'd58150,17'd68443,17'd65859,17'd57267,17'd53950,17'd66349,17'd54705,17'd56689,17'd69070,17'd69071,17'd58402,17'd55582,17'd56582,17'd58522,17'd56020,17'd65734,17'd65982,17'd56021,17'd54803,17'd56241,17'd64144,17'd64144,17'd56904,17'd54803,17'd57505,17'd69072,17'd69073,17'd69074,17'd69075,17'd69076,17'd69077,17'd68977,17'd69078,17'd68978,17'd68875,17'd69079,17'd69080,17'd68879,17'd69081,17'd69082,17'd69083,17'd68881,17'd61464,17'd69084,17'd69085,17'd69086,17'd69087,17'd69088,17'd68989,17'd69089,17'd68775,17'd68990,17'd69090,17'd69091,17'd69092,17'd17111,17'd69093,17'd69094,17'd36477,17'd8716,17'd69095,17'd45812,17'd8728,17'd8725,17'd8878,17'd15684,17'd23859,17'd9195,17'd8576,17'd16803,17'd14938,17'd8738,17'd69096,17'd69097,17'd69098,17'd53258,17'd132,17'd130,17'd133,17'd11541,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd52492,17'd52812,17'd68893,17'd69099,17'd68895,17'd35154,17'd35156,17'd31497,17'd22160,17'd22326,17'd51552,17'd58821,17'd58824,17'd65138,17'd67889,17'd69100,17'd69101,17'd69102,17'd67004,17'd69103,17'd67249,17'd67382,17'd67251,17'd67383,17'd61759,17'd69104,17'd69105,17'd61240,17'd60588,17'd61762,17'd61768,17'd63607,17'd58210,17'd50645,17'd64730,17'd50650,17'd69106,17'd57205,17'd30424,17'd23731,17'd69107,17'd24414,17'd28975,17'd29100,17'd24088,17'd25439,17'd24086,17'd29099,17'd69006,17'd45381,17'd22856,17'd32660,17'd31498,17'd69108,17'd69109,17'd69110,17'd41129,17'd62169,17'd69111,17'd69112,17'd68707,17'd69113,17'd69114,17'd69115,17'd68606,17'd69116,17'd69117,17'd69118,17'd69119,17'd68812,17'd16714,17'd69120,17'd69121,17'd69122,17'd69123,17'd69124,17'd69125,17'd11993,17'd8615,17'd8614,17'd13672,17'd8762,17'd8917,17'd12139,17'd69126,17'd15464,17'd69127,17'd68401,17'd14561,17'd9221,17'd7174,17'd68822,17'd69028,17'd69128,17'd9932,17'd9394,17'd8780,17'd27696,17'd68510,17'd68824,17'd69129,17'd69130,17'd69131,17'd69132,17'd69133,17'd69134,17'd69135,17'd69136,17'd69137,17'd69034,17'd69138,17'd69139,17'd69140,17'd67548,17'd67420,17'd65163,17'd69141,17'd64628,17'd64628,17'd64902,17'd64902,17'd69142,17'd68058,17'd65815,17'd65164,17'd65039,17'd69143,17'd66321,17'd64109,17'd63965,17'd64529,17'd68292,17'd68292,17'd68517,17'd67923,17'd69144,17'd68519,17'd68519,17'd68519,17'd68944,17'd68944,17'd68944,17'd69145,17'd69145,17'd68833,17'd68833,17'd64650,17'd64526,17'd64386,17'd63106,17'd63372,17'd63372,17'd63105,17'd63105,17'd64386,17'd64386,17'd63106,17'd63106,17'd68295,17'd68183,17'd68295,17'd68183,17'd63241,17'd68946,17'd63241,17'd63241,17'd63105,17'd63105,17'd64386,17'd63105,17'd63105,17'd64386,17'd63106,17'd63106,17'd65830,17'd65566,17'd64531,17'd15483,17'd66434,17'd67428,17'd13688,17'd13175,17'd13570,17'd14175,17'd69146,17'd16255,17'd68416,17'd66536,17'd65286,17'd67422,17'd63377,17'd64653,17'd63965,17'd64109,17'd64109,17'd64527,17'd64527,17'd64109,17'd64110,17'd65306,17'd65306,17'd64241,17'd64921,17'd67439,17'd68632,17'd69147,17'd67673,17'd66199,17'd66198,17'd69143,17'd63110,17'd15734,17'd62976,17'd18269,17'd69148,17'd62977,17'd69149,17'd48385,17'd8481,17'd69047,17'd60628,17'd57615,17'd57489,17'd69150,17'd57748,17'd69151,17'd69152,17'd20270,17'd801,17'd69153,17'd69154,17'd2251
},
'{
17'd14744,17'd4893,17'd4737,17'd4086,17'd3901,17'd2934,17'd2935,17'd3250,17'd1688,17'd1688,17'd1127,17'd14,17'd14,17'd14,17'd1127,17'd4247,17'd10535,17'd2422,17'd69155,17'd64929,17'd69156,17'd69157,17'd66686,17'd67446,17'd67687,17'd66690,17'd67571,17'd68852,17'd69158,17'd69158,17'd69159,17'd69160,17'd67180,17'd66686,17'd66088,17'd68313,17'd67815,17'd69161,17'd9270,17'd64125,17'd9422,17'd3748,17'd1128,17'd10,17'd10,17'd3905,17'd16,17'd1416,17'd1127,17'd4247,17'd1688,17'd1688,17'd3252,17'd3251,17'd3428,17'd15496,17'd3901,17'd3901,17'd2934,17'd3101,17'd52621,17'd3429,17'd2596,17'd1415,17'd30,17'd30,17'd1129,17'd1129,17'd2941,17'd2941,17'd3104,17'd3104,17'd3435,17'd5658,17'd5657,17'd11889,17'd11211,17'd10409,17'd7228,17'd7064,17'd7228,17'd7730,17'd6281,17'd5662,17'd5384,17'd66694,17'd68428,17'd69162,17'd69163,17'd69164,17'd69165,17'd69166,17'd69167,17'd39347,17'd69168,17'd38351,17'd69169,17'd69170,17'd25913,17'd69171,17'd42660,17'd13215,17'd69066,17'd69067,17'd68971,17'd68094,17'd13098,17'd12068,17'd20435,17'd24198,17'd9578,17'd9441,17'd10114,17'd9303,17'd5089,17'd4925,17'd4610,17'd4291,17'd59512,17'd52782,17'd68096,17'd59012,17'd57012,17'd56343,17'd53810,17'd54021,17'd57773,17'd58649,17'd69172,17'd65603,17'd58399,17'd55576,17'd55576,17'd64820,17'd54992,17'd56028,17'd57395,17'd55182,17'd63405,17'd55582,17'd56580,17'd56688,17'd65735,17'd56021,17'd57387,17'd58401,17'd55092,17'd55183,17'd68098,17'd55676,17'd55184,17'd65733,17'd3777,17'd69173,17'd69174,17'd69175,17'd69176,17'd69077,17'd69177,17'd69178,17'd68978,17'd69179,17'd69180,17'd69181,17'd68981,17'd69182,17'd69183,17'd69184,17'd68881,17'd61336,17'd69185,17'd69186,17'd69187,17'd69188,17'd69088,17'd69189,17'd68989,17'd15280,17'd69190,17'd69191,17'd69192,17'd69092,17'd69193,17'd69194,17'd69195,17'd69196,17'd69197,17'd69198,17'd48001,17'd8571,17'd11966,17'd24368,17'd24999,17'd23859,17'd26154,17'd26155,17'd61747,17'd7621,17'd8263,17'd17857,17'd68890,17'd69199,17'd53258,17'd132,17'd130,17'd133,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd52245,17'd69200,17'd21070,17'd69201,17'd21382,17'd51563,17'd35154,17'd32498,17'd22507,17'd33311,17'd37116,17'd23736,17'd23734,17'd55228,17'd56507,17'd52815,17'd60360,17'd69202,17'd50644,17'd69203,17'd69204,17'd69205,17'd66627,17'd67887,17'd67130,17'd60717,17'd66629,17'd62784,17'd61900,17'd57833,17'd50728,17'd59085,17'd64730,17'd51553,17'd67256,17'd62797,17'd53405,17'd30424,17'd30879,17'd28849,17'd31047,17'd26280,17'd28975,17'd45493,17'd36701,17'd35577,17'd35166,17'd30579,17'd55227,17'd22851,17'd22157,17'd44825,17'd50073,17'd69206,17'd45622,17'd69207,17'd42019,17'd69208,17'd69209,17'd69210,17'd69211,17'd69212,17'd69213,17'd69214,17'd69016,17'd69215,17'd69216,17'd68811,17'd69119,17'd68812,17'd68921,17'd69217,17'd69218,17'd69218,17'd69219,17'd69220,17'd9773,17'd8295,17'd8294,17'd8294,17'd8293,17'd12137,17'd8763,17'd11988,17'd69221,17'd15212,17'd69222,17'd25876,17'd14158,17'd8292,17'd10235,17'd68926,17'd68927,17'd69223,17'd9394,17'd9394,17'd28184,17'd27696,17'd68510,17'd69224,17'd69225,17'd69226,17'd69227,17'd69228,17'd69229,17'd69230,17'd69231,17'd69232,17'd69233,17'd69234,17'd69235,17'd69236,17'd66784,17'd67160,17'd65683,17'd65037,17'd69141,17'd69141,17'd69141,17'd64628,17'd69237,17'd67918,17'd67791,17'd65164,17'd68290,17'd67422,17'd63246,17'd63377,17'd64527,17'd64109,17'd65703,17'd64529,17'd68292,17'd68517,17'd68059,17'd69144,17'd68519,17'd68519,17'd68519,17'd68944,17'd68944,17'd68944,17'd69145,17'd69145,17'd68945,17'd68833,17'd69238,17'd64650,17'd64526,17'd64526,17'd63962,17'd63962,17'd64386,17'd64526,17'd64526,17'd64526,17'd63962,17'd63962,17'd68295,17'd68183,17'd68295,17'd68183,17'd63241,17'd63241,17'd63105,17'd63105,17'd64386,17'd63105,17'd64386,17'd63105,17'd63105,17'd63106,17'd63962,17'd66197,17'd65830,17'd64244,17'd68834,17'd69239,17'd67428,17'd67428,17'd14175,17'd13570,17'd13570,17'd62576,17'd67038,17'd69240,17'd68741,17'd64630,17'd67422,17'd69241,17'd63657,17'd64653,17'd67793,17'd64109,17'd64109,17'd64109,17'd64109,17'd63965,17'd65306,17'd65306,17'd64241,17'd64921,17'd66320,17'd68187,17'd69147,17'd69147,17'd69039,17'd69242,17'd69243,17'd67422,17'd66678,17'd15734,17'd62976,17'd65058,17'd18382,17'd63111,17'd46354,17'd4056,17'd8481,17'd68954,17'd60628,17'd59909,17'd69244,17'd69245,17'd54776,17'd69246,17'd2411,17'd772,17'd801,17'd69153,17'd69247,17'd2251
},
'{
17'd7049,17'd64660,17'd4737,17'd4086,17'd3901,17'd2934,17'd2935,17'd3250,17'd1688,17'd1688,17'd1127,17'd14,17'd14,17'd14,17'd1127,17'd4247,17'd1831,17'd2422,17'd68075,17'd69248,17'd69249,17'd69250,17'd67939,17'd67685,17'd69251,17'd67181,17'd66939,17'd67813,17'd69158,17'd69252,17'd68424,17'd69253,17'd66690,17'd69254,17'd66554,17'd65959,17'd69156,17'd7547,17'd10922,17'd69255,17'd65450,17'd1276,17'd1128,17'd808,17'd10,17'd4089,17'd16,17'd17,17'd1127,17'd1127,17'd1689,17'd1688,17'd2422,17'd3101,17'd34512,17'd15358,17'd3427,17'd3427,17'd3101,17'd3101,17'd52621,17'd2258,17'd1414,17'd1415,17'd1414,17'd1414,17'd30,17'd30,17'd3254,17'd3254,17'd2941,17'd3104,17'd3435,17'd3435,17'd5657,17'd5804,17'd11211,17'd6904,17'd7063,17'd7063,17'd7064,17'd7228,17'd7392,17'd6111,17'd5976,17'd4898,17'd69256,17'd69257,17'd69258,17'd69259,17'd69260,17'd69261,17'd69262,17'd69263,17'd69264,17'd38094,17'd69265,17'd69266,17'd69267,17'd7263,17'd8850,17'd42348,17'd13098,17'd68862,17'd68764,17'd69268,17'd69068,17'd12961,17'd10698,17'd9845,17'd9705,17'd9578,17'd68095,17'd10114,17'd6304,17'd5088,17'd5688,17'd4768,17'd4769,17'd59513,17'd58759,17'd68096,17'd52710,17'd52850,17'd58519,17'd53950,17'd54020,17'd64820,17'd55776,17'd54252,17'd58031,17'd55668,17'd53950,17'd58272,17'd54993,17'd69269,17'd56240,17'd65207,17'd63405,17'd69270,17'd69271,17'd60539,17'd65605,17'd56241,17'd55092,17'd56582,17'd56026,17'd69272,17'd69272,17'd55183,17'd55280,17'd57268,17'd3620,17'd69073,17'd69273,17'd69274,17'd69275,17'd69276,17'd69277,17'd69178,17'd68978,17'd69278,17'd69080,17'd69279,17'd69280,17'd69281,17'd69282,17'd69283,17'd69284,17'd69285,17'd69286,17'd69287,17'd69288,17'd69188,17'd69289,17'd69290,17'd68989,17'd15544,17'd69291,17'd69292,17'd69293,17'd11100,17'd10707,17'd69294,17'd69295,17'd69296,17'd69297,17'd8239,17'd10858,17'd24862,17'd35514,17'd11966,17'd24999,17'd29637,17'd26259,17'd13256,17'd11279,17'd14269,17'd20615,17'd55527,17'd69298,17'd65766,17'd20188,17'd132,17'd1481,17'd1481,17'd132,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd131,17'd20626,17'd69299,17'd69300,17'd69301,17'd69302,17'd47067,17'd42602,17'd21697,17'd35153,17'd22330,17'd32008,17'd29827,17'd23918,17'd30127,17'd24421,17'd39133,17'd59858,17'd69303,17'd64874,17'd69304,17'd69100,17'd69305,17'd63896,17'd63756,17'd63756,17'd69306,17'd58585,17'd69307,17'd59582,17'd68594,17'd52161,17'd57967,17'd50563,17'd58459,17'd33801,17'd24087,17'd24086,17'd23564,17'd29972,17'd34299,17'd45163,17'd24086,17'd35999,17'd23921,17'd35166,17'd36414,17'd36543,17'd23219,17'd69308,17'd22166,17'd32664,17'd47939,17'd48158,17'd47057,17'd69309,17'd69310,17'd69311,17'd69312,17'd69313,17'd69314,17'd69315,17'd69316,17'd69317,17'd69318,17'd69319,17'd69320,17'd69321,17'd68812,17'd68718,17'd69020,17'd69322,17'd69323,17'd69323,17'd14705,17'd10369,17'd11165,17'd11994,17'd13400,17'd15459,17'd69324,17'd12282,17'd8917,17'd18480,17'd69221,17'd17055,17'd66656,17'd16479,17'd12885,17'd7172,17'd10235,17'd12301,17'd68927,17'd69223,17'd26219,17'd26219,17'd28184,17'd27696,17'd68510,17'd69325,17'd69326,17'd69131,17'd69327,17'd69227,17'd69132,17'd69328,17'd69329,17'd69330,17'd69331,17'd69332,17'd69333,17'd69236,17'd66784,17'd67160,17'd65551,17'd64505,17'd69141,17'd69141,17'd69141,17'd64902,17'd69334,17'd69335,17'd69336,17'd66788,17'd67440,17'd63378,17'd64652,17'd64109,17'd64527,17'd64109,17'd65703,17'd65703,17'd67423,17'd67923,17'd68059,17'd68059,17'd68182,17'd68060,17'd68519,17'd68944,17'd68944,17'd68944,17'd69337,17'd69337,17'd69145,17'd69145,17'd69145,17'd69338,17'd69339,17'd69339,17'd64650,17'd64650,17'd69338,17'd69338,17'd69338,17'd69338,17'd64526,17'd64386,17'd64386,17'd63105,17'd63372,17'd62969,17'd62969,17'd63372,17'd63106,17'd63106,17'd63106,17'd63372,17'd69340,17'd69340,17'd63106,17'd63106,17'd63962,17'd66197,17'd65830,17'd68834,17'd15232,17'd67428,17'd67429,17'd62447,17'd69341,17'd13570,17'd14175,17'd62449,17'd16255,17'd68416,17'd66536,17'd64767,17'd67422,17'd68415,17'd63657,17'd63657,17'd67793,17'd67793,17'd64109,17'd64109,17'd63965,17'd63965,17'd65306,17'd65306,17'd64921,17'd65055,17'd67439,17'd68632,17'd69147,17'd68837,17'd68633,17'd66198,17'd63511,17'd67440,17'd62852,17'd69342,17'd67290,17'd14175,17'd62855,17'd67166,17'd69343,17'd49196,17'd5932,17'd50002,17'd58008,17'd57749,17'd69344,17'd69345,17'd629,17'd3095,17'd1679,17'd607,17'd2778,17'd69346,17'd1548,17'd253
},
'{
17'd67065,17'd64392,17'd14443,17'd4893,17'd13943,17'd3751,17'd2593,17'd2784,17'd2422,17'd1688,17'd4247,17'd14,17'd14,17'd14,17'd14,17'd1127,17'd1688,17'd3250,17'd7371,17'd69347,17'd65713,17'd68849,17'd66554,17'd66443,17'd69348,17'd67303,17'd67449,17'd68640,17'd68080,17'd69252,17'd68308,17'd69055,17'd69349,17'd67687,17'd67446,17'd69350,17'd68849,17'd8043,17'd10665,17'd6433,17'd10544,17'd1277,17'd18,17'd808,17'd10,17'd20404,17'd18,17'd1277,17'd1127,17'd1127,17'd1689,17'd1688,17'd2422,17'd2422,17'd3251,17'd37047,17'd3427,17'd3427,17'd3101,17'd3101,17'd52621,17'd3429,17'd2596,17'd1415,17'd1415,17'd1414,17'd30,17'd30,17'd31,17'd3254,17'd2941,17'd2941,17'd3104,17'd3435,17'd5657,17'd5804,17'd6746,17'd10408,17'd9970,17'd7063,17'd7064,17'd6907,17'd7227,17'd10672,17'd11738,17'd69351,17'd33055,17'd69352,17'd69353,17'd69354,17'd69355,17'd69356,17'd69357,17'd69358,17'd69359,17'd69360,17'd69361,17'd6783,17'd69362,17'd6942,17'd7760,17'd8699,17'd9847,17'd11766,17'd13608,17'd69268,17'd69068,17'd21970,17'd12068,17'd11765,17'd10120,17'd10118,17'd29181,17'd28669,17'd6304,17'd6138,17'd5088,17'd4610,17'd4768,17'd4769,17'd69363,17'd58641,17'd68096,17'd52710,17'd53370,17'd66457,17'd54254,17'd54171,17'd59646,17'd65328,17'd66226,17'd57772,17'd58272,17'd54614,17'd56446,17'd69364,17'd69365,17'd55907,17'd67472,17'd67593,17'd67593,17'd69366,17'd67472,17'd63543,17'd56026,17'd59013,17'd60657,17'd60657,17'd56026,17'd55183,17'd55380,17'd65733,17'd57381,17'd68446,17'd69367,17'd69368,17'd69369,17'd69370,17'd69371,17'd69372,17'd68978,17'd69276,17'd69181,17'd69373,17'd69182,17'd69374,17'd69375,17'd69376,17'd68881,17'd69377,17'd60814,17'd69378,17'd69379,17'd69380,17'd69289,17'd17706,17'd68989,17'd15544,17'd69291,17'd14787,17'd16672,17'd69381,17'd20302,17'd69382,17'd69383,17'd69384,17'd69385,17'd69386,17'd8414,17'd25147,17'd11531,17'd8572,17'd9046,17'd29920,17'd26259,17'd13256,17'd11279,17'd14269,17'd19784,17'd69387,17'd69388,17'd10869,17'd20188,17'd132,17'd130,17'd1197,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd131,17'd5593,17'd20629,17'd69389,17'd69390,17'd69301,17'd69391,17'd51382,17'd43428,17'd52171,17'd46099,17'd22328,17'd23387,17'd23565,17'd23733,17'd23918,17'd29376,17'd24421,17'd34112,17'd59453,17'd56507,17'd51074,17'd50819,17'd63473,17'd65376,17'd59861,17'd68701,17'd58207,17'd67256,17'd51735,17'd57839,17'd56966,17'd29527,17'd29528,17'd29241,17'd23733,17'd23918,17'd23565,17'd29242,17'd28976,17'd26397,17'd23920,17'd35721,17'd39134,17'd42161,17'd42610,17'd43986,17'd34759,17'd30580,17'd69392,17'd22002,17'd35154,17'd48058,17'd69393,17'd69394,17'd21549,17'd69395,17'd69396,17'd69397,17'd68601,17'd25743,17'd28627,17'd69398,17'd69399,17'd69400,17'd68613,17'd69401,17'd68613,17'd68919,17'd69402,17'd69403,17'd69323,17'd69404,17'd69405,17'd69406,17'd69407,17'd9774,17'd9649,17'd9230,17'd15209,17'd15459,17'd8294,17'd8763,17'd18480,17'd11552,17'd25763,17'd69408,17'd69409,17'd20108,17'd7173,17'd68822,17'd69028,17'd69128,17'd11430,17'd26219,17'd26219,17'd28184,17'd27696,17'd68510,17'd69410,17'd69411,17'd69131,17'd69412,17'd69327,17'd69228,17'd69413,17'd69329,17'd69414,17'd69415,17'd69416,17'd69333,17'd69236,17'd69140,17'd67160,17'd65551,17'd69141,17'd69417,17'd69418,17'd69418,17'd64628,17'd69419,17'd69420,17'd68299,17'd63378,17'd63964,17'd63808,17'd64527,17'd64109,17'd64527,17'd64109,17'd65570,17'd65703,17'd67423,17'd67923,17'd68059,17'd68059,17'd68060,17'd68060,17'd68519,17'd68944,17'd68944,17'd68944,17'd69337,17'd69337,17'd69145,17'd69145,17'd69145,17'd69145,17'd69421,17'd69421,17'd69238,17'd69238,17'd69338,17'd69338,17'd69338,17'd69422,17'd64526,17'd64386,17'd63105,17'd63105,17'd62969,17'd62969,17'd63372,17'd63106,17'd63962,17'd63962,17'd63106,17'd63372,17'd69340,17'd68521,17'd63962,17'd63962,17'd66197,17'd66197,17'd68834,17'd16959,17'd67428,17'd67429,17'd67429,17'd62447,17'd69341,17'd14175,17'd69341,17'd62449,17'd17543,17'd68741,17'd64630,17'd67421,17'd69241,17'd67932,17'd64111,17'd69423,17'd68297,17'd67793,17'd64109,17'd63965,17'd64654,17'd64654,17'd64241,17'd67436,17'd65055,17'd67296,17'd67672,17'd69424,17'd68837,17'd69425,17'd69426,17'd66074,17'd63511,17'd67440,17'd62852,17'd14734,17'd67290,17'd69341,17'd62855,17'd69427,17'd69428,17'd59620,17'd7191,17'd40715,17'd51580,17'd58245,17'd54877,17'd1265,17'd2249,17'd2764,17'd260,17'd271,17'd2778,17'd69153,17'd402,17'd69429
},
'{
17'd69430,17'd5376,17'd64660,17'd4893,17'd4086,17'd3427,17'd3101,17'd3252,17'd1831,17'd1831,17'd4247,17'd1127,17'd14,17'd14,17'd14,17'd1127,17'd1688,17'd1688,17'd2422,17'd11887,17'd64396,17'd67683,17'd66441,17'd66443,17'd69431,17'd69432,17'd68526,17'd69433,17'd68424,17'd69252,17'd69434,17'd69159,17'd69435,17'd69436,17'd66554,17'd66089,17'd68965,17'd8344,17'd11069,17'd9270,17'd64125,17'd1830,17'd19,17'd11,17'd10,17'd10,17'd18,17'd1277,17'd14,17'd1967,17'd1127,17'd4247,17'd1688,17'd1831,17'd14070,17'd38864,17'd34512,17'd34512,17'd3251,17'd3101,17'd52621,17'd3429,17'd2596,17'd2936,17'd1415,17'd1415,17'd1414,17'd30,17'd31,17'd31,17'd2941,17'd2941,17'd3104,17'd3435,17'd5657,17'd5804,17'd6746,17'd6599,17'd6600,17'd6747,17'd69437,17'd7390,17'd8048,17'd10408,17'd69438,17'd69439,17'd69440,17'd69441,17'd69442,17'd69443,17'd69444,17'd69445,17'd46250,17'd69358,17'd7920,17'd38479,17'd69446,17'd69447,17'd69448,17'd38480,17'd69449,17'd36764,17'd16042,17'd69450,17'd11482,17'd12366,17'd69451,17'd69451,17'd12364,17'd12364,17'd22285,17'd11916,17'd29181,17'd28669,17'd9985,17'd8846,17'd6137,17'd5998,17'd4768,17'd4291,17'd65979,17'd69452,17'd58266,17'd66347,17'd59012,17'd57012,17'd53447,17'd58029,17'd54433,17'd59646,17'd57126,17'd65734,17'd56804,17'd58649,17'd56446,17'd54894,17'd65082,17'd59930,17'd55780,17'd57508,17'd63689,17'd63405,17'd55182,17'd55182,17'd55378,17'd57277,17'd69453,17'd69454,17'd56023,17'd64420,17'd55184,17'd57773,17'd52933,17'd69455,17'd69456,17'd69457,17'd69458,17'd69459,17'd69460,17'd69461,17'd69462,17'd69276,17'd69463,17'd69464,17'd69465,17'd69466,17'd69467,17'd69468,17'd69469,17'd69470,17'd61332,17'd69471,17'd69472,17'd69473,17'd69474,17'd17706,17'd69475,17'd15156,17'd69476,17'd69477,17'd69478,17'd10953,17'd20302,17'd69479,17'd69480,17'd69481,17'd69482,17'd8094,17'd24042,17'd8579,17'd9887,17'd8571,17'd8724,17'd9046,17'd12425,17'd13256,17'd59708,17'd14269,17'd63185,17'd15953,17'd69483,17'd10869,17'd53258,17'd130,17'd130,17'd356,17'd132,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd136,17'd136,17'd130,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd5593,17'd20623,17'd65635,17'd69484,17'd69485,17'd69486,17'd51222,17'd51382,17'd42602,17'd21694,17'd35157,17'd23570,17'd42611,17'd23565,17'd23564,17'd34137,17'd34137,17'd23564,17'd28722,17'd23731,17'd24249,17'd30431,17'd29375,17'd29527,17'd29527,17'd29375,17'd30431,17'd24249,17'd23917,17'd30879,17'd28722,17'd23732,17'd23733,17'd23733,17'd31502,17'd29099,17'd23566,17'd23387,17'd23387,17'd26396,17'd23211,17'd23736,17'd34298,17'd36139,17'd32202,17'd40523,17'd22157,17'd69487,17'd69488,17'd22000,17'd51562,17'd47749,17'd69489,17'd69490,17'd69491,17'd69492,17'd43446,17'd69493,17'd69494,17'd69495,17'd69496,17'd69497,17'd69498,17'd68917,17'd68717,17'd69499,17'd69500,17'd68919,17'd69501,17'd69322,17'd69502,17'd69503,17'd69504,17'd69505,17'd69506,17'd69507,17'd69508,17'd8297,17'd9380,17'd69509,17'd12283,17'd9642,17'd11988,17'd17641,17'd25620,17'd69510,17'd17168,17'd8611,17'd7175,17'd11850,17'd68927,17'd69223,17'd11430,17'd26219,17'd26219,17'd28184,17'd9933,17'd68622,17'd69511,17'd69512,17'd69513,17'd69412,17'd69327,17'd69514,17'd69515,17'd69516,17'd69517,17'd69518,17'd69416,17'd69333,17'd69236,17'd69519,17'd69520,17'd65285,17'd69141,17'd69417,17'd69418,17'd69521,17'd65552,17'd69335,17'd69522,17'd63964,17'd66073,17'd66676,17'd66437,17'd65569,17'd65570,17'd65570,17'd65570,17'd65703,17'd67423,17'd67923,17'd68059,17'd69523,17'd69524,17'd68182,17'd68060,17'd69525,17'd69525,17'd68944,17'd69337,17'd69337,17'd69337,17'd69145,17'd69145,17'd69145,17'd69145,17'd69145,17'd69338,17'd69338,17'd69338,17'd69526,17'd69526,17'd69422,17'd69422,17'd67044,17'd67046,17'd63105,17'd63105,17'd62969,17'd63372,17'd68295,17'd68295,17'd63106,17'd63106,17'd63106,17'd63106,17'd69340,17'd68521,17'd69527,17'd63962,17'd66197,17'd65950,17'd16959,17'd15999,17'd67429,17'd67428,17'd67290,17'd62576,17'd62576,17'd62576,17'd62449,17'd67427,17'd17543,17'd65689,17'd69528,17'd68740,17'd68415,17'd69243,17'd64388,17'd69529,17'd69530,17'd69531,17'd64109,17'd63965,17'd64654,17'd64922,17'd64241,17'd64789,17'd65831,17'd67439,17'd68632,17'd69424,17'd68947,17'd68633,17'd66199,17'd66075,17'd64528,17'd65951,17'd62851,17'd15483,17'd15618,17'd15618,17'd69532,17'd69533,17'd47767,17'd4553,17'd5494,17'd55166,17'd69534,17'd69535,17'd18144,17'd232,17'd5050,17'd1668,17'd425,17'd642,17'd255,17'd69536,17'd1683,17'd69537
},
'{
17'd69538,17'd5645,17'd9959,17'd6730,17'd4086,17'd3901,17'd3427,17'd3101,17'd2422,17'd1831,17'd1688,17'd1127,17'd14,17'd14,17'd14,17'd1127,17'd1831,17'd1831,17'd10535,17'd6265,17'd63977,17'd65840,17'd66553,17'd66686,17'd69431,17'd69431,17'd67181,17'd66812,17'd69539,17'd69252,17'd69158,17'd68308,17'd68426,17'd68644,17'd66686,17'd66089,17'd67450,17'd68853,17'd7220,17'd66942,17'd12783,17'd63118,17'd1,17'd1128,17'd10,17'd808,17'd20404,17'd18,17'd14,17'd14,17'd1127,17'd4247,17'd1688,17'd1688,17'd3252,17'd38864,17'd37047,17'd34512,17'd3251,17'd3101,17'd52621,17'd3429,17'd2596,17'd2936,17'd1415,17'd1415,17'd1414,17'd1414,17'd30,17'd31,17'd3255,17'd2941,17'd2941,17'd3435,17'd3756,17'd5804,17'd6746,17'd6439,17'd6904,17'd6747,17'd6601,17'd7390,17'd8048,17'd7556,17'd7731,17'd69540,17'd69541,17'd3443,17'd69542,17'd69543,17'd69544,17'd69545,17'd69546,17'd69547,17'd25125,17'd7920,17'd69548,17'd69446,17'd69549,17'd38095,17'd37970,17'd36057,17'd13612,17'd29182,17'd10288,17'd11235,17'd12364,17'd21970,17'd21970,17'd12364,17'd12683,17'd12536,17'd10432,17'd68095,17'd10114,17'd6304,17'd8846,17'd5251,17'd5250,17'd4126,17'd4124,17'd59512,17'd52782,17'd58759,17'd52549,17'd59012,17'd52850,17'd53447,17'd54348,17'd69550,17'd54705,17'd68663,17'd68663,17'd55900,17'd65733,17'd57773,17'd65470,17'd55776,17'd64825,17'd55490,17'd63543,17'd57278,17'd58408,17'd65332,17'd64146,17'd60916,17'd64284,17'd69551,17'd55486,17'd67472,17'd59516,17'd69552,17'd69553,17'd69554,17'd69555,17'd69457,17'd69369,17'd69556,17'd69557,17'd69558,17'd69462,17'd69276,17'd69463,17'd69559,17'd69374,17'd69560,17'd69561,17'd69562,17'd69563,17'd60561,17'd69564,17'd62493,17'd69565,17'd69566,17'd69567,17'd17706,17'd69475,17'd15156,17'd15792,17'd69568,17'd69569,17'd69570,17'd52121,17'd69571,17'd8712,17'd69572,17'd69573,17'd8096,17'd18566,17'd12588,17'd19923,17'd8574,17'd8572,17'd12425,17'd24368,17'd32121,17'd59708,17'd14391,17'd69574,17'd55620,17'd69575,17'd69199,17'd53258,17'd132,17'd132,17'd134,17'd132,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd136,17'd136,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd11541,17'd20622,17'd20624,17'd69576,17'd69577,17'd52323,17'd69578,17'd51301,17'd53485,17'd42440,17'd34457,17'd39441,17'd32513,17'd29686,17'd23386,17'd23565,17'd23384,17'd29243,17'd29102,17'd23562,17'd34884,17'd29100,17'd28975,17'd23731,17'd24086,17'd30879,17'd28975,17'd28975,17'd28975,17'd28975,17'd28722,17'd30275,17'd23732,17'd23920,17'd30127,17'd23736,17'd30579,17'd29829,17'd29974,17'd45165,17'd57195,17'd22328,17'd45492,17'd44944,17'd48712,17'd49487,17'd34110,17'd59726,17'd53416,17'd21527,17'd52594,17'd69579,17'd69580,17'd69581,17'd69582,17'd69583,17'd69584,17'd69585,17'd69586,17'd69587,17'd17645,17'd67268,17'd69588,17'd69216,17'd68717,17'd69589,17'd69500,17'd69590,17'd69591,17'd69592,17'd69593,17'd69593,17'd69594,17'd69595,17'd69596,17'd69597,17'd10771,17'd8297,17'd9079,17'd15209,17'd69598,17'd10202,17'd11694,17'd17641,17'd69599,17'd69600,17'd69601,17'd7496,17'd10235,17'd11850,17'd69028,17'd69128,17'd11430,17'd10777,17'd10777,17'd10514,17'd9933,17'd68622,17'd69511,17'd69512,17'd69513,17'd69602,17'd69603,17'd69604,17'd69515,17'd69605,17'd69517,17'd69606,17'd69607,17'd69608,17'd69236,17'd69519,17'd67548,17'd65551,17'd69417,17'd69609,17'd69418,17'd65163,17'd68058,17'd69610,17'd64242,17'd66676,17'd66072,17'd66437,17'd66437,17'd65569,17'd65570,17'd65703,17'd65703,17'd65703,17'd67423,17'd67923,17'd68059,17'd69523,17'd69524,17'd68182,17'd68182,17'd69525,17'd69525,17'd68944,17'd69337,17'd69337,17'd69337,17'd69145,17'd69145,17'd69145,17'd69145,17'd69338,17'd69338,17'd69338,17'd69338,17'd69422,17'd69422,17'd69611,17'd69340,17'd63105,17'd63105,17'd63105,17'd63105,17'd63372,17'd63372,17'd68295,17'd68295,17'd63372,17'd63106,17'd63962,17'd69527,17'd68521,17'd64387,17'd69527,17'd66197,17'd65950,17'd62851,17'd17179,17'd14734,17'd67428,17'd62447,17'd62576,17'd62576,17'd67290,17'd62576,17'd67427,17'd16255,17'd65689,17'd65040,17'd69336,17'd68181,17'd68415,17'd66198,17'd64388,17'd69612,17'd69530,17'd69531,17'd64110,17'd65306,17'd64241,17'd64241,17'd64789,17'd64789,17'd67296,17'd68187,17'd69424,17'd68632,17'd69425,17'd69426,17'd66199,17'd67560,17'd63809,17'd63378,17'd62971,17'd62851,17'd64531,17'd62448,17'd67429,17'd69613,17'd39790,17'd10906,17'd3710,17'd6404,17'd54325,17'd69614,17'd38071,17'd1263,17'd604,17'd1668,17'd1111,17'd642,17'd408,17'd69615,17'd1682,17'd20867
},
'{
17'd69616,17'd6263,17'd9959,17'd4736,17'd4244,17'd4892,17'd3427,17'd3251,17'd3252,17'd1831,17'd1689,17'd1689,17'd14,17'd15,17'd0,17'd14,17'd1689,17'd1688,17'd17917,17'd2422,17'd69617,17'd65712,17'd69618,17'd67684,17'd67939,17'd69619,17'd67940,17'd69620,17'd69433,17'd67944,17'd69621,17'd68754,17'd68197,17'd69620,17'd67940,17'd69350,17'd65960,17'd9417,17'd8664,17'd7547,17'd67306,17'd64668,17'd0,17'd806,17'd20,17'd21,17'd11,17'd19,17'd3905,17'd17,17'd1416,17'd2257,17'd1688,17'd1689,17'd3250,17'd2935,17'd37047,17'd3101,17'd3252,17'd3252,17'd2426,17'd2426,17'd2257,17'd1414,17'd17,17'd17,17'd17,17'd17,17'd289,17'd30,17'd30,17'd3255,17'd3254,17'd4249,17'd3756,17'd6278,17'd6746,17'd5972,17'd27592,17'd9817,17'd7390,17'd7390,17'd7390,17'd7227,17'd7391,17'd7562,17'd69622,17'd69623,17'd69624,17'd69625,17'd69626,17'd69627,17'd65853,17'd65744,17'd24979,17'd37591,17'd25514,17'd69628,17'd6943,17'd69549,17'd69549,17'd38219,17'd7920,17'd40269,17'd9706,17'd10698,17'd43467,17'd43467,17'd20436,17'd10698,17'd69629,17'd12683,17'd13096,17'd21190,17'd30059,17'd10946,17'd6304,17'd8692,17'd8376,17'd7421,17'd7095,17'd6934,17'd4290,17'd52029,17'd52284,17'd69630,17'd16030,17'd47972,17'd55483,17'd54093,17'd56446,17'd54993,17'd56020,17'd66830,17'd65328,17'd55776,17'd63845,17'd56446,17'd69631,17'd55485,17'd55490,17'd63543,17'd63689,17'd69632,17'd69633,17'd61441,17'd58768,17'd61190,17'd1319,17'd61187,17'd56580,17'd63542,17'd69634,17'd69635,17'd69636,17'd69637,17'd69638,17'd69639,17'd69640,17'd69641,17'd69642,17'd69643,17'd69644,17'd69645,17'd69646,17'd69647,17'd69648,17'd69649,17'd69650,17'd69651,17'd61081,17'd62492,17'd69652,17'd69566,17'd15028,17'd15155,17'd69653,17'd15279,17'd14496,17'd13618,17'd19145,17'd26026,17'd23506,17'd49312,17'd45928,17'd69654,17'd69655,17'd35645,17'd8580,17'd9745,17'd21208,17'd12865,17'd8573,17'd30672,17'd23341,17'd19923,17'd59321,17'd63319,17'd69574,17'd7634,17'd69656,17'd23696,17'd13901,17'd5593,17'd5593,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd132,17'd132,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd131,17'd11541,17'd51987,17'd20764,17'd51806,17'd69657,17'd69658,17'd69659,17'd69660,17'd69661,17'd69662,17'd69663,17'd35157,17'd44702,17'd35455,17'd30882,17'd30730,17'd23384,17'd24902,17'd30879,17'd23731,17'd24086,17'd23732,17'd23564,17'd23564,17'd30275,17'd28722,17'd30879,17'd23731,17'd23917,17'd24087,17'd24087,17'd23920,17'd29099,17'd29827,17'd23923,17'd30128,17'd23215,17'd23389,17'd55132,17'd22674,17'd22008,17'd31192,17'd50577,17'd69664,17'd41584,17'd69665,17'd69666,17'd68685,17'd69667,17'd51810,17'd69668,17'd69669,17'd69670,17'd69671,17'd69672,17'd69673,17'd69674,17'd69675,17'd29858,17'd69676,17'd69677,17'd69678,17'd69679,17'd69680,17'd69499,17'd68718,17'd68814,17'd69681,17'd69682,17'd69683,17'd69684,17'd69685,17'd69686,17'd8924,17'd69687,17'd8620,17'd9231,17'd69688,17'd12889,17'd15971,17'd17510,17'd15839,17'd67652,17'd25621,17'd69689,17'd12885,17'd69690,17'd11850,17'd12301,17'd69028,17'd69691,17'd11430,17'd10641,17'd27932,17'd10515,17'd69692,17'd68825,17'd69029,17'd69512,17'd69602,17'd69693,17'd69694,17'd69515,17'd69695,17'd69696,17'd69697,17'd69698,17'd69699,17'd69700,17'd68052,17'd69519,17'd66786,17'd69701,17'd69701,17'd63939,17'd69702,17'd67918,17'd67792,17'd67423,17'd69703,17'd69144,17'd68060,17'd66677,17'd65570,17'd65570,17'd65570,17'd65570,17'd65703,17'd67423,17'd66677,17'd68060,17'd68059,17'd69523,17'd69704,17'd69523,17'd69523,17'd69705,17'd69706,17'd68519,17'd68944,17'd68945,17'd68833,17'd68833,17'd68945,17'd68945,17'd68945,17'd69145,17'd69145,17'd69707,17'd69708,17'd68520,17'd68521,17'd69340,17'd69709,17'd63105,17'd62969,17'd63372,17'd63372,17'd68295,17'd68295,17'd63106,17'd63962,17'd63962,17'd63962,17'd63962,17'd63962,17'd63807,17'd63807,17'd66197,17'd65308,17'd64390,17'd17179,17'd62576,17'd67289,17'd67291,17'd67291,17'd14583,17'd14583,17'd14734,17'd14976,17'd15734,17'd65816,17'd65688,17'd67287,17'd68740,17'd69710,17'd67800,17'd67932,17'd63511,17'd69531,17'd67793,17'd67793,17'd64110,17'd64241,17'd64241,17'd67436,17'd64789,17'd69711,17'd68298,17'd69147,17'd69147,17'd68947,17'd68633,17'd68633,17'd67295,17'd67295,17'd66929,17'd68297,17'd64527,17'd69712,17'd62851,17'd62698,17'd67925,17'd69713,17'd69714,17'd10906,17'd69715,17'd53293,17'd2391,17'd5195,17'd1262,17'd1666,17'd26595,17'd191,17'd644,17'd259,17'd69716,17'd69717,17'd595,17'd22100
},
'{
17'd69616,17'd5198,17'd5377,17'd69718,17'd4427,17'd4244,17'd3901,17'd3427,17'd2935,17'd2422,17'd1689,17'd1689,17'd14,17'd15,17'd2,17'd1127,17'd1689,17'd1688,17'd17917,17'd1831,17'd69719,17'd63976,17'd66808,17'd67810,17'd66207,17'd66440,17'd69254,17'd69720,17'd66939,17'd68852,17'd68529,17'd68641,17'd68530,17'd69435,17'd68962,17'd69721,17'd66088,17'd69722,17'd9417,17'd9546,17'd6894,17'd69723,17'd3249,17'd3,17'd25,17'd2598,17'd10,17'd11,17'd18,17'd18,17'd17,17'd2257,17'd1688,17'd1688,17'd3250,17'd2935,17'd34512,17'd3251,17'd14070,17'd3252,17'd2426,17'd2258,17'd2257,17'd1415,17'd17,17'd17,17'd17,17'd17,17'd289,17'd289,17'd30,17'd30,17'd3255,17'd3255,17'd3756,17'd11210,17'd11889,17'd6746,17'd27592,17'd10672,17'd7227,17'd7390,17'd7390,17'd7227,17'd69724,17'd10409,17'd11891,17'd69725,17'd69726,17'd69727,17'd69728,17'd69729,17'd69730,17'd69731,17'd8385,17'd69732,17'd69732,17'd25126,17'd69359,17'd69733,17'd69734,17'd69733,17'd25804,17'd8384,17'd24523,17'd9580,17'd69735,17'd69735,17'd69735,17'd9988,17'd12537,17'd12683,17'd12818,17'd12817,17'd10287,17'd10117,17'd10114,17'd8846,17'd7422,17'd7099,17'd7097,17'd7584,17'd6629,17'd4128,17'd4770,17'd65466,17'd66347,17'd47864,17'd57120,17'd57013,17'd48932,17'd58400,17'd59646,17'd57126,17'd59515,17'd59515,17'd55775,17'd54993,17'd68664,17'd68665,17'd55093,17'd56689,17'd63406,17'd55582,17'd57647,17'd57275,17'd58893,17'd57391,17'd60176,17'd58653,17'd63403,17'd69736,17'd69737,17'd69738,17'd69739,17'd69740,17'd69741,17'd69639,17'd69742,17'd69641,17'd69743,17'd69744,17'd69279,17'd69745,17'd69746,17'd69747,17'd69748,17'd69749,17'd69750,17'd60814,17'd69751,17'd62611,17'd69752,17'd69753,17'd15028,17'd15155,17'd16185,17'd16420,17'd13861,17'd13110,17'd11099,17'd24982,17'd9716,17'd69754,17'd69755,17'd69756,17'd69757,17'd17730,17'd17353,17'd69758,17'd8249,17'd24043,17'd8414,17'd8575,17'd30672,17'd8418,17'd58316,17'd63451,17'd69759,17'd66603,17'd69760,17'd65240,17'd11152,17'd5593,17'd5593,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd20466,17'd69761,17'd69762,17'd69763,17'd52420,17'd20919,17'd69764,17'd69765,17'd69766,17'd52594,17'd42602,17'd22510,17'd31345,17'd45986,17'd33944,17'd23572,17'd23217,17'd30128,17'd29530,17'd35865,17'd23387,17'd30128,17'd23923,17'd23923,17'd29827,17'd23566,17'd34137,17'd23918,17'd23920,17'd29241,17'd29241,17'd31502,17'd23923,17'd23217,17'd22679,17'd22678,17'd32344,17'd22162,17'd22335,17'd22684,17'd50818,17'd34879,17'd69767,17'd69768,17'd51067,17'd54139,17'd54214,17'd69769,17'd69770,17'd69771,17'd69772,17'd69773,17'd22022,17'd69774,17'd69775,17'd69776,17'd30615,17'd69777,17'd69778,17'd69779,17'd69780,17'd69781,17'd69679,17'd69680,17'd69499,17'd17157,17'd68921,17'd69782,17'd69783,17'd69783,17'd69784,17'd69685,17'd69785,17'd8620,17'd69786,17'd8624,17'd8462,17'd69688,17'd12745,17'd15971,17'd17510,17'd8764,17'd14710,17'd25621,17'd21302,17'd8454,17'd7666,17'd11850,17'd12301,17'd69028,17'd69691,17'd69691,17'd69787,17'd27932,17'd27933,17'd69692,17'd68825,17'd69029,17'd69512,17'd69602,17'd69788,17'd69789,17'd69515,17'd69329,17'd69790,17'd69790,17'd69791,17'd69698,17'd69792,17'd69793,17'd69035,17'd66786,17'd69794,17'd69794,17'd69795,17'd67035,17'd67919,17'd65570,17'd68059,17'd69796,17'd69144,17'd68060,17'd66677,17'd65570,17'd64109,17'd63965,17'd65703,17'd65703,17'd67423,17'd68060,17'd68182,17'd68059,17'd69523,17'd69797,17'd69523,17'd69798,17'd69706,17'd69706,17'd68944,17'd68944,17'd68945,17'd68833,17'd68833,17'd68833,17'd68833,17'd68833,17'd69338,17'd69338,17'd69799,17'd69799,17'd68521,17'd63807,17'd63373,17'd63242,17'd63372,17'd63372,17'd63372,17'd63106,17'd68295,17'd68295,17'd63106,17'd63106,17'd63962,17'd63962,17'd63962,17'd63962,17'd63807,17'd63243,17'd65308,17'd65441,17'd17415,17'd65705,17'd62976,17'd67289,17'd67291,17'd14434,17'd67557,17'd14583,17'd14734,17'd65705,17'd68416,17'd68741,17'd64507,17'd65164,17'd68949,17'd69710,17'd67932,17'd68415,17'd69531,17'd69531,17'd67793,17'd64110,17'd66929,17'd67436,17'd67436,17'd64789,17'd69800,17'd67439,17'd69424,17'd69147,17'd68837,17'd69425,17'd68633,17'd68633,17'd67295,17'd67172,17'd69801,17'd67793,17'd63965,17'd63964,17'd62970,17'd67554,17'd64788,17'd66195,17'd60399,17'd11048,17'd58626,17'd4558,17'd3247,17'd1261,17'd4727,17'd3743,17'd26595,17'd191,17'd970,17'd259,17'd17787,17'd69802,17'd1097,17'd2112
},
'{
17'd69803,17'd10397,17'd5377,17'd9959,17'd4427,17'd4892,17'd3427,17'd3427,17'd2935,17'd2422,17'd1688,17'd1689,17'd1127,17'd14,17'd2,17'd1127,17'd1688,17'd1689,17'd2594,17'd1831,17'd69804,17'd64928,17'd66439,17'd67938,17'd66089,17'd66442,17'd69805,17'd67569,17'd67449,17'd67813,17'd68754,17'd68309,17'd68643,17'd69806,17'd69807,17'd67940,17'd67939,17'd69808,17'd69809,17'd9265,17'd6896,17'd10799,17'd10668,17'd1,17'd16389,17'd1128,17'd10,17'd11,17'd18,17'd18,17'd17,17'd22965,17'd4247,17'd1688,17'd3250,17'd2422,17'd3101,17'd3251,17'd14188,17'd3252,17'd2258,17'd2258,17'd2257,17'd1415,17'd1416,17'd17,17'd3905,17'd18,17'd29,17'd289,17'd809,17'd30,17'd3255,17'd3255,17'd3756,17'd6278,17'd5803,17'd5803,17'd26971,17'd10672,17'd9817,17'd6907,17'd69810,17'd7390,17'd7063,17'd7730,17'd12037,17'd69811,17'd69812,17'd69813,17'd69353,17'd69814,17'd69815,17'd15903,17'd64158,17'd36764,17'd37323,17'd69816,17'd63421,17'd69446,17'd63421,17'd69817,17'd38887,17'd8547,17'd9013,17'd9443,17'd24523,17'd24523,17'd24523,17'd9845,17'd22285,17'd12818,17'd13096,17'd11916,17'd10287,17'd10117,17'd68095,17'd9985,17'd8073,17'd8070,17'd42795,17'd7095,17'd6629,17'd4289,17'd59390,17'd59264,17'd68438,17'd53082,17'd69818,17'd58648,17'd66457,17'd54020,17'd66570,17'd65080,17'd66830,17'd57014,17'd65202,17'd54992,17'd54893,17'd64947,17'd55901,17'd60172,17'd56688,17'd55907,17'd55582,17'd55182,17'd58885,17'd63279,17'd69819,17'd68327,17'd63277,17'd69820,17'd69821,17'd69822,17'd69823,17'd69824,17'd69825,17'd69639,17'd69826,17'd69827,17'd69828,17'd69829,17'd69464,17'd69830,17'd69831,17'd69832,17'd69833,17'd69834,17'd69835,17'd60203,17'd69836,17'd69837,17'd69838,17'd69839,17'd15921,17'd15278,17'd15410,17'd15408,17'd13860,17'd12964,17'd69840,17'd54034,17'd69841,17'd69842,17'd69843,17'd69844,17'd49428,17'd14005,17'd18203,17'd33716,17'd7946,17'd53035,17'd8416,17'd23342,17'd11137,17'd53035,17'd22996,17'd10482,17'd54650,17'd69845,17'd69846,17'd10349,17'd7979,17'd131,17'd135,17'd130,17'd130,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd128,17'd132,17'd131,17'd20623,17'd52247,17'd52737,17'd69847,17'd20771,17'd69848,17'd69849,17'd21226,17'd69668,17'd69850,17'd47652,17'd51066,17'd42603,17'd22511,17'd33162,17'd21846,17'd23394,17'd22324,17'd22325,17'd33311,17'd22332,17'd22504,17'd22330,17'd36986,17'd23218,17'd23215,17'd29686,17'd23566,17'd29376,17'd23387,17'd23388,17'd22328,17'd22860,17'd34281,17'd69851,17'd47746,17'd35709,17'd47160,17'd50898,17'd69852,17'd52004,17'd46777,17'd54583,17'd51468,17'd52754,17'd69853,17'd69854,17'd69855,17'd69856,17'd69857,17'd69858,17'd69859,17'd69860,17'd69861,17'd69862,17'd69863,17'd22715,17'd69864,17'd69865,17'd69866,17'd69867,17'd69868,17'd69869,17'd68717,17'd69018,17'd69870,17'd69871,17'd69872,17'd69783,17'd69784,17'd69685,17'd69785,17'd69873,17'd8622,17'd9382,17'd69874,17'd69688,17'd12888,17'd14558,17'd69875,17'd8764,17'd14710,17'd69876,17'd20841,17'd8454,17'd7666,17'd11850,17'd68823,17'd68823,17'd11573,17'd11430,17'd27932,17'd10515,17'd68928,17'd69692,17'd68825,17'd69877,17'd69878,17'd69879,17'd69880,17'd69789,17'd69694,17'd69329,17'd69881,17'd69790,17'd69791,17'd69882,17'd69883,17'd69793,17'd69035,17'd66179,17'd69794,17'd64367,17'd64088,17'd69884,17'd68740,17'd65570,17'd68059,17'd69796,17'd69144,17'd68060,17'd67423,17'd65703,17'd65570,17'd65703,17'd68292,17'd67423,17'd67923,17'd67923,17'd68059,17'd68182,17'd68059,17'd69524,17'd69523,17'd69797,17'd69706,17'd69885,17'd68944,17'd69337,17'd68833,17'd68833,17'd68833,17'd68833,17'd68833,17'd68520,17'd68520,17'd69422,17'd69422,17'd69422,17'd69340,17'd63373,17'd63106,17'd63372,17'd63372,17'd63106,17'd63106,17'd63962,17'd63962,17'd63962,17'd63106,17'd63106,17'd63106,17'd63962,17'd63962,17'd63962,17'd65702,17'd66197,17'd65308,17'd62853,17'd65705,17'd62576,17'd67290,17'd67290,17'd14583,17'd67557,17'd15618,17'd14583,17'd14976,17'd15734,17'd65816,17'd68741,17'd65039,17'd69886,17'd69887,17'd69887,17'd68415,17'd69241,17'd69531,17'd69531,17'd64110,17'd65306,17'd67436,17'd67436,17'd64789,17'd65056,17'd67439,17'd69888,17'd69889,17'd69424,17'd67672,17'd69039,17'd66320,17'd67295,17'd65055,17'd64921,17'd64110,17'd65306,17'd64529,17'd66073,17'd63242,17'd62848,17'd67294,17'd17292,17'd38580,17'd38202,17'd5028,17'd12914,17'd4422,17'd3743,17'd1394,17'd604,17'd411,17'd1111,17'd970,17'd259,17'd41005,17'd69890,17'd258,17'd9942
},
'{
17'd69891,17'd6262,17'd5960,17'd5377,17'd4087,17'd4244,17'd3901,17'd3427,17'd3101,17'd2784,17'd3250,17'd1688,17'd1127,17'd14,17'd2,17'd1127,17'd1688,17'd1689,17'd4247,17'd1831,17'd6260,17'd69892,17'd64119,17'd67567,17'd66088,17'd66207,17'd69805,17'd69893,17'd68526,17'd67571,17'd68852,17'd68309,17'd69894,17'd68643,17'd68197,17'd66937,17'd66686,17'd69350,17'd65959,17'd69809,17'd8515,17'd6738,17'd9967,17'd63116,17'd1276,17'd11,17'd11,17'd808,17'd19,17'd18,17'd17,17'd22965,17'd4247,17'd1688,17'd3250,17'd3250,17'd2784,17'd3251,17'd38864,17'd3252,17'd2597,17'd2258,17'd2257,17'd1415,17'd1416,17'd17,17'd3905,17'd18,17'd29,17'd29,17'd809,17'd30,17'd3754,17'd3255,17'd3434,17'd3910,17'd5804,17'd5803,17'd27445,17'd10672,17'd7730,17'd9277,17'd69895,17'd7559,17'd6905,17'd9970,17'd69438,17'd69896,17'd69623,17'd69897,17'd69898,17'd69899,17'd69900,17'd69901,17'd65744,17'd35631,17'd37322,17'd69359,17'd63421,17'd69902,17'd63421,17'd69817,17'd25804,17'd8385,17'd28670,17'd9162,17'd66346,17'd66346,17'd69903,17'd24522,17'd12067,17'd13096,17'd12067,17'd10120,17'd24198,17'd9578,17'd29181,17'd68095,17'd9985,17'd65462,17'd69904,17'd67466,17'd68321,17'd62998,17'd62353,17'd59643,17'd3298,17'd3301,17'd58396,17'd69905,17'd53163,17'd54350,17'd54020,17'd65470,17'd59515,17'd65202,17'd60171,17'd55184,17'd60172,17'd55901,17'd69820,17'd69906,17'd60172,17'd54892,17'd63403,17'd55582,17'd61189,17'd57921,17'd57783,17'd55090,17'd69907,17'd69906,17'd69908,17'd69909,17'd69910,17'd69911,17'd69912,17'd69913,17'd69914,17'd69914,17'd69828,17'd69915,17'd69559,17'd69916,17'd69647,17'd69917,17'd69918,17'd69919,17'd69920,17'd69921,17'd69922,17'd69923,17'd69924,17'd69839,17'd15660,17'd15543,17'd16420,17'd69925,17'd69926,17'd19768,17'd22984,17'd51782,17'd69927,17'd69842,17'd69928,17'd69929,17'd69930,17'd69931,17'd11968,17'd17354,17'd9350,17'd7945,17'd8418,17'd15945,17'd8413,17'd8250,17'd9051,17'd12729,17'd69932,17'd69933,17'd69934,17'd10187,17'd53258,17'd131,17'd132,17'd129,17'd130,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd130,17'd130,17'd132,17'd131,17'd52069,17'd69935,17'd52737,17'd69936,17'd67993,17'd69937,17'd69938,17'd69939,17'd21235,17'd69940,17'd69941,17'd52593,17'd52681,17'd51911,17'd68686,17'd69942,17'd69943,17'd69944,17'd21851,17'd22013,17'd47358,17'd47358,17'd30880,17'd22861,17'd22158,17'd30426,17'd22677,17'd23038,17'd33311,17'd22333,17'd22861,17'd22336,17'd22002,17'd47160,17'd53569,17'd69945,17'd69946,17'd69947,17'd69948,17'd69949,17'd54214,17'd69950,17'd53991,17'd54848,17'd21231,17'd69951,17'd69952,17'd69953,17'd69954,17'd69955,17'd69956,17'd69957,17'd69958,17'd69959,17'd69960,17'd69961,17'd29716,17'd69962,17'd69963,17'd69867,17'd69964,17'd69589,17'd69965,17'd69018,17'd69966,17'd69872,17'd69783,17'd69783,17'd69967,17'd15837,17'd69968,17'd69687,17'd8772,17'd9382,17'd69874,17'd69688,17'd12447,17'd8916,17'd69875,17'd8764,17'd14846,17'd27691,17'd67411,17'd7993,17'd10235,17'd11850,17'd68823,17'd68927,17'd69691,17'd11430,17'd27932,17'd27932,17'd27933,17'd69692,17'd68825,17'd69129,17'd69969,17'd69970,17'd69971,17'd69788,17'd69694,17'd69516,17'd69881,17'd69972,17'd69697,17'd69973,17'd69974,17'd69975,17'd69976,17'd66305,17'd69794,17'd69977,17'd64226,17'd69334,17'd69610,17'd66677,17'd68059,17'd69524,17'd68059,17'd68060,17'd67423,17'd65703,17'd65703,17'd64529,17'd69978,17'd67423,17'd68060,17'd67923,17'd68059,17'd68182,17'd68182,17'd69144,17'd69523,17'd69523,17'd69706,17'd69706,17'd68944,17'd69337,17'd68520,17'd68521,17'd68520,17'd68520,17'd68520,17'd68520,17'd68520,17'd68520,17'd68521,17'd68521,17'd63373,17'd63373,17'd63106,17'd63106,17'd63106,17'd63962,17'd63962,17'd63962,17'd63962,17'd63962,17'd63106,17'd63106,17'd63962,17'd63962,17'd69527,17'd69527,17'd65702,17'd65308,17'd65441,17'd67426,17'd62576,17'd67290,17'd67290,17'd62576,17'd14583,17'd15618,17'd15618,17'd14734,17'd14976,17'd68416,17'd66791,17'd66536,17'd68290,17'd68949,17'd69710,17'd69887,17'd69241,17'd69979,17'd69531,17'd63511,17'd64110,17'd65306,17'd67436,17'd64789,17'd64789,17'd69711,17'd67931,17'd69980,17'd69889,17'd68632,17'd67673,17'd68633,17'd66320,17'd66320,17'd65055,17'd64921,17'd65307,17'd67920,17'd65570,17'd65181,17'd63807,17'd64526,17'd67433,17'd69981,17'd37958,17'd12773,17'd69982,17'd57610,17'd5372,17'd3743,17'd781,17'd604,17'd605,17'd605,17'd970,17'd259,17'd261,17'd47670,17'd271,17'd19493
},
'{
17'd29754,17'd6262,17'd5643,17'd5199,17'd4087,17'd3902,17'd4892,17'd6420,17'd3101,17'd2935,17'd2422,17'd1688,17'd1127,17'd14,17'd2,17'd466,17'd4247,17'd1689,17'd1689,17'd1688,17'd3250,17'd68191,17'd63817,17'd69249,17'd66692,17'd66208,17'd67446,17'd69983,17'd67303,17'd66940,17'd67690,17'd68196,17'd69252,17'd69984,17'd67690,17'd69349,17'd67940,17'd69985,17'd66089,17'd9675,17'd8515,17'd7053,17'd11735,17'd63257,17'd17187,17'd979,17'd1128,17'd25,17'd11,17'd18,17'd17,17'd1416,17'd4247,17'd1688,17'd3250,17'd2781,17'd3250,17'd14188,17'd38864,17'd3252,17'd2597,17'd2258,17'd2597,17'd1415,17'd1416,17'd3905,17'd3905,17'd18,17'd652,17'd652,17'd289,17'd289,17'd3755,17'd3595,17'd5209,17'd3910,17'd5804,17'd5803,17'd6746,17'd10408,17'd10672,17'd7228,17'd7559,17'd69986,17'd69987,17'd7064,17'd69988,17'd69989,17'd11892,17'd25115,17'd69990,17'd69991,17'd69992,17'd69993,17'd69994,17'd24979,17'd69816,17'd69359,17'd63421,17'd69995,17'd69996,17'd69997,17'd25804,17'd24979,17'd38218,17'd28670,17'd69998,17'd67702,17'd67702,17'd67465,17'd24198,17'd10120,17'd9845,17'd9705,17'd9579,17'd24522,17'd29181,17'd10115,17'd66105,17'd63834,17'd69999,17'd63535,17'd63134,17'd6477,17'd6775,17'd6315,17'd6150,17'd5841,17'd4771,17'd63139,17'd63139,17'd54094,17'd53880,17'd54093,17'd55775,17'd57126,17'd60171,17'd64419,17'd59516,17'd54892,17'd70000,17'd55901,17'd64000,17'd54803,17'd60299,17'd63141,17'd65207,17'd58159,17'd57782,17'd70001,17'd65739,17'd55185,17'd70002,17'd70003,17'd70004,17'd70005,17'd70006,17'd70007,17'd69914,17'd69914,17'd69828,17'd70008,17'd69374,17'd70009,17'd70010,17'd70011,17'd70012,17'd70013,17'd69470,17'd70014,17'd62893,17'd69924,17'd70015,17'd69839,17'd15790,17'd17218,17'd17705,17'd14786,17'd13983,17'd12225,17'd21196,17'd54640,17'd70016,17'd70017,17'd70018,17'd70019,17'd70020,17'd7615,17'd16802,17'd25152,17'd17129,17'd7784,17'd10608,17'd9196,17'd25147,17'd17128,17'd70021,17'd53981,17'd70022,17'd70023,17'd69934,17'd11540,17'd68231,17'd134,17'd130,17'd141,17'd130,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd128,17'd134,17'd131,17'd52245,17'd20627,17'd52883,17'd66484,17'd52812,17'd21222,17'd52496,17'd69938,17'd52059,17'd70024,17'd70025,17'd70026,17'd70027,17'd69302,17'd70028,17'd21526,17'd54296,17'd21999,17'd51726,17'd46678,17'd51164,17'd46571,17'd42305,17'd41584,17'd50740,17'd33646,17'd41728,17'd33160,17'd33314,17'd70029,17'd51543,17'd46455,17'd46860,17'd70030,17'd70031,17'd70032,17'd70033,17'd68579,17'd21382,17'd70034,17'd21234,17'd70035,17'd66730,17'd21522,17'd69849,17'd52496,17'd70036,17'd70037,17'd70038,17'd70039,17'd70040,17'd70041,17'd70042,17'd70043,17'd70044,17'd26804,17'd70045,17'd68497,17'd68917,17'd70046,17'd70047,17'd69402,17'd70048,17'd70049,17'd70050,17'd69683,17'd70051,17'd69967,17'd15838,17'd70052,17'd8622,17'd70053,17'd9382,17'd8623,17'd69688,17'd69598,17'd11987,17'd10201,17'd8614,17'd14415,17'd69689,17'd11986,17'd7993,17'd10235,17'd11850,17'd68823,17'd11573,17'd11430,17'd11430,17'd27932,17'd10515,17'd68928,17'd69692,17'd68825,17'd69877,17'd70054,17'd69879,17'd69880,17'd69788,17'd69693,17'd69516,17'd70055,17'd69790,17'd69697,17'd69882,17'd70056,17'd69975,17'd70057,17'd66061,17'd69701,17'd64226,17'd66064,17'd66663,17'd63966,17'd66072,17'd68059,17'd69524,17'd68059,17'd67923,17'd68292,17'd67423,17'd67553,17'd70058,17'd70059,17'd68293,17'd70060,17'd70060,17'd68059,17'd68182,17'd68182,17'd69144,17'd69523,17'd69523,17'd68518,17'd68518,17'd70061,17'd69338,17'd69611,17'd70062,17'd64386,17'd64386,17'd64386,17'd64526,17'd63962,17'd63962,17'd63962,17'd63962,17'd63106,17'd63106,17'd63106,17'd63106,17'd63106,17'd63962,17'd63962,17'd69527,17'd63962,17'd63962,17'd63962,17'd63962,17'd63807,17'd64387,17'd64387,17'd67924,17'd65308,17'd64390,17'd65571,17'd69342,17'd67290,17'd67290,17'd14583,17'd67557,17'd14583,17'd67557,17'd69342,17'd69342,17'd65705,17'd68416,17'd70063,17'd64507,17'd68740,17'd69887,17'd67932,17'd68415,17'd67422,17'd67422,17'd63377,17'd63658,17'd63657,17'd63809,17'd64921,17'd64921,17'd67295,17'd67296,17'd70064,17'd70065,17'd69424,17'd67673,17'd66320,17'd66320,17'd65831,17'd65831,17'd65056,17'd65056,17'd70066,17'd70067,17'd66677,17'd68061,17'd68520,17'd70068,17'd67048,17'd15484,17'd37959,17'd70069,17'd10257,17'd7211,17'd5371,17'd604,17'd604,17'd1111,17'd643,17'd643,17'd643,17'd206,17'd3746,17'd3746,17'd643,17'd3900
},
'{
17'd7369,17'd7369,17'd5375,17'd5644,17'd5201,17'd4087,17'd3902,17'd4428,17'd3427,17'd2935,17'd2784,17'd2422,17'd1688,17'd14,17'd2,17'd1127,17'd1689,17'd1689,17'd1689,17'd1688,17'd1688,17'd2592,17'd66090,17'd70070,17'd65843,17'd70071,17'd66329,17'd69983,17'd69251,17'd69720,17'd67572,17'd68643,17'd70072,17'd68080,17'd70073,17'd70074,17'd68644,17'd70075,17'd66208,17'd69722,17'd65845,17'd7378,17'd7890,17'd70076,17'd9969,17'd5969,17'd1128,17'd25,17'd10,17'd11,17'd18,17'd17,17'd1127,17'd4247,17'd1688,17'd2781,17'd2781,17'd3252,17'd14188,17'd14070,17'd2258,17'd2597,17'd2597,17'd1414,17'd1416,17'd3905,17'd3905,17'd18,17'd652,17'd652,17'd29,17'd29,17'd3755,17'd3433,17'd5209,17'd5208,17'd3910,17'd5804,17'd6746,17'd70077,17'd11345,17'd9817,17'd7559,17'd7896,17'd69986,17'd7559,17'd7391,17'd69438,17'd5662,17'd5815,17'd70078,17'd70079,17'd70080,17'd70081,17'd46797,17'd70082,17'd70083,17'd70084,17'd63421,17'd69996,17'd70085,17'd70086,17'd37322,17'd36923,17'd24979,17'd8222,17'd69358,17'd68434,17'd70087,17'd67702,17'd67465,17'd24522,17'd9579,17'd9579,17'd9579,17'd24522,17'd24522,17'd29181,17'd68435,17'd50192,17'd63839,17'd63840,17'd64943,17'd6476,17'd42060,17'd6319,17'd43602,17'd64416,17'd3296,17'd3302,17'd3635,17'd59141,17'd53812,17'd68973,17'd54253,17'd55775,17'd59515,17'd64419,17'd68097,17'd64553,17'd59516,17'd58522,17'd70000,17'd70088,17'd70089,17'd54703,17'd55779,17'd55582,17'd56023,17'd69070,17'd55181,17'd54893,17'd70090,17'd70091,17'd70092,17'd70093,17'd70094,17'd70095,17'd70096,17'd70097,17'd70098,17'd70099,17'd70100,17'd70101,17'd70102,17'd70103,17'd70104,17'd70105,17'd60328,17'd70106,17'd70107,17'd69924,17'd70015,17'd70108,17'd15790,17'd17218,17'd70109,17'd70110,17'd13339,17'd10705,17'd55407,17'd50300,17'd49722,17'd70111,17'd70112,17'd70113,17'd70114,17'd70115,17'd14681,17'd14937,17'd15192,17'd17129,17'd14527,17'd8417,17'd19923,17'd9197,17'd70116,17'd9353,17'd70117,17'd70118,17'd70119,17'd70120,17'd21679,17'd720,17'd136,17'd138,17'd130,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd132,17'd131,17'd131,17'd52245,17'd52069,17'd65124,17'd67992,17'd65362,17'd70121,17'd22844,17'd21682,17'd70122,17'd70123,17'd52496,17'd70124,17'd70125,17'd70126,17'd70127,17'd21394,17'd70128,17'd55049,17'd70129,17'd70130,17'd51384,17'd21387,17'd21384,17'd52964,17'd47161,17'd47161,17'd52160,17'd51922,17'd52160,17'd47161,17'd21705,17'd51980,17'd21537,17'd53492,17'd21524,17'd70131,17'd70132,17'd70133,17'd70134,17'd70135,17'd70136,17'd70137,17'd70138,17'd70139,17'd68892,17'd68467,17'd51972,17'd70140,17'd70141,17'd70142,17'd70143,17'd70144,17'd70145,17'd70146,17'd70147,17'd68269,17'd70148,17'd68810,17'd70046,17'd70047,17'd70048,17'd69870,17'd70149,17'd70050,17'd69683,17'd70051,17'd70150,17'd70151,17'd69687,17'd9080,17'd70053,17'd9382,17'd8623,17'd69874,17'd69598,17'd11987,17'd11016,17'd8614,17'd14297,17'd70152,17'd11551,17'd7173,17'd10235,17'd68926,17'd68927,17'd11573,17'd11430,17'd11430,17'd27932,17'd27932,17'd27933,17'd69692,17'd68825,17'd69129,17'd69969,17'd70153,17'd70154,17'd69788,17'd69693,17'd70155,17'd70055,17'd70156,17'd70157,17'd70158,17'd70159,17'd70160,17'd70161,17'd66304,17'd69701,17'd67037,17'd64507,17'd63378,17'd67671,17'd66928,17'd68059,17'd68059,17'd67923,17'd67923,17'd68292,17'd67423,17'd67921,17'd70162,17'd70162,17'd70163,17'd70164,17'd70164,17'd68059,17'd68182,17'd68059,17'd68059,17'd69523,17'd69523,17'd68518,17'd68518,17'd70165,17'd69338,17'd69611,17'd70062,17'd63241,17'd63105,17'd63105,17'd63372,17'd63106,17'd63106,17'd63962,17'd63962,17'd63106,17'd63106,17'd63106,17'd63962,17'd63962,17'd63962,17'd63962,17'd69527,17'd63962,17'd63962,17'd63962,17'd63962,17'd64387,17'd64387,17'd64387,17'd66435,17'd65441,17'd65571,17'd67426,17'd14734,17'd67290,17'd67290,17'd14583,17'd67557,17'd67557,17'd69342,17'd69342,17'd62701,17'd69240,17'd70166,17'd66306,17'd66535,17'd68181,17'd69887,17'd67932,17'd69241,17'd67422,17'd67422,17'd63377,17'd64528,17'd63657,17'd63809,17'd64921,17'd64921,17'd66320,17'd68187,17'd70167,17'd70167,17'd67672,17'd69039,17'd66320,17'd66320,17'd66077,17'd65831,17'd69800,17'd65056,17'd70067,17'd70168,17'd67923,17'd66319,17'd69338,17'd67044,17'd66070,17'd7364,17'd70169,17'd70170,17'd70171,17'd5940,17'd11337,17'd192,17'd191,17'd605,17'd206,17'd206,17'd643,17'd2779,17'd3746,17'd206,17'd1687,17'd1550
},
'{
17'd7883,17'd7369,17'd5375,17'd5790,17'd5201,17'd4426,17'd3902,17'd4892,17'd3427,17'd3101,17'd2784,17'd2422,17'd1688,17'd1127,17'd2,17'd466,17'd1127,17'd1689,17'd3250,17'd1689,17'd4247,17'd1831,17'd13186,17'd64122,17'd67062,17'd68638,17'd70071,17'd66555,17'd70172,17'd67940,17'd69620,17'd67572,17'd69252,17'd70173,17'd69984,17'd70174,17'd69620,17'd67940,17'd67939,17'd70175,17'd70176,17'd9963,17'd70177,17'd70178,17'd65584,17'd14442,17'd19,17'd10,17'd10,17'd11,17'd18,17'd16,17'd14,17'd4247,17'd1688,17'd1689,17'd2781,17'd2422,17'd14070,17'd14070,17'd52621,17'd3752,17'd2596,17'd1414,17'd17,17'd3905,17'd20404,17'd1128,17'd1128,17'd1128,17'd652,17'd652,17'd4091,17'd3908,17'd3433,17'd5208,17'd3910,17'd6278,17'd11889,17'd11211,17'd6279,17'd7730,17'd6905,17'd7729,17'd69986,17'd69895,17'd7560,17'd10409,17'd6281,17'd5062,17'd70179,17'd70180,17'd70181,17'd70182,17'd70183,17'd70184,17'd70185,17'd69628,17'd70084,17'd69359,17'd37975,17'd37975,17'd37974,17'd37322,17'd69816,17'd38887,17'd70082,17'd65744,17'd70087,17'd8544,17'd8695,17'd8695,17'd9306,17'd9306,17'd9578,17'd24522,17'd24198,17'd30059,17'd10117,17'd10946,17'd49201,17'd64275,17'd64680,17'd67587,17'd6478,17'd6319,17'd6320,17'd42797,17'd62224,17'd62354,17'd2982,17'd2989,17'd61436,17'd60652,17'd70186,17'd66349,17'd65470,17'd59515,17'd64682,17'd64553,17'd60539,17'd57128,17'd70187,17'd70188,17'd60540,17'd55907,17'd56582,17'd60656,17'd67472,17'd70189,17'd64283,17'd70190,17'd70191,17'd70192,17'd70193,17'd70194,17'd70195,17'd70196,17'd70096,17'd70197,17'd70198,17'd70199,17'd70200,17'd70201,17'd69917,17'd70202,17'd70203,17'd70204,17'd60446,17'd70205,17'd70107,17'd70206,17'd70015,17'd70108,17'd15790,17'd17218,17'd14786,17'd14644,17'd14234,17'd26025,17'd53532,17'd28444,17'd70207,17'd47581,17'd70208,17'd70209,17'd70210,17'd70211,17'd7790,17'd25005,17'd7617,17'd7787,17'd7947,17'd16072,17'd10028,17'd23688,17'd70212,17'd70213,17'd70214,17'd70215,17'd70216,17'd70120,17'd16811,17'd70217,17'd136,17'd138,17'd130,17'd128,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd131,17'd131,17'd131,17'd132,17'd128,17'd130,17'd130,17'd130,17'd132,17'd11541,17'd11541,17'd11541,17'd131,17'd11541,17'd20625,17'd69935,17'd69200,17'd20767,17'd70218,17'd70219,17'd52661,17'd52578,17'd69577,17'd70220,17'd51535,17'd53640,17'd70221,17'd70222,17'd70223,17'd70224,17'd70225,17'd51808,17'd68894,17'd70226,17'd70227,17'd70228,17'd21383,17'd53207,17'd51991,17'd53493,17'd52326,17'd70229,17'd54848,17'd70230,17'd52814,17'd70231,17'd70232,17'd70233,17'd68893,17'd70234,17'd70235,17'd70236,17'd21681,17'd70237,17'd67992,17'd67992,17'd70238,17'd70239,17'd70240,17'd70241,17'd35323,17'd70242,17'd70243,17'd70244,17'd70245,17'd69498,17'd68916,17'd69118,17'd70046,17'd70047,17'd70048,17'd70246,17'd70149,17'd70050,17'd69593,17'd70247,17'd70150,17'd15590,17'd69687,17'd9080,17'd9515,17'd9382,17'd8623,17'd8462,17'd12283,17'd11987,17'd70248,17'd8614,17'd14297,17'd70249,17'd9639,17'd7495,17'd6551,17'd68621,17'd68927,17'd11573,17'd11430,17'd11315,17'd27932,17'd10515,17'd68928,17'd69692,17'd68825,17'd70250,17'd70251,17'd70252,17'd70253,17'd69788,17'd69971,17'd70155,17'd70254,17'd70255,17'd70256,17'd70257,17'd70159,17'd69235,17'd70258,17'd66060,17'd69701,17'd64227,17'd66790,17'd66435,17'd70259,17'd68519,17'd68518,17'd68518,17'd68060,17'd67923,17'd68517,17'd67923,17'd68293,17'd70260,17'd70261,17'd70262,17'd70262,17'd70263,17'd70264,17'd70264,17'd70060,17'd70060,17'd69523,17'd69523,17'd68518,17'd68519,17'd70061,17'd69145,17'd67045,17'd67044,17'd63105,17'd63105,17'd63372,17'd63106,17'd63106,17'd65950,17'd65950,17'd66197,17'd63106,17'd63106,17'd63106,17'd63962,17'd63807,17'd64387,17'd64387,17'd64387,17'd64387,17'd64387,17'd64387,17'd64387,17'd64387,17'd64387,17'd63963,17'd65702,17'd65571,17'd15734,17'd62449,17'd62576,17'd14583,17'd14583,17'd67557,17'd67557,17'd67426,17'd69342,17'd14976,17'd68836,17'd65816,17'd65040,17'd70265,17'd70266,17'd68181,17'd69887,17'd68415,17'd69241,17'd67792,17'd67792,17'd63658,17'd64528,17'd63809,17'd63809,17'd64921,17'd65831,17'd67439,17'd70167,17'd69424,17'd68632,17'd69039,17'd66076,17'd66320,17'd67296,17'd70267,17'd69800,17'd70268,17'd70268,17'd70269,17'd70168,17'd68517,17'd68519,17'd70270,17'd66193,17'd70271,17'd70272,17'd70273,17'd70274,17'd5183,17'd8185,17'd11337,17'd192,17'd1667,17'd1243,17'd271,17'd207,17'd272,17'd269,17'd70275,17'd1124,17'd70276,17'd14316
},
'{
17'd8509,17'd7883,17'd7046,17'd5790,17'd5376,17'd5201,17'd4087,17'd4244,17'd3901,17'd2934,17'd2593,17'd2784,17'd3250,17'd1689,17'd14,17'd1127,17'd1967,17'd3250,17'd3250,17'd1689,17'd4247,17'd17917,17'd70277,17'd70278,17'd65839,17'd67938,17'd66208,17'd67939,17'd70279,17'd70280,17'd70281,17'd66939,17'd69434,17'd69054,17'd70282,17'd70283,17'd69349,17'd67688,17'd70284,17'd66332,17'd70285,17'd69156,17'd70286,17'd6591,17'd70287,17'd17187,17'd979,17'd1128,17'd10,17'd11,17'd18,17'd18,17'd2,17'd4247,17'd1688,17'd1689,17'd2781,17'd3250,17'd3252,17'd14070,17'd10547,17'd3752,17'd2596,17'd1414,17'd17,17'd3905,17'd20404,17'd20404,17'd1128,17'd1128,17'd652,17'd28,17'd4431,17'd3908,17'd3433,17'd3595,17'd3910,17'd3910,17'd5804,17'd68646,17'd6279,17'd10672,17'd6747,17'd70288,17'd7896,17'd69895,17'd7390,17'd6747,17'd7063,17'd5522,17'd70289,17'd70290,17'd70291,17'd70292,17'd70293,17'd46365,17'd70294,17'd69628,17'd69628,17'd6943,17'd37974,17'd38096,17'd37970,17'd38095,17'd69360,17'd70295,17'd39054,17'd69263,17'd28206,17'd8384,17'd8849,17'd8849,17'd9161,17'd9306,17'd9578,17'd9578,17'd24522,17'd10118,17'd10117,17'd10431,17'd10114,17'd9985,17'd70296,17'd65325,17'd6637,17'd6632,17'd44281,17'd6311,17'd43201,17'd70297,17'd60532,17'd2825,17'd2990,17'd3959,17'd70298,17'd69552,17'd70299,17'd54705,17'd60172,17'd56689,17'd69907,17'd70300,17'd56911,17'd70301,17'd70302,17'd56352,17'd70303,17'd62876,17'd55282,17'd63544,17'd54803,17'd70304,17'd70305,17'd70192,17'd70306,17'd70307,17'd70308,17'd70309,17'd70310,17'd70197,17'd70198,17'd70311,17'd70312,17'd70313,17'd70011,17'd70314,17'd70315,17'd70316,17'd59814,17'd70317,17'd70318,17'd70206,17'd70319,17'd70108,17'd15790,17'd15277,17'd15277,17'd70320,17'd70321,17'd10133,17'd51952,17'd70322,17'd70323,17'd70324,17'd70325,17'd70326,17'd37849,17'd70327,17'd9623,17'd13377,17'd14680,17'd14385,17'd17482,17'd53836,17'd17850,17'd70328,17'd70329,17'd70330,17'd70331,17'd70332,17'd70216,17'd9494,17'd9360,17'd70217,17'd136,17'd138,17'd130,17'd128,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd132,17'd130,17'd130,17'd128,17'd132,17'd132,17'd132,17'd132,17'd128,17'd130,17'd131,17'd20623,17'd20625,17'd22665,17'd24056,17'd52884,17'd66125,17'd70333,17'd70334,17'd70121,17'd22844,17'd68353,17'd70335,17'd70336,17'd68232,17'd70337,17'd70338,17'd51822,17'd70339,17'd70225,17'd70340,17'd70341,17'd70342,17'd21391,17'd70343,17'd66862,17'd67361,17'd70344,17'd21380,17'd70025,17'd70345,17'd70346,17'd67232,17'd68353,17'd70347,17'd70348,17'd65771,17'd20465,17'd131,17'd11541,17'd133,17'd131,17'd70349,17'd70350,17'd70351,17'd70352,17'd38302,17'd70353,17'd70354,17'd70355,17'd18107,17'd70356,17'd70357,17'd70358,17'd70359,17'd69591,17'd70360,17'd70246,17'd70149,17'd69593,17'd69784,17'd70247,17'd70361,17'd70362,17'd8622,17'd9080,17'd9515,17'd9382,17'd8624,17'd8462,17'd12283,17'd11987,17'd70248,17'd14958,17'd14297,17'd70363,17'd9220,17'd7666,17'd11850,17'd68823,17'd11573,17'd11573,17'd11430,17'd69787,17'd27932,17'd27932,17'd27933,17'd69692,17'd68825,17'd70364,17'd69412,17'd70153,17'd70154,17'd69788,17'd69971,17'd70154,17'd70365,17'd70255,17'd70366,17'd70367,17'd70368,17'd69235,17'd70369,17'd70370,17'd69794,17'd65289,17'd62971,17'd68833,17'd68518,17'd68519,17'd68518,17'd68518,17'd68060,17'd67923,17'd68517,17'd67923,17'd70164,17'd70260,17'd70371,17'd70372,17'd70371,17'd70263,17'd70264,17'd70263,17'd70164,17'd70060,17'd69524,17'd69523,17'd68519,17'd68944,17'd69145,17'd69145,17'd69338,17'd69339,17'd64526,17'd64526,17'd63962,17'd63962,17'd66197,17'd66197,17'd66197,17'd66197,17'd63372,17'd63106,17'd63106,17'd63962,17'd63807,17'd64387,17'd64387,17'd64387,17'd64387,17'd64919,17'd64919,17'd64919,17'd64919,17'd64387,17'd63243,17'd65308,17'd65571,17'd65705,17'd62576,17'd62576,17'd14583,17'd67557,17'd67557,17'd69342,17'd17179,17'd62975,17'd62975,17'd70373,17'd66306,17'd64507,17'd70374,17'd70375,17'd70376,17'd68949,17'd69241,17'd69241,17'd67792,17'd69610,17'd64528,17'd63657,17'd63809,17'd64921,17'd65055,17'd66320,17'd68298,17'd70065,17'd70377,17'd68947,17'd69039,17'd66076,17'd67296,17'd67439,17'd70267,17'd69800,17'd70268,17'd70268,17'd70269,17'd70378,17'd70379,17'd69704,17'd69706,17'd70380,17'd65943,17'd70381,17'd70382,17'd12923,17'd49009,17'd70383,17'd11337,17'd604,17'd1823,17'd1243,17'd271,17'd271,17'd641,17'd2779,17'd3747,17'd972,17'd70276,17'd14316
},
'{
17'd8509,17'd7046,17'd6262,17'd5643,17'd5377,17'd5201,17'd5646,17'd4244,17'd3592,17'd2934,17'd2593,17'd2935,17'd2422,17'd1689,17'd14,17'd1127,17'd1689,17'd3750,17'd2781,17'd3250,17'd4247,17'd2594,17'd1688,17'd12652,17'd64537,17'd70384,17'd66327,17'd69350,17'd66326,17'd66936,17'd69436,17'd69720,17'd68528,17'd69434,17'd70385,17'd70283,17'd69435,17'd68427,17'd69619,17'd68964,17'd70386,17'd68853,17'd70387,17'd7051,17'd63520,17'd63118,17'd17,17'd19,17'd1128,17'd10,17'd19,17'd18,17'd2,17'd2595,17'd2594,17'd1127,17'd1688,17'd1967,17'd2781,17'd14070,17'd12195,17'd3429,17'd2596,17'd2257,17'd17,17'd3905,17'd1128,17'd11,17'd11,17'd11,17'd27,17'd28,17'd29,17'd289,17'd3595,17'd3433,17'd5208,17'd3910,17'd6278,17'd11889,17'd11737,17'd6279,17'd6904,17'd8048,17'd70388,17'd70388,17'd6906,17'd6601,17'd7388,17'd70389,17'd70390,17'd70391,17'd70392,17'd70393,17'd70394,17'd70395,17'd70396,17'd25126,17'd25126,17'd36194,17'd37723,17'd37974,17'd37973,17'd38222,17'd6784,17'd69361,17'd69549,17'd69817,17'd7425,17'd8222,17'd40269,17'd8849,17'd69903,17'd9442,17'd9441,17'd10116,17'd10116,17'd10116,17'd10116,17'd10116,17'd10114,17'd9303,17'd6304,17'd8692,17'd8070,17'd7097,17'd6638,17'd41780,17'd70397,17'd53817,17'd53817,17'd53612,17'd62226,17'd2650,17'd70398,17'd70399,17'd70400,17'd69906,17'd64000,17'd58522,17'd55584,17'd70401,17'd70402,17'd58659,17'd54990,17'd55779,17'd70403,17'd56457,17'd58152,17'd56351,17'd70404,17'd70405,17'd70406,17'd70407,17'd70408,17'd70409,17'd70410,17'd70411,17'd70412,17'd70413,17'd68672,17'd70414,17'd70201,17'd70415,17'd70011,17'd70416,17'd70417,17'd70418,17'd61989,17'd70419,17'd70420,17'd70421,17'd70422,17'd70423,17'd16298,17'd15277,17'd14786,17'd19025,17'd10704,17'd70424,17'd50401,17'd70425,17'd70426,17'd70427,17'd70428,17'd47882,17'd70429,17'd70430,17'd18451,17'd7790,17'd63446,17'd7788,17'd12120,17'd17482,17'd23688,17'd70431,17'd70432,17'd70433,17'd70434,17'd70435,17'd70436,17'd18696,17'd6368,17'd70437,17'd70438,17'd139,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd130,17'd130,17'd130,17'd130,17'd132,17'd11541,17'd11541,17'd52069,17'd52069,17'd69761,17'd52247,17'd69762,17'd70238,17'd70439,17'd52736,17'd70440,17'd67614,17'd70441,17'd51538,17'd70442,17'd52813,17'd52317,17'd70443,17'd70444,17'd70445,17'd70446,17'd70447,17'd51453,17'd70448,17'd70449,17'd21073,17'd69764,17'd67232,17'd51820,17'd51729,17'd65635,17'd23017,17'd20624,17'd11683,17'd131,17'd131,17'd131,17'd11541,17'd133,17'd131,17'd70349,17'd70450,17'd70451,17'd70452,17'd70453,17'd18467,17'd70454,17'd70455,17'd70456,17'd68915,17'd70457,17'd69869,17'd70458,17'd69591,17'd70360,17'd69403,17'd69871,17'd69783,17'd70051,17'd70459,17'd70460,17'd70362,17'd8622,17'd8771,17'd9515,17'd9515,17'd8623,17'd9231,17'd12283,17'd8762,17'd11161,17'd11161,17'd14715,17'd70461,17'd8292,17'd7175,17'd11850,17'd68823,17'd11573,17'd11708,17'd11315,17'd69787,17'd27932,17'd27933,17'd69692,17'd68928,17'd68825,17'd70364,17'd69879,17'd70252,17'd69880,17'd70154,17'd69971,17'd70154,17'd70462,17'd70463,17'd70464,17'd70257,17'd70159,17'd69235,17'd70465,17'd70466,17'd69794,17'd70467,17'd70468,17'd69338,17'd70469,17'd70469,17'd68518,17'd70259,17'd68517,17'd68517,17'd69144,17'd68059,17'd70264,17'd70262,17'd70470,17'd70471,17'd70472,17'd70473,17'd70473,17'd70474,17'd70264,17'd70264,17'd69524,17'd69523,17'd69706,17'd69706,17'd68944,17'd69338,17'd69340,17'd69340,17'd64650,17'd64526,17'd63962,17'd63962,17'd66197,17'd65950,17'd65950,17'd65950,17'd64387,17'd64387,17'd64387,17'd64387,17'd68520,17'd68520,17'd65054,17'd65054,17'd66072,17'd65054,17'd64387,17'd64387,17'd63963,17'd63963,17'd63963,17'd65308,17'd17179,17'd67427,17'd62576,17'd62576,17'd67557,17'd15618,17'd67426,17'd69342,17'd65705,17'd62701,17'd66322,17'd68741,17'd65040,17'd66063,17'd70374,17'd70475,17'd69887,17'd68949,17'd69241,17'd69241,17'd69241,17'd69241,17'd63511,17'd63511,17'd64653,17'd65055,17'd65831,17'd67439,17'd69424,17'd69889,17'd68947,17'd70476,17'd70477,17'd70477,17'd67296,17'd67439,17'd70478,17'd69711,17'd70479,17'd70480,17'd70481,17'd70378,17'd70060,17'd69523,17'd70482,17'd70483,17'd70483,17'd70484,17'd70485,17'd11336,17'd49008,17'd35907,17'd5371,17'd5050,17'd1823,17'd1243,17'd607,17'd271,17'd260,17'd206,17'd1829,17'd205,17'd14066,17'd1381
},
'{
17'd8509,17'd8509,17'd7046,17'd6422,17'd70486,17'd5376,17'd4735,17'd4427,17'd13943,17'd3751,17'd2783,17'd2593,17'd2784,17'd2781,17'd1689,17'd1689,17'd2781,17'd9968,17'd9968,17'd3750,17'd4247,17'd4247,17'd1127,17'd9968,17'd70487,17'd68751,17'd65957,17'd65959,17'd66327,17'd66205,17'd70280,17'd68962,17'd68423,17'd68308,17'd70488,17'd69055,17'd69435,17'd69620,17'd67446,17'd68304,17'd70285,17'd8512,17'd8191,17'd7218,17'd9270,17'd63259,17'd1415,17'd19,17'd11,17'd808,17'd19,17'd18,17'd0,17'd2,17'd2594,17'd4247,17'd1688,17'd1967,17'd2781,17'd3252,17'd10547,17'd3429,17'd2597,17'd2257,17'd17,17'd18,17'd19,17'd11,17'd11,17'd11,17'd27,17'd27,17'd652,17'd289,17'd3595,17'd3433,17'd5209,17'd5208,17'd6278,17'd11889,17'd11890,17'd6279,17'd10408,17'd69724,17'd8521,17'd70388,17'd6906,17'd6749,17'd8047,17'd68854,17'd70489,17'd70490,17'd70290,17'd70491,17'd70492,17'd70493,17'd70494,17'd69816,17'd25126,17'd36057,17'd37723,17'd37974,17'd69360,17'd38222,17'd70495,17'd70495,17'd38222,17'd69360,17'd69816,17'd7760,17'd8547,17'd8849,17'd67079,17'd65855,17'd28669,17'd9441,17'd9441,17'd9441,17'd9441,17'd9441,17'd10114,17'd10695,17'd6304,17'd6138,17'd6137,17'd8541,17'd68437,17'd7914,17'd42662,17'd6155,17'd70496,17'd53885,17'd53689,17'd60164,17'd70497,17'd70498,17'd70499,17'd70000,17'd70500,17'd55285,17'd70501,17'd70502,17'd62102,17'd58772,17'd63405,17'd63689,17'd61310,17'd66110,17'd70503,17'd60299,17'd54805,17'd70504,17'd70505,17'd70506,17'd70507,17'd70508,17'd70509,17'd70510,17'd70412,17'd70511,17'd70512,17'd70513,17'd70514,17'd70103,17'd70012,17'd70515,17'd70516,17'd70517,17'd69921,17'd70518,17'd70519,17'd70421,17'd70520,17'd70521,17'd17217,17'd70522,17'd19143,17'd70523,17'd9854,17'd70524,17'd28085,17'd70525,17'd70526,17'd70527,17'd70528,17'd70529,17'd7128,17'd38494,17'd67223,17'd53634,17'd9890,17'd15440,17'd11968,17'd10179,17'd22825,17'd70530,17'd70531,17'd70532,17'd70533,17'd70534,17'd70535,17'd70536,17'd6829,17'd70537,17'd70538,17'd127,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd130,17'd130,17'd130,17'd130,17'd132,17'd131,17'd131,17'd11541,17'd11541,17'd11541,17'd20623,17'd20465,17'd20625,17'd20625,17'd20629,17'd70539,17'd22148,17'd70540,17'd70541,17'd21222,17'd21070,17'd52071,17'd68893,17'd52418,17'd70542,17'd70542,17'd70542,17'd70543,17'd70544,17'd21223,17'd21682,17'd70545,17'd70546,17'd52053,17'd20626,17'd15823,17'd133,17'd131,17'd131,17'd134,17'd134,17'd132,17'd132,17'd133,17'd131,17'd70349,17'd70547,17'd70548,17'd70549,17'd70550,17'd70551,17'd70552,17'd70553,17'd70554,17'd70555,17'd70556,17'd70557,17'd70558,17'd68815,17'd69020,17'd69217,17'd69872,17'd70559,17'd70051,17'd70459,17'd70460,17'd10637,17'd8622,17'd8622,17'd9515,17'd9515,17'd8623,17'd9231,17'd69598,17'd11987,17'd11161,17'd8613,17'd70461,17'd70560,17'd7171,17'd6551,17'd10512,17'd68927,17'd11573,17'd70561,17'd69787,17'd69787,17'd28306,17'd28306,17'd27933,17'd33993,17'd68931,17'd70364,17'd69879,17'd70153,17'd70154,17'd70154,17'd69971,17'd70562,17'd70462,17'd70563,17'd70564,17'd70565,17'd70566,17'd69333,17'd67544,17'd70567,17'd70568,17'd70569,17'd70468,17'd69145,17'd70570,17'd70469,17'd66928,17'd66928,17'd67923,17'd68517,17'd69144,17'd68059,17'd70264,17'd70262,17'd70471,17'd70471,17'd70571,17'd70571,17'd70571,17'd70473,17'd70572,17'd70263,17'd69524,17'd69523,17'd69705,17'd69705,17'd68519,17'd69337,17'd68520,17'd68520,17'd64526,17'd64526,17'd63962,17'd63962,17'd66197,17'd66197,17'd66197,17'd66197,17'd64387,17'd64387,17'd64387,17'd64387,17'd68833,17'd68833,17'd65054,17'd65054,17'd65054,17'd65054,17'd64919,17'd66435,17'd66435,17'd63963,17'd63243,17'd62851,17'd67426,17'd62449,17'd62576,17'd62576,17'd67557,17'd15618,17'd67426,17'd67426,17'd62975,17'd70573,17'd70373,17'd65688,17'd66063,17'd67791,17'd70574,17'd70375,17'd70575,17'd68949,17'd69241,17'd69241,17'd68415,17'd68415,17'd63657,17'd64388,17'd64921,17'd66320,17'd67439,17'd67931,17'd69424,17'd69424,17'd69425,17'd70576,17'd70477,17'd70477,17'd67296,17'd67296,17'd70478,17'd70479,17'd70577,17'd70480,17'd70481,17'd70578,17'd70579,17'd70580,17'd70581,17'd70582,17'd70483,17'd70583,17'd36904,17'd11335,17'd70584,17'd35907,17'd5371,17'd5050,17'd1823,17'd1243,17'd607,17'd607,17'd260,17'd260,17'd606,17'd205,17'd2256,17'd1381
},
'{
17'd8509,17'd7046,17'd6262,17'd5643,17'd5376,17'd5645,17'd4735,17'd4087,17'd13943,17'd3901,17'd3901,17'd2593,17'd2784,17'd3250,17'd3750,17'd9815,17'd70277,17'd13186,17'd63257,17'd12503,17'd1689,17'd4247,17'd1127,17'd2781,17'd63518,17'd64665,17'd69249,17'd68849,17'd65959,17'd66086,17'd66205,17'd69436,17'd68193,17'd69055,17'd70585,17'd68310,17'd67814,17'd69620,17'd66941,17'd66327,17'd69809,17'd70586,17'd7886,17'd69161,17'd70587,17'd10543,17'd3249,17'd1,17'd19,17'd808,17'd979,17'd18,17'd0,17'd0,17'd1127,17'd2594,17'd1688,17'd1689,17'd1689,17'd1688,17'd2426,17'd2426,17'd2597,17'd1414,17'd1416,17'd18,17'd19,17'd979,17'd11,17'd11,17'd11,17'd10,17'd28,17'd29,17'd3595,17'd3433,17'd3254,17'd3255,17'd3756,17'd12655,17'd11890,17'd6279,17'd10408,17'd9276,17'd8521,17'd8198,17'd6906,17'd8199,17'd69724,17'd70588,17'd12037,17'd70589,17'd70590,17'd70591,17'd70080,17'd70592,17'd70593,17'd69817,17'd69628,17'd36922,17'd37322,17'd6943,17'd69264,17'd70594,17'd52206,17'd38093,17'd37838,17'd37320,17'd70595,17'd70596,17'd25260,17'd8383,17'd70087,17'd69167,17'd65727,17'd28669,17'd28669,17'd68095,17'd68095,17'd28669,17'd9842,17'd9842,17'd9303,17'd9303,17'd6138,17'd5088,17'd6627,17'd5085,17'd6639,17'd6313,17'd70397,17'd6012,17'd70597,17'd70598,17'd70599,17'd70600,17'd2993,17'd70601,17'd61056,17'd70602,17'd70603,17'd67084,17'd70604,17'd61189,17'd69632,17'd63405,17'd61440,17'd62876,17'd56581,17'd54704,17'd60421,17'd70605,17'd70606,17'd70607,17'd70608,17'd70609,17'd70610,17'd70510,17'd70611,17'd70612,17'd68873,17'd70200,17'd69917,17'd70613,17'd70104,17'd70614,17'd70615,17'd70616,17'd70014,17'd70617,17'd70519,17'd70421,17'd70520,17'd70521,17'd16183,17'd15407,17'd14644,17'd15153,17'd14232,17'd51028,17'd70618,17'd47978,17'd70619,17'd70620,17'd70621,17'd70622,17'd70623,17'd70624,17'd14006,17'd22135,17'd9890,17'd15440,17'd15693,17'd70625,17'd70626,17'd70627,17'd70628,17'd70629,17'd70630,17'd70631,17'd70632,17'd8276,17'd5465,17'd125,17'd355,17'd70217,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd5593,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd11541,17'd52069,17'd52664,17'd52492,17'd51715,17'd52498,17'd69200,17'd20767,17'd51624,17'd52736,17'd51624,17'd51624,17'd20766,17'd22148,17'd69935,17'd20627,17'd52069,17'd11541,17'd131,17'd132,17'd1481,17'd1480,17'd1481,17'd132,17'd130,17'd130,17'd132,17'd132,17'd133,17'd11541,17'd70349,17'd70633,17'd70634,17'd70635,17'd70636,17'd22370,17'd70637,17'd70638,17'd70639,17'd68809,17'd70640,17'd70641,17'd70642,17'd70643,17'd69020,17'd70644,17'd70645,17'd70559,17'd70051,17'd70646,17'd70647,17'd10374,17'd8771,17'd8622,17'd9515,17'd9515,17'd70648,17'd9380,17'd69598,17'd11987,17'd7833,17'd8613,17'd70461,17'd20993,17'd7171,17'd6551,17'd68823,17'd68927,17'd11180,17'd11315,17'd69787,17'd70649,17'd28305,17'd28183,17'd33993,17'd70650,17'd68933,17'd70651,17'd69879,17'd70153,17'd70154,17'd70154,17'd70652,17'd70653,17'd70462,17'd70654,17'd70655,17'd70656,17'd70657,17'd70658,17'd70659,17'd70660,17'd70661,17'd25367,17'd63110,17'd68833,17'd70469,17'd70662,17'd68519,17'd66928,17'd67923,17'd68517,17'd69144,17'd68059,17'd70264,17'd70262,17'd70472,17'd70571,17'd70663,17'd70664,17'd70663,17'd70571,17'd70665,17'd70470,17'd70666,17'd70667,17'd69524,17'd69523,17'd68519,17'd68944,17'd68833,17'd66317,17'd64387,17'd64387,17'd64387,17'd63807,17'd63807,17'd64387,17'd64387,17'd64387,17'd68833,17'd68833,17'd68833,17'd68833,17'd66319,17'd66319,17'd66319,17'd66319,17'd65181,17'd65054,17'd66435,17'd67049,17'd66435,17'd63375,17'd62851,17'd62850,17'd69342,17'd62449,17'd67557,17'd67557,17'd15999,17'd15483,17'd67426,17'd17179,17'd62701,17'd70373,17'd65040,17'd66063,17'd67791,17'd70668,17'd70669,17'd70670,17'd68290,17'd68290,17'd68415,17'd68415,17'd67932,17'd67800,17'd64921,17'd64921,17'd65055,17'd67296,17'd67931,17'd70167,17'd69424,17'd67673,17'd69039,17'd68633,17'd67437,17'd70477,17'd69711,17'd69711,17'd70671,17'd70671,17'd70577,17'd70480,17'd70481,17'd70672,17'd70673,17'd70674,17'd70675,17'd70582,17'd70676,17'd70677,17'd11061,17'd5776,17'd70584,17'd35907,17'd5372,17'd4084,17'd410,17'd1243,17'd260,17'd260,17'd260,17'd259,17'd425,17'd972,17'd1244,17'd1381
},
'{
17'd8509,17'd7046,17'd7368,17'd5375,17'd5792,17'd5645,17'd4735,17'd5201,17'd4893,17'd5204,17'd4086,17'd2783,17'd2782,17'd2592,17'd9968,17'd70678,17'd70679,17'd70680,17'd11608,17'd63386,17'd9815,17'd1688,17'd1688,17'd3250,17'd11887,17'd70681,17'd67816,17'd68755,17'd69809,17'd66206,17'd70682,17'd68964,17'd67941,17'd70683,17'd69806,17'd70684,17'd70685,17'd66813,17'd66814,17'd68964,17'd67179,17'd9130,17'd8515,17'd12033,17'd6591,17'd11607,17'd9684,17'd1967,17'd18,17'd10,17'd979,17'd19,17'd0,17'd0,17'd1127,17'd4247,17'd1688,17'd1688,17'd1689,17'd1689,17'd2258,17'd2426,17'd2258,17'd2596,17'd1414,17'd16,17'd979,17'd979,17'd11,17'd11,17'd11,17'd10,17'd287,17'd288,17'd3755,17'd3595,17'd3254,17'd3254,17'd3756,17'd11210,17'd11737,17'd6279,17'd10408,17'd9685,17'd70686,17'd8198,17'd6907,17'd6907,17'd70687,17'd70688,17'd7562,17'd70689,17'd70690,17'd70691,17'd70692,17'd70693,17'd67461,17'd70694,17'd63421,17'd70695,17'd37322,17'd69359,17'd69733,17'd70696,17'd70495,17'd38221,17'd70697,17'd70698,17'd70699,17'd37975,17'd70700,17'd68540,17'd70701,17'd70702,17'd70703,17'd70703,17'd8380,17'd8380,17'd8847,17'd9985,17'd9985,17'd9985,17'd6304,17'd9303,17'd9303,17'd5089,17'd4925,17'd5250,17'd7089,17'd6475,17'd6319,17'd53690,17'd70704,17'd70705,17'd70706,17'd70707,17'd70708,17'd70709,17'd70710,17'd62097,17'd54891,17'd70502,17'd67199,17'd57133,17'd61188,17'd61188,17'd61310,17'd56911,17'd54802,17'd70711,17'd60536,17'd70712,17'd70606,17'd70713,17'd70714,17'd70715,17'd69640,17'd70716,17'd70717,17'd70718,17'd70719,17'd70720,17'd70103,17'd70314,17'd70721,17'd70316,17'd70722,17'd70723,17'd70205,17'd70420,17'd70724,17'd70519,17'd70520,17'd70521,17'd15659,17'd14644,17'd70725,17'd70726,17'd11923,17'd27723,17'd70727,17'd47678,17'd47494,17'd70728,17'd70729,17'd70730,17'd70731,17'd70624,17'd7456,17'd22135,17'd9890,17'd15692,17'd10995,17'd70732,17'd70733,17'd70734,17'd70735,17'd70736,17'd70737,17'd70738,17'd70739,17'd70740,17'd70741,17'd70742,17'd70743,17'd70744,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd5593,17'd131,17'd131,17'd132,17'd132,17'd132,17'd134,17'd131,17'd131,17'd131,17'd131,17'd11541,17'd11541,17'd131,17'd131,17'd131,17'd131,17'd20623,17'd20623,17'd11541,17'd131,17'd132,17'd130,17'd136,17'd136,17'd129,17'd129,17'd70438,17'd70438,17'd130,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd11541,17'd70349,17'd70745,17'd70746,17'd70747,17'd70748,17'd70749,17'd70750,17'd70751,17'd67398,17'd69116,17'd70752,17'd70753,17'd70643,17'd70643,17'd70754,17'd70755,17'd70756,17'd70757,17'd70758,17'd70759,17'd70760,17'd70761,17'd8771,17'd8622,17'd9515,17'd9515,17'd9381,17'd15458,17'd14841,17'd11987,17'd7832,17'd7833,17'd11423,17'd10883,17'd7171,17'd6385,17'd68823,17'd11573,17'd11430,17'd11315,17'd69787,17'd70649,17'd28305,17'd28183,17'd33993,17'd33993,17'd70762,17'd69131,17'd69602,17'd70153,17'd70154,17'd70763,17'd70562,17'd70653,17'd70764,17'd70654,17'd70655,17'd70765,17'd70766,17'd70767,17'd70768,17'd70660,17'd64901,17'd25232,17'd68840,17'd63243,17'd70165,17'd70570,17'd68519,17'd66928,17'd67923,17'd68517,17'd69144,17'd69144,17'd70263,17'd70262,17'd70472,17'd70571,17'd70663,17'd70664,17'd70664,17'd70664,17'd70663,17'd70571,17'd70769,17'd70770,17'd69524,17'd69524,17'd68519,17'd66318,17'd66317,17'd66436,17'd66317,17'd64919,17'd64919,17'd64387,17'd64387,17'd64919,17'd64919,17'd68833,17'd68833,17'd68833,17'd68833,17'd66319,17'd66319,17'd66318,17'd66318,17'd66319,17'd65054,17'd66072,17'd66073,17'd64530,17'd69712,17'd63375,17'd62850,17'd62700,17'd14734,17'd62449,17'd15618,17'd15618,17'd15999,17'd15999,17'd67426,17'd68836,17'd70373,17'd65040,17'd66063,17'd67791,17'd70668,17'd70668,17'd70668,17'd70668,17'd70771,17'd68290,17'd68415,17'd68415,17'd67932,17'd66198,17'd64921,17'd67295,17'd66320,17'd67439,17'd70167,17'd70772,17'd68632,17'd68633,17'd69426,17'd69039,17'd67437,17'd70477,17'd70773,17'd69711,17'd70479,17'd70671,17'd70577,17'd70774,17'd70481,17'd70672,17'd70775,17'd70572,17'd70675,17'd70582,17'd70776,17'd60625,17'd11335,17'd5630,17'd35907,17'd5372,17'd6407,17'd4084,17'd1243,17'd970,17'd260,17'd260,17'd259,17'd1666,17'd605,17'd971,17'd1244,17'd1381
},
'{
17'd7046,17'd7046,17'd7368,17'd5198,17'd5645,17'd5645,17'd4735,17'd5201,17'd6730,17'd5204,17'd4086,17'd2783,17'd6424,17'd7371,17'd9968,17'd63257,17'd13302,17'd70777,17'd70777,17'd70778,17'd63257,17'd7371,17'd2422,17'd3250,17'd6265,17'd63518,17'd66693,17'd69249,17'd65844,17'd68752,17'd65843,17'd70779,17'd70780,17'd68962,17'd67304,17'd70684,17'd67690,17'd66812,17'd70781,17'd66208,17'd65957,17'd9126,17'd7220,17'd7547,17'd13064,17'd10799,17'd69723,17'd9815,17'd17,17'd11,17'd3748,17'd19,17'd2,17'd2,17'd2,17'd466,17'd2594,17'd2594,17'd1689,17'd1967,17'd2597,17'd12194,17'd2426,17'd2597,17'd1414,17'd17,17'd19,17'd979,17'd10,17'd11,17'd10,17'd10,17'd287,17'd28,17'd29,17'd30,17'd3254,17'd3254,17'd3255,17'd6278,17'd11211,17'd6439,17'd9555,17'd9555,17'd9685,17'd69724,17'd7390,17'd69810,17'd7390,17'd7227,17'd9970,17'd70782,17'd70783,17'd70784,17'd70785,17'd70786,17'd70787,17'd70788,17'd70789,17'd69733,17'd6943,17'd6943,17'd70790,17'd70696,17'd69168,17'd70791,17'd38606,17'd70697,17'd37837,17'd70792,17'd70793,17'd68860,17'd69996,17'd69995,17'd70794,17'd70794,17'd8071,17'd8379,17'd8220,17'd8847,17'd8847,17'd64275,17'd64275,17'd64275,17'd64275,17'd6136,17'd5088,17'd5688,17'd70795,17'd7089,17'd63137,17'd70796,17'd70797,17'd70798,17'd63157,17'd70598,17'd70799,17'd5093,17'd2996,17'd70800,17'd65987,17'd62727,17'd66110,17'd56242,17'd56242,17'd56352,17'd56352,17'd64145,17'd60422,17'd60537,17'd70801,17'd70802,17'd70803,17'd70804,17'd70805,17'd70806,17'd69640,17'd70807,17'd70807,17'd69828,17'd70808,17'd70809,17'd70613,17'd70810,17'd70811,17'd70812,17'd70813,17'd70814,17'd70815,17'd70519,17'd70816,17'd70520,17'd70817,17'd16892,17'd15659,17'd14785,17'd14643,17'd26024,17'd26988,17'd27965,17'd48567,17'd47493,17'd30362,17'd70818,17'd70729,17'd7281,17'd70731,17'd70819,17'd70820,17'd24714,17'd7619,17'd15193,17'd15060,17'd70821,17'd70822,17'd70823,17'd70824,17'd70825,17'd70826,17'd70827,17'd70828,17'd70829,17'd70830,17'd70831,17'd70832,17'd70833,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd131,17'd131,17'd131,17'd131,17'd132,17'd130,17'd130,17'd132,17'd131,17'd131,17'd132,17'd132,17'd134,17'd134,17'd134,17'd134,17'd134,17'd20466,17'd131,17'd131,17'd131,17'd132,17'd132,17'd128,17'd138,17'd128,17'd132,17'd131,17'd133,17'd542,17'd133,17'd132,17'd130,17'd130,17'd130,17'd130,17'd1481,17'd11541,17'd70349,17'd70834,17'd70835,17'd70836,17'd70837,17'd70838,17'd70839,17'd70840,17'd70841,17'd70842,17'd70843,17'd70844,17'd16591,17'd69020,17'd69403,17'd69871,17'd70845,17'd70846,17'd70847,17'd70848,17'd70849,17'd10772,17'd8771,17'd8622,17'd70850,17'd70850,17'd9381,17'd14411,17'd14841,17'd9506,17'd7832,17'd7498,17'd10883,17'd10499,17'd70851,17'd6551,17'd68823,17'd11573,17'd11430,17'd11315,17'd11181,17'd11181,17'd28183,17'd28183,17'd68929,17'd70650,17'd69031,17'd70651,17'd69412,17'd70153,17'd70154,17'd70763,17'd70653,17'd70653,17'd70764,17'd70654,17'd70852,17'd70853,17'd70766,17'd70767,17'd70768,17'd67030,17'd70854,17'd70855,17'd70856,17'd62971,17'd70857,17'd70570,17'd68519,17'd68519,17'd68060,17'd68517,17'd68517,17'd69144,17'd70263,17'd70572,17'd70665,17'd70571,17'd70663,17'd70664,17'd70858,17'd70859,17'd70860,17'd70663,17'd70769,17'd70861,17'd70770,17'd69524,17'd68519,17'd66318,17'd66072,17'd66676,17'd67049,17'd66435,17'd64919,17'd64919,17'd66319,17'd66319,17'd66319,17'd66319,17'd68833,17'd68833,17'd68944,17'd68944,17'd66318,17'd70862,17'd68060,17'd68060,17'd66677,17'd66437,17'd67671,17'd64530,17'd63656,17'd62852,17'd62700,17'd67425,17'd69342,17'd67426,17'd15483,17'd15483,17'd15483,17'd15999,17'd67425,17'd68836,17'd70166,17'd65553,17'd64506,17'd67918,17'd70863,17'd70863,17'd70864,17'd70865,17'd68290,17'd68290,17'd68949,17'd69887,17'd69243,17'd66198,17'd67295,17'd70477,17'd67437,17'd68187,17'd70065,17'd70065,17'd67672,17'd69426,17'd66199,17'd67674,17'd67296,17'd66320,17'd70773,17'd70773,17'd70866,17'd70866,17'd70867,17'd70868,17'd70869,17'd70775,17'd70470,17'd70572,17'd70870,17'd70871,17'd27822,17'd27949,17'd9123,17'd4423,17'd5372,17'd5372,17'd2740,17'd191,17'd803,17'd643,17'd206,17'd643,17'd606,17'd425,17'd971,17'd1272,17'd1244,17'd1381
},
'{
17'd6423,17'd6423,17'd6262,17'd10397,17'd5645,17'd5376,17'd4735,17'd4735,17'd4893,17'd4737,17'd64251,17'd63384,17'd63255,17'd68191,17'd68075,17'd11887,17'd70872,17'd70872,17'd70873,17'd70872,17'd70874,17'd63256,17'd2592,17'd2781,17'd2781,17'd63257,17'd64122,17'd69050,17'd66808,17'd69051,17'd68313,17'd70875,17'd70876,17'd70877,17'd66813,17'd68530,17'd70073,17'd70878,17'd67182,17'd67692,17'd9417,17'd69056,17'd8515,17'd7886,17'd67574,17'd6894,17'd67306,17'd70777,17'd0,17'd1128,17'd979,17'd979,17'd0,17'd2,17'd2,17'd2,17'd2594,17'd2594,17'd1688,17'd1689,17'd2597,17'd2426,17'd2426,17'd2258,17'd2257,17'd1415,17'd16,17'd979,17'd10,17'd10,17'd10,17'd10,17'd287,17'd70879,17'd2118,17'd809,17'd3254,17'd3254,17'd3255,17'd3755,17'd6598,17'd5972,17'd9555,17'd9555,17'd9685,17'd9685,17'd70687,17'd69810,17'd7390,17'd7063,17'd7557,17'd70880,17'd70881,17'd70882,17'd70883,17'd70884,17'd69900,17'd70885,17'd70886,17'd70887,17'd37974,17'd37056,17'd70084,17'd70295,17'd70888,17'd37972,17'd6947,17'd38606,17'd37838,17'd38351,17'd70889,17'd70890,17'd70793,17'd70891,17'd70085,17'd7424,17'd70892,17'd8377,17'd8377,17'd8072,17'd8072,17'd65462,17'd65462,17'd65462,17'd69999,17'd69999,17'd5998,17'd5998,17'd5250,17'd4923,17'd3947,17'd3138,17'd70893,17'd70894,17'd53816,17'd60788,17'd64014,17'd70895,17'd70896,17'd70897,17'd70898,17'd70899,17'd70900,17'd70901,17'd64145,17'd56456,17'd70501,17'd60299,17'd60170,17'd63542,17'd64551,17'd70902,17'd70903,17'd70904,17'd70905,17'd70906,17'd70907,17'd70807,17'd70908,17'd68875,17'd70909,17'd70910,17'd70314,17'd70810,17'd70105,17'd70911,17'd70912,17'd60943,17'd70815,17'd70519,17'd70816,17'd70520,17'd70913,17'd16532,17'd16183,17'd70914,17'd20039,17'd11097,17'd70915,17'd70916,17'd70917,17'd47284,17'd70918,17'd70919,17'd70920,17'd70921,17'd70922,17'd70923,17'd70924,17'd24714,17'd15439,17'd70925,17'd59840,17'd70926,17'd70927,17'd70928,17'd70929,17'd70930,17'd70931,17'd70932,17'd70933,17'd70934,17'd70935,17'd70936,17'd70937,17'd355,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd131,17'd132,17'd130,17'd130,17'd128,17'd128,17'd11541,17'd11541,17'd131,17'd131,17'd130,17'd130,17'd130,17'd132,17'd131,17'd131,17'd132,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd131,17'd11541,17'd11541,17'd11541,17'd134,17'd134,17'd130,17'd130,17'd130,17'd131,17'd131,17'd133,17'd133,17'd131,17'd131,17'd135,17'd129,17'd130,17'd130,17'd130,17'd131,17'd53482,17'd70938,17'd70939,17'd70940,17'd70941,17'd70942,17'd70943,17'd70944,17'd70945,17'd70946,17'd70641,17'd68716,17'd69019,17'd69020,17'd69403,17'd69592,17'd70845,17'd70846,17'd70847,17'd70848,17'd70947,17'd10772,17'd8771,17'd9080,17'd70850,17'd70648,17'd70948,17'd14411,17'd70949,17'd9506,17'd7833,17'd70950,17'd70461,17'd10883,17'd69690,17'd70951,17'd68823,17'd11573,17'd11430,17'd11315,17'd27932,17'd11181,17'd28183,17'd28183,17'd68929,17'd33993,17'd70762,17'd69226,17'd69602,17'd70153,17'd70154,17'd70763,17'd70653,17'd70952,17'd70764,17'd70953,17'd70954,17'd70955,17'd70956,17'd70957,17'd70958,17'd67030,17'd70959,17'd70960,17'd70961,17'd66678,17'd70857,17'd70570,17'd68519,17'd68519,17'd68060,17'd68517,17'd68517,17'd68517,17'd70163,17'd70262,17'd70473,17'd70571,17'd70663,17'd70664,17'd70858,17'd70858,17'd70860,17'd70860,17'd70962,17'd70769,17'd70666,17'd69524,17'd68519,17'd65054,17'd64651,17'd66073,17'd66435,17'd66435,17'd64919,17'd64919,17'd66319,17'd66319,17'd69337,17'd69337,17'd66318,17'd68945,17'd68519,17'd68519,17'd68060,17'd67923,17'd67923,17'd67923,17'd67423,17'd67423,17'd67671,17'd63808,17'd66078,17'd62853,17'd67425,17'd70963,17'd67426,17'd67426,17'd16959,17'd15483,17'd15483,17'd67425,17'd68836,17'd70373,17'd70166,17'd65289,17'd68058,17'd67918,17'd70863,17'd70863,17'd70964,17'd70668,17'd70771,17'd68740,17'd69887,17'd69710,17'd66198,17'd69242,17'd70965,17'd70477,17'd68187,17'd68298,17'd70065,17'd70167,17'd67673,17'd69426,17'd66199,17'd67674,17'd67296,17'd66320,17'd69711,17'd69711,17'd70866,17'd70866,17'd70867,17'd70966,17'd70868,17'd70967,17'd70371,17'd70770,17'd70582,17'd70776,17'd29170,17'd58863,17'd5940,17'd4423,17'd5372,17'd6407,17'd26595,17'd411,17'd803,17'd643,17'd206,17'd643,17'd425,17'd605,17'd1272,17'd1272,17'd1381,17'd1244
},
'{
17'd6423,17'd6423,17'd6262,17'd10397,17'd5645,17'd5376,17'd4735,17'd4735,17'd64116,17'd70968,17'd70969,17'd70970,17'd11344,17'd11887,17'd12652,17'd12652,17'd70873,17'd70971,17'd67693,17'd70278,17'd70972,17'd63518,17'd6265,17'd2781,17'd2594,17'd3249,17'd63667,17'd64796,17'd67062,17'd66552,17'd68965,17'd65956,17'd70973,17'd70974,17'd67181,17'd69433,17'd68643,17'd67571,17'd66811,17'd66331,17'd70975,17'd70976,17'd70977,17'd10660,17'd8043,17'd7547,17'd6894,17'd63668,17'd67308,17'd18,17'd19,17'd3748,17'd3,17'd12,17'd2,17'd2,17'd4247,17'd4247,17'd4247,17'd1127,17'd2596,17'd2597,17'd2258,17'd2426,17'd2257,17'd1414,17'd17,17'd19,17'd808,17'd808,17'd10,17'd11,17'd979,17'd979,17'd288,17'd981,17'd3255,17'd3254,17'd3255,17'd3755,17'd6438,17'd6745,17'd6439,17'd10408,17'd10408,17'd10409,17'd70686,17'd8198,17'd70978,17'd6749,17'd7063,17'd7731,17'd70979,17'd70980,17'd70981,17'd70982,17'd70983,17'd65971,17'd70984,17'd70985,17'd37058,17'd37595,17'd37322,17'd70986,17'd70295,17'd70696,17'd37972,17'd37839,17'd38093,17'd39058,17'd70987,17'd70988,17'd52113,17'd38888,17'd70891,17'd70891,17'd70989,17'd70990,17'd7916,17'd64273,17'd64813,17'd64813,17'd70991,17'd69999,17'd69999,17'd64680,17'd69904,17'd5084,17'd4125,17'd52625,17'd4128,17'd3948,17'd70992,17'd6935,17'd6310,17'd53689,17'd70993,17'd70994,17'd70995,17'd70996,17'd4933,17'd70997,17'd70998,17'd70300,17'd56455,17'd57387,17'd58032,17'd70000,17'd59930,17'd66701,17'd70999,17'd71000,17'd71001,17'd71002,17'd71003,17'd69556,17'd71004,17'd71005,17'd71006,17'd71007,17'd71008,17'd71009,17'd71010,17'd71011,17'd71012,17'd71013,17'd71014,17'd62245,17'd70518,17'd70724,17'd70816,17'd70520,17'd70913,17'd16532,17'd16183,17'd71015,17'd14906,17'd26858,17'd28929,17'd71016,17'd71017,17'd71018,17'd71019,17'd71020,17'd71021,17'd71022,17'd43080,17'd70923,17'd70924,17'd18567,17'd53634,17'd25153,17'd52875,17'd71023,17'd71024,17'd71025,17'd71026,17'd71027,17'd71028,17'd71029,17'd71030,17'd71031,17'd71032,17'd71033,17'd71034,17'd71035,17'd136,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd131,17'd132,17'd130,17'd136,17'd136,17'd136,17'd132,17'd132,17'd134,17'd134,17'd128,17'd136,17'd130,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd135,17'd135,17'd1197,17'd719,17'd133,17'd131,17'd132,17'd135,17'd132,17'd132,17'd1197,17'd131,17'd71036,17'd71037,17'd71038,17'd71039,17'd71040,17'd71041,17'd71042,17'd71043,17'd71044,17'd70946,17'd71045,17'd68716,17'd68921,17'd70246,17'd71046,17'd71047,17'd71048,17'd71049,17'd71050,17'd71051,17'd70947,17'd10772,17'd8622,17'd9080,17'd70850,17'd70648,17'd70948,17'd14717,17'd15087,17'd15463,17'd7833,17'd7835,17'd70560,17'd10499,17'd71052,17'd70951,17'd68823,17'd11180,17'd11430,17'd11315,17'd27932,17'd11181,17'd28183,17'd28183,17'd68929,17'd68724,17'd69031,17'd68932,17'd69412,17'd70153,17'd70154,17'd71053,17'd70653,17'd70952,17'd71054,17'd71055,17'd71056,17'd71057,17'd71058,17'd71059,17'd71060,17'd70161,17'd71061,17'd64087,17'd63790,17'd66536,17'd71062,17'd70662,17'd68518,17'd68519,17'd67923,17'd68517,17'd71063,17'd71063,17'd70163,17'd70262,17'd70473,17'd70571,17'd71064,17'd70860,17'd71065,17'd71066,17'd71066,17'd70858,17'd71067,17'd71068,17'd71069,17'd69796,17'd68182,17'd71070,17'd63654,17'd63655,17'd63244,17'd64651,17'd66072,17'd66437,17'd66928,17'd68519,17'd69797,17'd69706,17'd68518,17'd68518,17'd68518,17'd71071,17'd69144,17'd69144,17'd68517,17'd67923,17'd68292,17'd67423,17'd66676,17'd63375,17'd65441,17'd62700,17'd65705,17'd67426,17'd67426,17'd15483,17'd65949,17'd65949,17'd67435,17'd62850,17'd65441,17'd68741,17'd65553,17'd71072,17'd68058,17'd71073,17'd70863,17'd71074,17'd70964,17'd70376,17'd68740,17'd68181,17'd69710,17'd71075,17'd66075,17'd66199,17'd69039,17'd69425,17'd71076,17'd71076,17'd71076,17'd67438,17'd68633,17'd66076,17'd71077,17'd71077,17'd65831,17'd65831,17'd69800,17'd69800,17'd71078,17'd70066,17'd70168,17'd70162,17'd70261,17'd70371,17'd71069,17'd70581,17'd71079,17'd35770,17'd28544,17'd58244,17'd5372,17'd1810,17'd6407,17'd192,17'd1098,17'd1685,17'd972,17'd1966,17'd1966,17'd1966,17'd205,17'd971,17'd1244,17'd1381,17'd1381,17'd1244
},
'{
17'd6423,17'd5375,17'd10397,17'd10397,17'd5645,17'd5376,17'd4735,17'd4735,17'd14744,17'd14443,17'd71080,17'd71081,17'd71082,17'd63517,17'd71083,17'd69617,17'd69617,17'd71084,17'd63820,17'd65188,17'd65068,17'd71085,17'd63256,17'd3250,17'd2594,17'd1967,17'd12652,17'd71086,17'd68751,17'd67683,17'd68965,17'd67683,17'd65956,17'd71087,17'd68644,17'd71088,17'd68643,17'd70073,17'd71089,17'd66445,17'd71090,17'd65957,17'd70976,17'd8974,17'd8975,17'd8043,17'd7547,17'd6740,17'd63258,17'd1277,17'd16,17'd3748,17'd650,17'd3,17'd0,17'd466,17'd4247,17'd1127,17'd1127,17'd1127,17'd1414,17'd1414,17'd2597,17'd2426,17'd2257,17'd2257,17'd1415,17'd1277,17'd3748,17'd808,17'd10,17'd11,17'd11,17'd979,17'd288,17'd981,17'd3255,17'd3254,17'd3255,17'd3255,17'd5207,17'd6437,17'd6903,17'd10408,17'd10408,17'd10409,17'd71091,17'd70687,17'd70978,17'd6906,17'd7559,17'd71092,17'd71093,17'd71094,17'd71095,17'd71096,17'd71097,17'd71098,17'd71099,17'd71100,17'd39201,17'd71101,17'd37056,17'd71102,17'd70891,17'd70891,17'd71103,17'd38094,17'd38093,17'd39058,17'd71104,17'd71105,17'd6642,17'd52205,17'd6783,17'd6783,17'd71106,17'd68656,17'd71107,17'd70990,17'd71108,17'd71108,17'd65325,17'd65325,17'd65325,17'd42795,17'd42795,17'd67466,17'd4122,17'd52029,17'd4922,17'd4290,17'd71109,17'd71110,17'd2986,17'd60532,17'd60163,17'd5415,17'd2658,17'd71111,17'd71112,17'd71113,17'd71114,17'd56809,17'd61056,17'd70711,17'd71115,17'd71116,17'd59930,17'd66701,17'd71117,17'd71118,17'd71001,17'd71002,17'd71119,17'd71120,17'd71121,17'd71122,17'd71123,17'd71124,17'd70200,17'd71125,17'd70810,17'd71126,17'd71127,17'd71128,17'd71129,17'd61080,17'd70419,17'd71130,17'd71131,17'd70520,17'd70816,17'd16892,17'd15659,17'd19633,17'd22466,17'd71132,17'd28210,17'd71133,17'd71134,17'd71135,17'd71136,17'd71137,17'd71138,17'd71139,17'd71140,17'd71141,17'd42227,17'd7293,17'd53634,17'd25414,17'd71142,17'd71143,17'd71144,17'd71145,17'd71146,17'd71147,17'd71148,17'd71149,17'd71150,17'd71151,17'd71152,17'd71153,17'd70937,17'd71154,17'd70438,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd131,17'd132,17'd130,17'd136,17'd136,17'd136,17'd130,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd132,17'd131,17'd11541,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd11541,17'd131,17'd131,17'd131,17'd131,17'd131,17'd134,17'd134,17'd132,17'd132,17'd1481,17'd133,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd1197,17'd5593,17'd71155,17'd71156,17'd71157,17'd71158,17'd71159,17'd71160,17'd28033,17'd71161,17'd71044,17'd71162,17'd71163,17'd68815,17'd68921,17'd71164,17'd71046,17'd69502,17'd71165,17'd71049,17'd71050,17'd71166,17'd71167,17'd10772,17'd8622,17'd9080,17'd70850,17'd70648,17'd71168,17'd14717,17'd14707,17'd9506,17'd13672,17'd8613,17'd70461,17'd10883,17'd7495,17'd6385,17'd68823,17'd11180,17'd11430,17'd11315,17'd27932,17'd11181,17'd28183,17'd28183,17'd68824,17'd68929,17'd70762,17'd68932,17'd69969,17'd70153,17'd71169,17'd71170,17'd71171,17'd70952,17'd71172,17'd71173,17'd71174,17'd71175,17'd71176,17'd71177,17'd71178,17'd70161,17'd71179,17'd70568,17'd25367,17'd66306,17'd64791,17'd70061,17'd68518,17'd66928,17'd67923,17'd68517,17'd71063,17'd71063,17'd70163,17'd70262,17'd70472,17'd70571,17'd71064,17'd70860,17'd71180,17'd71066,17'd71181,17'd71181,17'd70858,17'd71182,17'd71183,17'd69796,17'd68182,17'd71184,17'd71185,17'd71186,17'd65305,17'd65305,17'd67423,17'd68517,17'd69703,17'd69796,17'd69796,17'd69796,17'd69703,17'd69703,17'd69703,17'd69703,17'd69703,17'd69703,17'd68517,17'd68517,17'd67423,17'd67671,17'd63808,17'd62972,17'd62853,17'd67425,17'd67426,17'd67426,17'd15483,17'd15483,17'd65949,17'd15483,17'd67435,17'd62974,17'd66790,17'd65688,17'd69334,17'd69142,17'd71073,17'd71187,17'd70863,17'd71188,17'd70864,17'd70575,17'd67919,17'd68181,17'd71075,17'd68739,17'd66199,17'd66076,17'd67673,17'd68947,17'd71189,17'd71189,17'd71190,17'd69039,17'd66199,17'd67674,17'd71077,17'd66077,17'd65055,17'd69800,17'd71191,17'd71191,17'd70866,17'd70066,17'd70168,17'd70162,17'd70261,17'd70371,17'd70666,17'd71192,17'd65564,17'd31251,17'd31899,17'd16382,17'd5371,17'd5957,17'd5957,17'd604,17'd411,17'd971,17'd972,17'd205,17'd1966,17'd1966,17'd972,17'd424,17'd1381,17'd1381,17'd1381,17'd1244
},
'{
17'd5510,17'd6422,17'd10397,17'd10397,17'd5645,17'd5377,17'd5201,17'd4734,17'd5646,17'd4426,17'd71193,17'd65711,17'd65187,17'd67061,17'd71194,17'd63816,17'd65065,17'd64122,17'd71195,17'd71195,17'd71195,17'd63978,17'd71196,17'd6260,17'd4576,17'd5196,17'd70277,17'd71197,17'd64397,17'd71198,17'd69051,17'd66552,17'd71199,17'd69809,17'd66208,17'd71200,17'd66939,17'd68310,17'd69433,17'd71201,17'd70877,17'd71202,17'd71203,17'd9126,17'd10085,17'd71204,17'd8344,17'd7547,17'd64667,17'd10668,17'd1127,17'd3,17'd979,17'd19,17'd1277,17'd17,17'd1414,17'd2257,17'd27442,17'd22965,17'd466,17'd466,17'd4247,17'd10535,17'd10535,17'd4247,17'd14,17'd2,17'd16,17'd979,17'd10,17'd10,17'd1128,17'd11,17'd287,17'd70879,17'd3907,17'd3254,17'd2940,17'd3255,17'd4091,17'd6438,17'd6903,17'd10408,17'd10408,17'd10408,17'd9685,17'd70688,17'd8198,17'd70388,17'd7559,17'd9817,17'd70782,17'd71205,17'd71206,17'd71207,17'd71208,17'd69992,17'd71209,17'd71210,17'd71211,17'd37057,17'd71212,17'd37323,17'd69359,17'd69733,17'd69549,17'd71103,17'd38351,17'd38482,17'd6646,17'd39058,17'd6645,17'd71213,17'd6642,17'd52286,17'd52552,17'd71214,17'd64015,17'd64015,17'd64413,17'd6778,17'd7098,17'd7421,17'd7421,17'd7097,17'd41019,17'd7097,17'd67466,17'd60783,17'd6772,17'd71215,17'd3627,17'd3946,17'd59642,17'd2987,17'd3134,17'd2649,17'd4299,17'd3486,17'd54896,17'd1873,17'd71216,17'd71217,17'd61056,17'd71218,17'd54704,17'd70088,17'd55901,17'd71219,17'd71220,17'd71221,17'd71222,17'd71223,17'd71224,17'd71225,17'd71226,17'd71227,17'd71228,17'd71229,17'd71230,17'd71231,17'd71232,17'd71127,17'd70616,17'd62245,17'd61080,17'd71233,17'd71234,17'd71235,17'd71130,17'd71236,17'd17106,17'd16533,17'd16048,17'd71237,17'd71238,17'd29908,17'd71239,17'd30962,17'd31934,17'd71240,17'd71241,17'd71242,17'd71243,17'd71244,17'd42807,17'd71245,17'd71246,17'd71247,17'd18451,17'd71248,17'd71249,17'd70734,17'd71250,17'd71251,17'd71252,17'd71253,17'd71254,17'd71255,17'd71256,17'd71257,17'd71258,17'd71259,17'd71260,17'd127,17'd1480,17'd541,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd1481,17'd1481,17'd132,17'd132,17'd131,17'd131,17'd131,17'd132,17'd130,17'd1481,17'd356,17'd5593,17'd71261,17'd71262,17'd71263,17'd71264,17'd71265,17'd29272,17'd71266,17'd71267,17'd71268,17'd71269,17'd70458,17'd71270,17'd70246,17'd69122,17'd71271,17'd71272,17'd71273,17'd71049,17'd70847,17'd71274,17'd10215,17'd8772,17'd8771,17'd71275,17'd71276,17'd9079,17'd12147,17'd8153,17'd8149,17'd13672,17'd11296,17'd9371,17'd71277,17'd27929,17'd7826,17'd6217,17'd11036,17'd9932,17'd11430,17'd11315,17'd27932,17'd28305,17'd28183,17'd28183,17'd68510,17'd69692,17'd68724,17'd70651,17'd69969,17'd70153,17'd71169,17'd71169,17'd71278,17'd70764,17'd71055,17'd71279,17'd71280,17'd71281,17'd71282,17'd70956,17'd71283,17'd71284,17'd66177,17'd70568,17'd67665,17'd65688,17'd69712,17'd71062,17'd66072,17'd66318,17'd66928,17'd71285,17'd69144,17'd69144,17'd69524,17'd71286,17'd70470,17'd70769,17'd70571,17'd70663,17'd70860,17'd71180,17'd71287,17'd71066,17'd71288,17'd71182,17'd71068,17'd70471,17'd70264,17'd71289,17'd71290,17'd71185,17'd67423,17'd68517,17'd71291,17'd70260,17'd70371,17'd70572,17'd70572,17'd70262,17'd70163,17'd70162,17'd70261,17'd71292,17'd71292,17'd69703,17'd71285,17'd70259,17'd66437,17'd66317,17'd63963,17'd62850,17'd71293,17'd15999,17'd15483,17'd16959,17'd15348,17'd15348,17'd15483,17'd15483,17'd62853,17'd66790,17'd64507,17'd64903,17'd69142,17'd71294,17'd71295,17'd71294,17'd71296,17'd70668,17'd70575,17'd70376,17'd71297,17'd71298,17'd68739,17'd66199,17'd66320,17'd67296,17'd68187,17'd70167,17'd69889,17'd68632,17'd69039,17'd66076,17'd67674,17'd67674,17'd67296,17'd69711,17'd69711,17'd71299,17'd70479,17'd70671,17'd71299,17'd71300,17'd70269,17'd71301,17'd70371,17'd70666,17'd71302,17'd71303,17'd36904,17'd11061,17'd11335,17'd9123,17'd4880,17'd5957,17'd1667,17'd1111,17'd803,17'd803,17'd1687,17'd1829,17'd936,17'd205,17'd1244,17'd1381,17'd1381,17'd1382,17'd1381,17'd1244
},
'{
17'd5510,17'd6422,17'd5198,17'd5198,17'd5645,17'd5377,17'd5201,17'd4734,17'd5646,17'd5646,17'd71304,17'd71305,17'd71306,17'd71307,17'd71308,17'd71309,17'd64795,17'd64121,17'd64120,17'd65449,17'd71195,17'd71310,17'd67693,17'd71311,17'd6583,17'd5196,17'd6583,17'd71312,17'd63978,17'd67816,17'd66552,17'd69250,17'd65717,17'd68082,17'd65960,17'd66330,17'd66689,17'd68197,17'd67571,17'd71088,17'd67688,17'd71313,17'd71314,17'd71315,17'd9127,17'd9127,17'd65718,17'd8043,17'd71316,17'd9967,17'd3249,17'd2,17'd979,17'd808,17'd18,17'd16,17'd1415,17'd2257,17'd27442,17'd22965,17'd466,17'd466,17'd4247,17'd1831,17'd10535,17'd1688,17'd1127,17'd14,17'd17,17'd1277,17'd979,17'd10,17'd20,17'd11,17'd28,17'd288,17'd3907,17'd3254,17'd2940,17'd2941,17'd3255,17'd4431,17'd10093,17'd6903,17'd10408,17'd10408,17'd71317,17'd70688,17'd71318,17'd71319,17'd7559,17'd7064,17'd71320,17'd71321,17'd69623,17'd71322,17'd69543,17'd71323,17'd71324,17'd71325,17'd71326,17'd37460,17'd37723,17'd37594,17'd69549,17'd70295,17'd69549,17'd69360,17'd38094,17'd38093,17'd40275,17'd38482,17'd38482,17'd38891,17'd38891,17'd39504,17'd51419,17'd52285,17'd52552,17'd71327,17'd71328,17'd71328,17'd6778,17'd6778,17'd7420,17'd7420,17'd6780,17'd7097,17'd67587,17'd60783,17'd6772,17'd71329,17'd71215,17'd59643,17'd3623,17'd3624,17'd3295,17'd2989,17'd4130,17'd54174,17'd71330,17'd70601,17'd71331,17'd71217,17'd71332,17'd61836,17'd70187,17'd54892,17'd64000,17'd71219,17'd71333,17'd71334,17'd71335,17'd71336,17'd71337,17'd71338,17'd71339,17'd71340,17'd71341,17'd71342,17'd70910,17'd71343,17'd71344,17'd71345,17'd59418,17'd71346,17'd71233,17'd62125,17'd71347,17'd71348,17'd71130,17'd17106,17'd71349,17'd16533,17'd71350,17'd25663,17'd71351,17'd54639,17'd71352,17'd71017,17'd71353,17'd71354,17'd71355,17'd71356,17'd42805,17'd71357,17'd71358,17'd71359,17'd71246,17'd38903,17'd18451,17'd70116,17'd71360,17'd71361,17'd71362,17'd71363,17'd71364,17'd71365,17'd71366,17'd71367,17'd71368,17'd71369,17'd71370,17'd71371,17'd71372,17'd720,17'd1480,17'd541,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd1481,17'd1481,17'd132,17'd132,17'd131,17'd131,17'd131,17'd132,17'd1481,17'd20762,17'd541,17'd5593,17'd71373,17'd71374,17'd71375,17'd71376,17'd71377,17'd71378,17'd71379,17'd71380,17'd71268,17'd71162,17'd71163,17'd71381,17'd69120,17'd69121,17'd71272,17'd71382,17'd71383,17'd71384,17'd71385,17'd71274,17'd71386,17'd8773,17'd8622,17'd71275,17'd71276,17'd9079,17'd8464,17'd7996,17'd7995,17'd7832,17'd11296,17'd9640,17'd71387,17'd71388,17'd7175,17'd11849,17'd68823,17'd9932,17'd11430,17'd69787,17'd28306,17'd28305,17'd28183,17'd28183,17'd68510,17'd69692,17'd68724,17'd69129,17'd69969,17'd71389,17'd71169,17'd71390,17'd71391,17'd71392,17'd71393,17'd71394,17'd71395,17'd71396,17'd71397,17'd70656,17'd70767,17'd71398,17'd66423,17'd71399,17'd71400,17'd65421,17'd63510,17'd64530,17'd66072,17'd66437,17'd70259,17'd71285,17'd69703,17'd69144,17'd69796,17'd71286,17'd70470,17'd70471,17'd70571,17'd71401,17'd71402,17'd70860,17'd71403,17'd71065,17'd70858,17'd71404,17'd71405,17'd71068,17'd70264,17'd71406,17'd71407,17'd67794,17'd70059,17'd70261,17'd70260,17'd70371,17'd70473,17'd70473,17'd70473,17'd70775,17'd70869,17'd70868,17'd70261,17'd70261,17'd69703,17'd68517,17'd71285,17'd66804,17'd66317,17'd66435,17'd65308,17'd67435,17'd15483,17'd15999,17'd15483,17'd15483,17'd15348,17'd15483,17'd16959,17'd62700,17'd63110,17'd64904,17'd68736,17'd71408,17'd71409,17'd67550,17'd71410,17'd71411,17'd71187,17'd70668,17'd70575,17'd71412,17'd71413,17'd71414,17'd68948,17'd66076,17'd67296,17'd67439,17'd68298,17'd70065,17'd69424,17'd67672,17'd71415,17'd71416,17'd67674,17'd67674,17'd66320,17'd69711,17'd71299,17'd70479,17'd70479,17'd70479,17'd71417,17'd71418,17'd70378,17'd70260,17'd70371,17'd70770,17'd71419,17'd71420,17'd36903,17'd5183,17'd5776,17'd5630,17'd4880,17'd5957,17'd1667,17'd1396,17'd644,17'd644,17'd1687,17'd1124,17'd1966,17'd204,17'd1244,17'd1381,17'd1382,17'd1382,17'd1381,17'd1244
},
'{
17'd5790,17'd5790,17'd5643,17'd5198,17'd5645,17'd5377,17'd5202,17'd4735,17'd5646,17'd5646,17'd5202,17'd71421,17'd71422,17'd71307,17'd71308,17'd71423,17'd63976,17'd63977,17'd64929,17'd66693,17'd64397,17'd63979,17'd12928,17'd70278,17'd71424,17'd6583,17'd4886,17'd71425,17'd65188,17'd70070,17'd67183,17'd71426,17'd69056,17'd71427,17'd66206,17'd66208,17'd67688,17'd67063,17'd67572,17'd69435,17'd67181,17'd71428,17'd69808,17'd68082,17'd8664,17'd9129,17'd68755,17'd67815,17'd6894,17'd67306,17'd9684,17'd4247,17'd979,17'd16389,17'd1128,17'd19,17'd17,17'd1414,17'd2257,17'd2425,17'd4247,17'd1127,17'd1127,17'd4247,17'd1831,17'd1688,17'd1127,17'd1127,17'd17,17'd18,17'd10,17'd10,17'd21,17'd20,17'd27,17'd288,17'd3907,17'd3255,17'd2941,17'd2940,17'd1129,17'd3754,17'd6598,17'd10093,17'd10408,17'd10408,17'd10409,17'd10409,17'd69724,17'd8198,17'd7559,17'd7064,17'd6282,17'd71429,17'd71430,17'd71431,17'd69353,17'd71432,17'd71433,17'd67582,17'd71434,17'd6784,17'd71435,17'd69448,17'd69448,17'd69448,17'd69361,17'd69361,17'd6784,17'd38094,17'd6643,17'd38890,17'd38482,17'd38482,17'd71436,17'd38891,17'd39504,17'd51419,17'd49203,17'd51256,17'd68655,17'd71437,17'd66954,17'd66954,17'd7421,17'd42795,17'd42795,17'd43069,17'd5084,17'd5084,17'd6933,17'd4463,17'd4463,17'd4290,17'd71215,17'd59643,17'd63138,17'd3467,17'd2980,17'd2299,17'd54174,17'd2994,17'd71438,17'd71438,17'd71439,17'd71438,17'd54703,17'd56905,17'd59930,17'd66348,17'd71440,17'd68328,17'd71441,17'd71442,17'd71443,17'd71444,17'd71445,17'd71446,17'd71447,17'd71448,17'd71449,17'd71450,17'd70812,17'd71345,17'd60943,17'd71451,17'd71452,17'd71453,17'd71454,17'd9168,17'd9709,17'd17331,17'd16668,17'd23329,17'd19767,17'd71455,17'd71456,17'd52938,17'd47876,17'd71134,17'd71457,17'd71458,17'd71459,17'd71460,17'd71461,17'd71462,17'd71463,17'd71464,17'd7131,17'd7292,17'd15059,17'd71465,17'd71466,17'd71467,17'd71468,17'd71469,17'd71470,17'd71471,17'd71472,17'd71473,17'd71474,17'd71475,17'd71370,17'd71476,17'd71477,17'd128,17'd1481,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd1481,17'd1481,17'd132,17'd132,17'd131,17'd131,17'd131,17'd132,17'd356,17'd20762,17'd356,17'd5593,17'd71478,17'd71479,17'd71480,17'd71481,17'd71482,17'd71483,17'd71484,17'd71485,17'd71486,17'd71487,17'd71488,17'd71489,17'd71490,17'd69322,17'd69405,17'd69405,17'd71273,17'd71491,17'd71492,17'd71274,17'd71493,17'd71494,17'd9080,17'd9080,17'd71276,17'd9380,17'd8464,17'd7996,17'd7995,17'd13672,17'd9506,17'd8611,17'd71495,17'd71496,17'd6847,17'd6850,17'd11036,17'd9932,17'd11430,17'd11315,17'd27932,17'd28305,17'd28183,17'd28183,17'd68622,17'd69692,17'd68724,17'd71497,17'd71498,17'd71389,17'd71499,17'd71500,17'd71501,17'd70764,17'd71502,17'd71503,17'd71504,17'd71505,17'd71506,17'd70656,17'd71507,17'd69139,17'd66423,17'd65036,17'd66533,17'd65421,17'd71508,17'd69712,17'd66073,17'd66072,17'd70259,17'd71285,17'd71071,17'd71071,17'd69524,17'd69796,17'd70470,17'd70470,17'd70571,17'd71401,17'd71064,17'd70860,17'd71065,17'd71065,17'd71509,17'd70859,17'd70663,17'd70571,17'd70572,17'd70264,17'd70263,17'd70371,17'd71510,17'd71510,17'd71510,17'd70472,17'd70472,17'd70571,17'd71511,17'd71512,17'd71510,17'd70967,17'd70261,17'd70163,17'd68517,17'd68517,17'd70259,17'd66804,17'd64387,17'd63107,17'd62850,17'd71293,17'd15483,17'd15483,17'd15483,17'd15483,17'd15483,17'd16959,17'd65571,17'd62853,17'd68741,17'd65688,17'd65815,17'd70863,17'd71294,17'd71513,17'd71411,17'd71411,17'd71187,17'd70669,17'd70376,17'd69710,17'd71514,17'd68948,17'd66076,17'd67674,17'd67438,17'd68187,17'd70167,17'd70065,17'd67672,17'd67673,17'd67674,17'd66076,17'd67674,17'd67296,17'd69711,17'd70773,17'd65056,17'd69800,17'd71515,17'd70268,17'd70269,17'd70269,17'd70162,17'd70261,17'd71286,17'd71302,17'd71303,17'd36904,17'd11882,17'd4714,17'd8185,17'd4880,17'd5050,17'd5050,17'd1111,17'd425,17'd643,17'd644,17'd1124,17'd1124,17'd205,17'd204,17'd1244,17'd202,17'd1382,17'd1382,17'd1381,17'd1244
},
'{
17'd5644,17'd5790,17'd5643,17'd5643,17'd5645,17'd5377,17'd5202,17'd5201,17'd4426,17'd4426,17'd5201,17'd71304,17'd71516,17'd71307,17'd71517,17'd71518,17'd64120,17'd64121,17'd64929,17'd71195,17'd64397,17'd64254,17'd63979,17'd63820,17'd71311,17'd6583,17'd5196,17'd6096,17'd71519,17'd71195,17'd65582,17'd68853,17'd9265,17'd71520,17'd70875,17'd66088,17'd69436,17'd69720,17'd67304,17'd68426,17'd69620,17'd70877,17'd71090,17'd9675,17'd69056,17'd9130,17'd8513,17'd67815,17'd8043,17'd6737,17'd63668,17'd9815,17'd0,17'd10,17'd11,17'd19,17'd16,17'd1415,17'd2597,17'd2597,17'd1688,17'd1127,17'd1127,17'd1127,17'd1831,17'd1688,17'd4247,17'd4247,17'd1416,17'd16,17'd19,17'd10,17'd10,17'd11,17'd27,17'd28,17'd4431,17'd3755,17'd3254,17'd2940,17'd469,17'd1693,17'd3907,17'd10093,17'd10408,17'd10408,17'd10408,17'd6904,17'd8048,17'd71521,17'd69986,17'd6906,17'd8049,17'd71522,17'd5061,17'd71523,17'd71524,17'd71525,17'd71526,17'd71527,17'd71528,17'd71529,17'd71530,17'd71531,17'd69448,17'd71103,17'd6784,17'd6784,17'd69360,17'd71103,17'd70792,17'd6643,17'd38093,17'd38482,17'd71436,17'd38891,17'd71532,17'd49015,17'd49203,17'd46999,17'd53086,17'd71437,17'd71437,17'd66954,17'd7421,17'd42795,17'd42795,17'd43069,17'd8541,17'd5250,17'd44521,17'd4126,17'd44521,17'd60290,17'd4922,17'd62873,17'd63137,17'd3137,17'd3134,17'd60291,17'd71533,17'd71534,17'd71535,17'd71536,17'd71537,17'd71538,17'd71539,17'd56905,17'd54618,17'd65468,17'd71440,17'd4459,17'd71540,17'd71541,17'd71542,17'd71543,17'd71544,17'd71447,17'd71545,17'd71546,17'd71547,17'd71548,17'd71549,17'd71550,17'd61080,17'd71551,17'd71552,17'd71553,17'd71348,17'd9169,17'd9588,17'd16532,17'd16893,17'd16048,17'd20039,17'd10131,17'd71554,17'd71555,17'd71556,17'd71353,17'd71557,17'd71558,17'd71559,17'd71560,17'd6963,17'd71561,17'd71562,17'd71563,17'd71564,17'd71565,17'd25292,17'd71566,17'd71567,17'd71568,17'd71569,17'd71570,17'd71571,17'd71572,17'd71573,17'd71574,17'd71575,17'd71576,17'd71577,17'd71578,17'd139,17'd130,17'd130,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd1481,17'd130,17'd132,17'd132,17'd131,17'd131,17'd131,17'd132,17'd356,17'd1481,17'd133,17'd11683,17'd71579,17'd71580,17'd71581,17'd71582,17'd71583,17'd71584,17'd71585,17'd71586,17'd71587,17'd71487,17'd71488,17'd71588,17'd69322,17'd69871,17'd69502,17'd69684,17'd71383,17'd71384,17'd71385,17'd71274,17'd71589,17'd71386,17'd8773,17'd9080,17'd71276,17'd9380,17'd8464,17'd7996,17'd7995,17'd7832,17'd11296,17'd8611,17'd71590,17'd71388,17'd6848,17'd11849,17'd68823,17'd9932,17'd11430,17'd69787,17'd28306,17'd28305,17'd28183,17'd28183,17'd68622,17'd69692,17'd68724,17'd69129,17'd69969,17'd71389,17'd71499,17'd71500,17'd71501,17'd71591,17'd71592,17'd71593,17'd71594,17'd71595,17'd71506,17'd70656,17'd71507,17'd68941,17'd66423,17'd65036,17'd66662,17'd65687,17'd71596,17'd63510,17'd64651,17'd66072,17'd66928,17'd70259,17'd68518,17'd68518,17'd69523,17'd69524,17'd70572,17'd70470,17'd70472,17'd70571,17'd71401,17'd71402,17'd70860,17'd71065,17'd71509,17'd70858,17'd70664,17'd70663,17'd71068,17'd70471,17'd71597,17'd71598,17'd71599,17'd71600,17'd71600,17'd71401,17'd70571,17'd70571,17'd71601,17'd71512,17'd71510,17'd71602,17'd70260,17'd70163,17'd68517,17'd67923,17'd66437,17'd66073,17'd63243,17'd71603,17'd67435,17'd71293,17'd15483,17'd15483,17'd15483,17'd15999,17'd15483,17'd62700,17'd62853,17'd66678,17'd65688,17'd68736,17'd71604,17'd71605,17'd71606,17'd71411,17'd71411,17'd71607,17'd70863,17'd70669,17'd70670,17'd71608,17'd71609,17'd71416,17'd67674,17'd67558,17'd68187,17'd68298,17'd70167,17'd70167,17'd67673,17'd69039,17'd66076,17'd66076,17'd67674,17'd66320,17'd66320,17'd70773,17'd65056,17'd71191,17'd71515,17'd71610,17'd71611,17'd70868,17'd70260,17'd71286,17'd71612,17'd71613,17'd63652,17'd35487,17'd5183,17'd5940,17'd5371,17'd4881,17'd5050,17'd5050,17'd605,17'd425,17'd643,17'd643,17'd1124,17'd1966,17'd204,17'd424,17'd202,17'd1382,17'd1382,17'd1382,17'd1381,17'd2256
},
'{
17'd5199,17'd5199,17'd6421,17'd5053,17'd5645,17'd5376,17'd5202,17'd5202,17'd5646,17'd4087,17'd5201,17'd5202,17'd71614,17'd71306,17'd71517,17'd71309,17'd65579,17'd64120,17'd64929,17'd64929,17'd64397,17'd66693,17'd71195,17'd71615,17'd70278,17'd71424,17'd6583,17'd6583,17'd71311,17'd65067,17'd70070,17'd69249,17'd8513,17'd65844,17'd71616,17'd67179,17'd66332,17'd68531,17'd69620,17'd69435,17'd69435,17'd67688,17'd67692,17'd71617,17'd71618,17'd69056,17'd8662,17'd9265,17'd69249,17'd7052,17'd67306,17'd65314,17'd14,17'd12,17'd10,17'd10,17'd18,17'd1415,17'd10268,17'd3752,17'd3752,17'd2597,17'd1414,17'd1414,17'd2597,17'd2597,17'd2597,17'd2257,17'd1416,17'd17,17'd19,17'd10,17'd10,17'd10,17'd27,17'd28,17'd29,17'd981,17'd3255,17'd2940,17'd292,17'd12036,17'd11210,17'd10269,17'd11211,17'd10672,17'd6441,17'd6441,17'd6747,17'd6905,17'd69986,17'd7559,17'd6907,17'd71619,17'd71320,17'd71620,17'd69542,17'd71621,17'd71622,17'd71623,17'd71624,17'd68539,17'd71625,17'd71626,17'd70594,17'd70594,17'd70495,17'd6784,17'd69549,17'd69448,17'd71103,17'd38222,17'd38351,17'd38093,17'd38890,17'd71213,17'd39504,17'd49015,17'd49203,17'd46895,17'd51256,17'd53086,17'd71437,17'd66954,17'd6937,17'd71627,17'd67587,17'd43069,17'd8541,17'd8541,17'd70795,17'd70795,17'd5250,17'd44521,17'd5084,17'd67466,17'd63681,17'd61301,17'd3137,17'd3134,17'd60162,17'd4931,17'd2468,17'd4301,17'd2996,17'd71628,17'd56695,17'd57387,17'd59646,17'd53880,17'd59511,17'd71629,17'd71630,17'd71631,17'd71632,17'd71633,17'd71634,17'd71635,17'd71636,17'd71637,17'd71638,17'd71639,17'd71640,17'd70723,17'd71641,17'd61459,17'd71642,17'd71643,17'd10295,17'd9851,17'd16667,17'd16182,17'd22983,17'd27465,17'd70726,17'd11633,17'd71644,17'd71645,17'd71646,17'd71647,17'd71648,17'd45085,17'd71649,17'd71650,17'd71651,17'd71652,17'd71653,17'd71654,17'd71564,17'd71655,17'd71656,17'd71657,17'd71658,17'd71659,17'd71660,17'd71661,17'd71662,17'd71663,17'd71664,17'd71665,17'd71666,17'd71667,17'd71668,17'd71669,17'd138,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd1481,17'd20762,17'd130,17'd5593,17'd71670,17'd71671,17'd71672,17'd71673,17'd71674,17'd71675,17'd71676,17'd71677,17'd71678,17'd68504,17'd71679,17'd71680,17'd69322,17'd69872,17'd70050,17'd69404,17'd71681,17'd71049,17'd71682,17'd71051,17'd71683,17'd71684,17'd71685,17'd71686,17'd16116,17'd71687,17'd8464,17'd8464,17'd8153,17'd13672,17'd9373,17'd8611,17'd71590,17'd71496,17'd6847,17'd10512,17'd11036,17'd9932,17'd11430,17'd69787,17'd28305,17'd28305,17'd28183,17'd28183,17'd68622,17'd69692,17'd68724,17'd68930,17'd71498,17'd71389,17'd71499,17'd71500,17'd71688,17'd71689,17'd71690,17'd71691,17'd71692,17'd71693,17'd71175,17'd70765,17'd71694,17'd71695,17'd66177,17'd70661,17'd67036,17'd63639,17'd66538,17'd66078,17'd64651,17'd66072,17'd66928,17'd66928,17'd68519,17'd68518,17'd69523,17'd69523,17'd69796,17'd70666,17'd70572,17'd70769,17'd71068,17'd70663,17'd70663,17'd70859,17'd70859,17'd70858,17'd71696,17'd70664,17'd71401,17'd71697,17'd71698,17'd71698,17'd71401,17'd71401,17'd71401,17'd70663,17'd71064,17'd71064,17'd71511,17'd71699,17'd70775,17'd70371,17'd70260,17'd70261,17'd68517,17'd66928,17'd64919,17'd63963,17'd65950,17'd62850,17'd15483,17'd67426,17'd67426,17'd67426,17'd15483,17'd15483,17'd62700,17'd62700,17'd69240,17'd70166,17'd66063,17'd69334,17'd71073,17'd71187,17'd71607,17'd71607,17'd71607,17'd71700,17'd71700,17'd71701,17'd71702,17'd71514,17'd71703,17'd71704,17'd69039,17'd67672,17'd68298,17'd68298,17'd68298,17'd68298,17'd69039,17'd68633,17'd68633,17'd68633,17'd66320,17'd66320,17'd66320,17'd67295,17'd65055,17'd71191,17'd71515,17'd71300,17'd67921,17'd70162,17'd71292,17'd69796,17'd71613,17'd71705,17'd36903,17'd11061,17'd6889,17'd6415,17'd3391,17'd1261,17'd1667,17'd1823,17'd644,17'd643,17'd206,17'd643,17'd1966,17'd205,17'd424,17'd1272,17'd202,17'd1382,17'd1382,17'd1382,17'd1244,17'd13940
},
'{
17'd5199,17'd33216,17'd5199,17'd6421,17'd5645,17'd5376,17'd5202,17'd9959,17'd4578,17'd4426,17'd5201,17'd5201,17'd71706,17'd71305,17'd71707,17'd71308,17'd64119,17'd65581,17'd64396,17'd64121,17'd71195,17'd71195,17'd71708,17'd64397,17'd63980,17'd71311,17'd6583,17'd7711,17'd71424,17'd71709,17'd64397,17'd67816,17'd65845,17'd70176,17'd71710,17'd65842,17'd9807,17'd69350,17'd68644,17'd69620,17'd69435,17'd71711,17'd66209,17'd71712,17'd66210,17'd68082,17'd69809,17'd9674,17'd65718,17'd71713,17'd69161,17'd71714,17'd12929,17'd2,17'd10,17'd10,17'd19,17'd16,17'd2936,17'd10268,17'd3752,17'd2597,17'd1414,17'd1415,17'd2596,17'd2597,17'd2597,17'd2597,17'd1414,17'd1416,17'd18,17'd979,17'd10,17'd10,17'd27,17'd27,17'd28,17'd29,17'd3755,17'd2941,17'd292,17'd470,17'd11208,17'd10269,17'd11211,17'd10672,17'd6441,17'd6441,17'd6747,17'd6905,17'd7559,17'd7559,17'd7559,17'd7228,17'd6282,17'd71321,17'd71715,17'd71716,17'd71717,17'd71718,17'd71719,17'd71720,17'd71721,17'd71722,17'd71531,17'd70594,17'd38094,17'd38222,17'd69448,17'd70086,17'd69448,17'd69549,17'd38222,17'd52206,17'd51773,17'd51773,17'd52286,17'd52285,17'd49203,17'd46895,17'd51256,17'd51256,17'd53086,17'd71437,17'd71437,17'd6937,17'd6937,17'd67587,17'd7421,17'd42795,17'd43069,17'd5084,17'd70795,17'd70795,17'd5084,17'd5084,17'd67466,17'd64140,17'd63683,17'd63402,17'd3294,17'd2982,17'd2826,17'd4773,17'd71535,17'd70709,17'd71723,17'd71724,17'd71725,17'd64818,17'd53018,17'd71726,17'd71727,17'd71728,17'd71729,17'd71730,17'd71635,17'd71731,17'd71732,17'd71733,17'd71638,17'd71734,17'd71735,17'd71736,17'd71552,17'd71737,17'd71738,17'd71739,17'd9315,17'd9589,17'd16782,17'd16182,17'd71740,17'd71741,17'd10437,17'd12073,17'd32115,17'd71742,17'd71743,17'd71744,17'd71745,17'd71746,17'd71747,17'd71748,17'd71749,17'd71750,17'd71751,17'd71752,17'd71653,17'd71753,17'd63584,17'd71754,17'd71755,17'd71756,17'd71757,17'd71758,17'd71759,17'd71760,17'd71761,17'd71762,17'd71763,17'd71764,17'd71668,17'd71765,17'd138,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd1481,17'd1481,17'd132,17'd70349,17'd71766,17'd71767,17'd71768,17'd71769,17'd71770,17'd71771,17'd71772,17'd71773,17'd71774,17'd68504,17'd71679,17'd69681,17'd69682,17'd71775,17'd71776,17'd71273,17'd71777,17'd71384,17'd71778,17'd71779,17'd71780,17'd71781,17'd71782,17'd71686,17'd16116,17'd71783,17'd8464,17'd8464,17'd8153,17'd7832,17'd10362,17'd8611,17'd71590,17'd28649,17'd6847,17'd11851,17'd68823,17'd11430,17'd71784,17'd69787,17'd28305,17'd28305,17'd28183,17'd28183,17'd68510,17'd69692,17'd70650,17'd69029,17'd69969,17'd71389,17'd71499,17'd71785,17'd71786,17'd71787,17'd71788,17'd71789,17'd71790,17'd71791,17'd71792,17'd71793,17'd71694,17'd71695,17'd71794,17'd71795,17'd67036,17'd65555,17'd71796,17'd66789,17'd63244,17'd66072,17'd66437,17'd66928,17'd68518,17'd68518,17'd69523,17'd69523,17'd69524,17'd69524,17'd70674,17'd70674,17'd70572,17'd70769,17'd70769,17'd70962,17'd70962,17'd71797,17'd70664,17'd70664,17'd71401,17'd71697,17'd71697,17'd71401,17'd70663,17'd70663,17'd70663,17'd70663,17'd71064,17'd71064,17'd71511,17'd70473,17'd70572,17'd70262,17'd70262,17'd69703,17'd70259,17'd66072,17'd63243,17'd62971,17'd62850,17'd67435,17'd67426,17'd67426,17'd67426,17'd67426,17'd15483,17'd67426,17'd62853,17'd63110,17'd71798,17'd65421,17'd69334,17'd71073,17'd71294,17'd71294,17'd71607,17'd71607,17'd71700,17'd71701,17'd71701,17'd71702,17'd71799,17'd71800,17'd71801,17'd68738,17'd67673,17'd67672,17'd68298,17'd68298,17'd68187,17'd67438,17'd68633,17'd68633,17'd69039,17'd69039,17'd66320,17'd66320,17'd66320,17'd66320,17'd65831,17'd66077,17'd65056,17'd70269,17'd68293,17'd70261,17'd71286,17'd70482,17'd71802,17'd71803,17'd11882,17'd4714,17'd1946,17'd5372,17'd445,17'd1261,17'd1823,17'd1396,17'd643,17'd643,17'd643,17'd643,17'd205,17'd972,17'd1272,17'd952,17'd1382,17'd1382,17'd1382,17'd1382,17'd2256,17'd71804
},
'{
17'd29756,17'd30047,17'd5202,17'd4735,17'd4734,17'd5201,17'd5202,17'd9959,17'd4426,17'd5646,17'd5201,17'd5202,17'd7212,17'd71805,17'd71806,17'd71307,17'd71807,17'd65579,17'd64396,17'd64121,17'd70487,17'd71708,17'd64537,17'd65449,17'd13433,17'd70278,17'd71808,17'd7711,17'd2781,17'd11887,17'd67576,17'd64123,17'd67815,17'd8513,17'd69249,17'd71809,17'd68082,17'd9674,17'd70071,17'd66559,17'd71810,17'd71810,17'd66331,17'd71090,17'd9809,17'd9265,17'd68082,17'd8662,17'd68853,17'd67815,17'd7547,17'd13815,17'd11736,17'd3749,17'd1275,17'd8814,17'd11,17'd19,17'd17187,17'd10268,17'd3752,17'd2597,17'd1414,17'd1414,17'd2596,17'd2597,17'd2597,17'd2596,17'd1414,17'd1416,17'd3905,17'd19,17'd11,17'd10,17'd286,17'd27,17'd28,17'd288,17'd3907,17'd3754,17'd292,17'd2942,17'd3435,17'd6278,17'd11211,17'd10408,17'd6441,17'd6441,17'd6747,17'd6748,17'd71521,17'd7559,17'd7559,17'd7063,17'd7228,17'd71522,17'd71811,17'd71812,17'd71813,17'd70080,17'd71814,17'd71815,17'd71816,17'd71817,17'd71626,17'd71818,17'd38095,17'd38096,17'd69448,17'd69448,17'd70086,17'd70295,17'd68860,17'd70793,17'd71106,17'd39055,17'd52785,17'd52474,17'd52552,17'd47094,17'd52552,17'd52552,17'd52552,17'd71327,17'd53086,17'd71437,17'd6636,17'd6636,17'd53168,17'd53169,17'd6937,17'd71627,17'd42795,17'd69904,17'd8541,17'd8541,17'd7089,17'd7421,17'd71819,17'd65201,17'd6477,17'd63137,17'd71820,17'd2982,17'd71821,17'd2013,17'd71822,17'd54433,17'd64818,17'd59012,17'd58641,17'd71823,17'd71824,17'd71825,17'd71826,17'd71730,17'd71827,17'd71828,17'd71829,17'd71830,17'd71639,17'd71831,17'd71832,17'd61080,17'd71833,17'd62892,17'd63021,17'd71834,17'd10129,17'd17582,17'd24844,17'd71740,17'd16047,17'd15405,17'd9995,17'd29625,17'd71835,17'd33232,17'd35223,17'd71836,17'd71837,17'd71838,17'd71839,17'd71840,17'd6806,17'd71841,17'd71842,17'd71843,17'd71653,17'd71844,17'd71845,17'd71846,17'd71847,17'd71848,17'd71849,17'd71850,17'd71851,17'd71852,17'd71853,17'd71854,17'd71855,17'd71856,17'd71668,17'd71857,17'd136,17'd132,17'd2698,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd133,17'd133,17'd1481,17'd1481,17'd134,17'd71858,17'd71859,17'd71860,17'd71861,17'd71862,17'd71863,17'd71864,17'd71865,17'd71866,17'd71867,17'd68812,17'd71489,17'd71588,17'd69592,17'd71868,17'd71869,17'd71681,17'd71870,17'd71871,17'd71872,17'd71873,17'd71874,17'd71875,17'd71876,17'd71686,17'd9381,17'd71783,17'd13794,17'd13794,17'd8153,17'd11296,17'd14716,17'd8611,17'd71495,17'd28649,17'd6386,17'd11035,17'd11179,17'd11180,17'd11315,17'd69787,17'd28305,17'd28305,17'd28305,17'd28183,17'd68510,17'd69692,17'd70650,17'd69029,17'd69969,17'd71389,17'd71499,17'd71877,17'd71878,17'd71879,17'd71880,17'd71881,17'd71882,17'd71883,17'd71884,17'd71885,17'd71886,17'd71887,17'd71888,17'd71889,17'd26956,17'd64769,17'd65042,17'd65556,17'd63656,17'd66072,17'd66437,17'd66928,17'd68519,17'd68518,17'd68518,17'd68519,17'd69523,17'd69523,17'd69523,17'd69523,17'd69524,17'd70667,17'd70770,17'd71890,17'd71891,17'd71891,17'd71892,17'd71405,17'd71405,17'd71405,17'd71405,17'd71182,17'd71404,17'd71893,17'd71893,17'd71893,17'd70663,17'd70962,17'd70571,17'd70473,17'd70572,17'd70572,17'd69796,17'd69144,17'd66928,17'd64387,17'd65950,17'd62850,17'd16959,17'd17179,17'd67426,17'd69342,17'd69342,17'd69342,17'd17179,17'd65571,17'd67163,17'd68741,17'd63789,17'd71072,17'd71894,17'd71895,17'd71896,17'd71411,17'd71897,17'd71700,17'd71898,17'd71413,17'd71414,17'd71609,17'd71899,17'd71900,17'd68838,17'd71901,17'd67672,17'd68632,17'd69424,17'd68632,17'd67438,17'd67437,17'd68633,17'd69039,17'd67437,17'd67437,17'd66320,17'd66320,17'd66320,17'd67296,17'd66077,17'd69800,17'd71610,17'd70269,17'd70059,17'd71292,17'd71902,17'd71613,17'd63652,17'd36903,17'd2906,17'd3073,17'd5372,17'd5050,17'd1823,17'd1823,17'd1243,17'd970,17'd643,17'd643,17'd1124,17'd1124,17'd205,17'd971,17'd1244,17'd1381,17'd1382,17'd1382,17'd603,17'd952,17'd204,17'd71903
},
'{
17'd29756,17'd10533,17'd5202,17'd4735,17'd4734,17'd4735,17'd5202,17'd69718,17'd4427,17'd4578,17'd5201,17'd69718,17'd5377,17'd5377,17'd71904,17'd71306,17'd71905,17'd63975,17'd64396,17'd64121,17'd63977,17'd64120,17'd65713,17'd65581,17'd66693,17'd63820,17'd71311,17'd6096,17'd3750,17'd6265,17'd70874,17'd71086,17'd68751,17'd68853,17'd7378,17'd68848,17'd71906,17'd12189,17'd66088,17'd66331,17'd67182,17'd67573,17'd71907,17'd66089,17'd9547,17'd8978,17'd65958,17'd71618,17'd7718,17'd67815,17'd12191,17'd6739,17'd71908,17'd63260,17'd1,17'd806,17'd20,17'd11,17'd16,17'd1415,17'd2597,17'd2597,17'd2597,17'd1414,17'd2596,17'd2597,17'd2597,17'd2596,17'd1414,17'd1414,17'd17,17'd19,17'd19,17'd10,17'd286,17'd27,17'd28,17'd28,17'd18037,17'd3754,17'd470,17'd470,17'd3431,17'd6278,17'd6746,17'd10408,17'd10672,17'd6441,17'd6904,17'd6747,17'd8048,17'd8198,17'd7390,17'd7063,17'd7063,17'd7392,17'd71093,17'd71909,17'd71910,17'd71911,17'd71912,17'd71913,17'd71914,17'd39815,17'd52378,17'd71818,17'd38096,17'd37975,17'd69448,17'd69448,17'd69448,17'd70891,17'd70085,17'd63559,17'd70989,17'd71915,17'd71915,17'd39055,17'd52785,17'd52552,17'd52552,17'd52552,17'd52474,17'd52552,17'd71327,17'd53086,17'd53086,17'd46489,17'd51771,17'd53376,17'd53168,17'd53169,17'd71627,17'd42795,17'd8376,17'd8541,17'd7755,17'd8070,17'd7421,17'd71627,17'd64809,17'd71819,17'd66456,17'd3780,17'd71916,17'd71917,17'd3480,17'd53523,17'd59012,17'd48081,17'd63841,17'd71918,17'd71919,17'd71920,17'd71921,17'd71730,17'd71922,17'd71923,17'd71924,17'd70615,17'd71734,17'd71925,17'd71926,17'd71453,17'd71738,17'd71927,17'd71928,17'd10293,17'd16044,17'd17582,17'd24844,17'd16181,17'd16047,17'd26857,17'd26858,17'd30359,17'd71929,17'd34949,17'd71930,17'd71931,17'd71932,17'd71933,17'd71934,17'd71935,17'd71936,17'd71937,17'd71938,17'd71939,17'd7296,17'd71940,17'd71941,17'd71942,17'd71943,17'd71944,17'd71945,17'd71946,17'd71947,17'd71948,17'd71949,17'd71950,17'd71951,17'd71952,17'd71953,17'd71954,17'd136,17'd132,17'd2698,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd133,17'd133,17'd1481,17'd132,17'd5593,17'd71036,17'd71955,17'd71956,17'd71957,17'd71958,17'd71863,17'd71864,17'd71959,17'd71960,17'd71961,17'd68812,17'd71489,17'd69681,17'd70645,17'd70845,17'd71165,17'd71681,17'd71870,17'd71962,17'd71778,17'd71873,17'd71166,17'd71493,17'd71782,17'd71686,17'd9381,17'd14040,17'd8627,17'd8627,17'd7996,17'd7833,17'd7497,17'd8610,17'd71495,17'd28649,17'd6386,17'd71963,17'd11573,17'd11430,17'd69787,17'd70649,17'd28305,17'd28305,17'd28305,17'd28305,17'd28183,17'd69692,17'd70650,17'd69029,17'd69969,17'd71389,17'd71499,17'd71785,17'd71964,17'd71965,17'd71966,17'd71881,17'd71967,17'd71968,17'd71969,17'd71970,17'd70956,17'd71971,17'd71972,17'd71973,17'd71974,17'd63357,17'd15733,17'd63789,17'd71975,17'd66073,17'd66676,17'd66072,17'd66318,17'd68519,17'd68519,17'd68944,17'd68182,17'd68182,17'd68182,17'd69797,17'd69797,17'd69797,17'd69797,17'd71976,17'd71977,17'd71978,17'd71977,17'd70861,17'd70861,17'd71891,17'd71892,17'd71405,17'd71182,17'd71893,17'd71893,17'd71405,17'd71405,17'd70571,17'd70472,17'd70470,17'd70861,17'd70666,17'd69524,17'd68519,17'd64919,17'd63243,17'd62851,17'd62850,17'd67426,17'd67426,17'd67426,17'd69342,17'd14734,17'd69342,17'd17179,17'd67163,17'd68741,17'd65688,17'd66064,17'd69237,17'd71979,17'd71896,17'd71410,17'd71980,17'd71897,17'd71700,17'd71898,17'd71413,17'd71414,17'd71609,17'd71899,17'd71981,17'd71982,17'd71982,17'd67672,17'd68632,17'd69424,17'd68632,17'd67438,17'd70477,17'd69039,17'd69039,17'd67437,17'd67437,17'd66320,17'd66320,17'd67296,17'd67296,17'd67051,17'd69800,17'd71300,17'd70269,17'd70162,17'd71286,17'd71302,17'd71983,17'd60030,17'd58990,17'd2906,17'd5940,17'd5371,17'd3743,17'd1396,17'd1396,17'd1243,17'd259,17'd206,17'd643,17'd1124,17'd1124,17'd205,17'd424,17'd1381,17'd1381,17'd1382,17'd1382,17'd603,17'd952,17'd204,17'd71984
},
'{
17'd3903,17'd4244,17'd4087,17'd4426,17'd4735,17'd5201,17'd5202,17'd9959,17'd4427,17'd5646,17'd5646,17'd4087,17'd5202,17'd5201,17'd71985,17'd71986,17'd71987,17'd71194,17'd63976,17'd63976,17'd71988,17'd71989,17'd71990,17'd71990,17'd70070,17'd63979,17'd69723,17'd71424,17'd3250,17'd9815,17'd12503,17'd67576,17'd65712,17'd71713,17'd6895,17'd67305,17'd64537,17'd71713,17'd66210,17'd66207,17'd66444,17'd66814,17'd71991,17'd69350,17'd71992,17'd9674,17'd71618,17'd65841,17'd10660,17'd70977,17'd65583,17'd67574,17'd6735,17'd13065,17'd15,17'd1275,17'd20,17'd21,17'd1128,17'd1416,17'd1414,17'd2597,17'd2258,17'd2597,17'd2596,17'd2596,17'd2597,17'd2597,17'd1414,17'd1414,17'd1416,17'd4089,17'd19,17'd979,17'd808,17'd808,17'd287,17'd28,17'd288,17'd2118,17'd1693,17'd469,17'd3254,17'd5208,17'd5803,17'd6439,17'd10672,17'd6440,17'd6904,17'd9970,17'd9970,17'd7063,17'd8198,17'd8198,17'd8198,17'd7227,17'd70880,17'd71430,17'd71993,17'd68203,17'd71994,17'd71995,17'd71996,17'd71997,17'd52475,17'd52114,17'd70086,17'd70700,17'd38888,17'd71103,17'd71103,17'd69549,17'd70085,17'd7424,17'd7424,17'd69062,17'd71998,17'd71998,17'd39199,17'd39055,17'd71106,17'd70793,17'd70793,17'd71106,17'd68656,17'd68656,17'd49611,17'd39647,17'd53087,17'd71999,17'd53168,17'd6937,17'd7097,17'd7253,17'd8375,17'd8070,17'd8375,17'd8070,17'd7916,17'd71108,17'd71108,17'd72000,17'd72001,17'd68539,17'd72002,17'd72003,17'd72004,17'd63999,17'd72005,17'd13467,17'd6464,17'd72006,17'd72007,17'd72008,17'd71921,17'd72009,17'd72010,17'd72011,17'd71924,17'd70615,17'd72012,17'd72013,17'd72014,17'd71234,17'd71738,17'd71928,17'd11364,17'd10293,17'd9709,17'd17582,17'd72015,17'd25130,17'd26987,17'd9994,17'd72016,17'd72017,17'd71742,17'd35081,17'd7599,17'd72018,17'd72019,17'd43359,17'd38232,17'd72020,17'd72021,17'd72022,17'd71754,17'd72023,17'd72024,17'd72025,17'd72026,17'd72027,17'd72028,17'd72029,17'd72030,17'd71945,17'd72031,17'd72032,17'd72033,17'd72034,17'd72035,17'd72036,17'd71953,17'd72037,17'd20762,17'd130,17'd132,17'd135,17'd134,17'd132,17'd132,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd133,17'd133,17'd1481,17'd130,17'd132,17'd72038,17'd72039,17'd72040,17'd72041,17'd72042,17'd72043,17'd72044,17'd72045,17'd72046,17'd72047,17'd68919,17'd71489,17'd69403,17'd72048,17'd72049,17'd72050,17'd71165,17'd72051,17'd72052,17'd72053,17'd72054,17'd71780,17'd72055,17'd72056,17'd70850,17'd9381,17'd71783,17'd8627,17'd8627,17'd14037,17'd7498,17'd10362,17'd8454,17'd9068,17'd72057,17'd6385,17'd11572,17'd11180,17'd11430,17'd69787,17'd70649,17'd28534,17'd28534,17'd28534,17'd28183,17'd68510,17'd69692,17'd72058,17'd68931,17'd69512,17'd71389,17'd72059,17'd72060,17'd72061,17'd72062,17'd72063,17'd72064,17'd72065,17'd72066,17'd71969,17'd72067,17'd72068,17'd72069,17'd72070,17'd72071,17'd27941,17'd14580,17'd64509,17'd72072,17'd66678,17'd63244,17'd66676,17'd66437,17'd66072,17'd66318,17'd66928,17'd70259,17'd66928,17'd68519,17'd68519,17'd68519,17'd68519,17'd68519,17'd68519,17'd69706,17'd69797,17'd71976,17'd71976,17'd71976,17'd71976,17'd70581,17'd70581,17'd72073,17'd72074,17'd72074,17'd72074,17'd72074,17'd70675,17'd70770,17'd70770,17'd70770,17'd70675,17'd71302,17'd69706,17'd69337,17'd63807,17'd65950,17'd68834,17'd68834,17'd15483,17'd15999,17'd69342,17'd69342,17'd70963,17'd67425,17'd68836,17'd66322,17'd72075,17'd68736,17'd69142,17'd69037,17'd71979,17'd69036,17'd72076,17'd71980,17'd72077,17'd72078,17'd71898,17'd71413,17'd71414,17'd71609,17'd72079,17'd72080,17'd71982,17'd68837,17'd69147,17'd69147,17'd67672,17'd67673,17'd69039,17'd69039,17'd67437,17'd67437,17'd66320,17'd66320,17'd66320,17'd67296,17'd67439,17'd67439,17'd67296,17'd69711,17'd71610,17'd70059,17'd69703,17'd69524,17'd72081,17'd71420,17'd36903,17'd11882,17'd9123,17'd5371,17'd5050,17'd3743,17'd1823,17'd1396,17'd259,17'd259,17'd206,17'd206,17'd1124,17'd1828,17'd971,17'd1272,17'd1245,17'd202,17'd202,17'd422,17'd603,17'd424,17'd205,17'd1966
},
'{
17'd9960,17'd3903,17'd4427,17'd4426,17'd5201,17'd5201,17'd5202,17'd9959,17'd4736,17'd4426,17'd5646,17'd4087,17'd5202,17'd4735,17'd5377,17'd72082,17'd72083,17'd71905,17'd63975,17'd63976,17'd72084,17'd72085,17'd72086,17'd72087,17'd65449,17'd66693,17'd12928,17'd70778,17'd6265,17'd7371,17'd12503,17'd63519,17'd71708,17'd67816,17'd7052,17'd6739,17'd64120,17'd69050,17'd8663,17'd69722,17'd70071,17'd66331,17'd72088,17'd71090,17'd69722,17'd8817,17'd9130,17'd72089,17'd72090,17'd72091,17'd68645,17'd65583,17'd13576,17'd65189,17'd64125,17'd1,17'd20,17'd21,17'd20,17'd20404,17'd17,17'd2596,17'd2258,17'd2597,17'd2596,17'd2596,17'd2596,17'd2597,17'd2257,17'd1414,17'd1414,17'd17,17'd18,17'd19,17'd10,17'd10,17'd28,17'd652,17'd29,17'd288,17'd31,17'd1129,17'd3254,17'd3255,17'd6278,17'd11211,17'd70077,17'd10672,17'd6904,17'd6904,17'd9970,17'd7227,17'd70687,17'd70687,17'd8048,17'd7063,17'd71092,17'd72092,17'd72093,17'd72094,17'd72095,17'd72096,17'd72097,17'd72098,17'd70889,17'd38094,17'd70295,17'd69062,17'd52785,17'd52205,17'd38095,17'd71435,17'd70086,17'd70700,17'd70085,17'd70085,17'd70891,17'd70891,17'd38888,17'd38888,17'd71106,17'd68860,17'd72099,17'd68860,17'd68860,17'd63559,17'd70989,17'd72100,17'd72101,17'd72102,17'd72101,17'd66954,17'd7421,17'd7089,17'd68437,17'd8375,17'd8376,17'd8375,17'd8376,17'd71108,17'd72103,17'd72104,17'd72105,17'd72106,17'd68654,17'd64941,17'd59265,17'd58644,17'd8539,17'd5090,17'd72107,17'd72108,17'd72109,17'd72008,17'd72110,17'd72111,17'd72112,17'd72011,17'd70614,17'd71549,17'd72113,17'd72114,17'd72115,17'd71643,17'd71834,17'd72116,17'd11364,17'd10293,17'd16891,17'd16667,17'd16782,17'd25131,17'd15787,17'd72117,17'd72118,17'd8393,17'd72119,17'd72120,17'd72121,17'd72122,17'd72123,17'd72124,17'd72125,17'd72126,17'd72127,17'd72128,17'd72129,17'd72130,17'd72131,17'd72132,17'd72133,17'd71025,17'd72134,17'd72135,17'd72136,17'd72137,17'd72138,17'd72139,17'd72140,17'd72141,17'd72142,17'd72143,17'd71953,17'd70742,17'd20762,17'd130,17'd132,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd133,17'd133,17'd1481,17'd132,17'd5593,17'd72144,17'd72145,17'd72146,17'd72147,17'd26692,17'd72148,17'd72044,17'd72045,17'd72149,17'd72150,17'd68919,17'd71489,17'd72151,17'd69682,17'd72049,17'd72050,17'd71049,17'd72152,17'd72153,17'd72154,17'd72054,17'd71780,17'd71683,17'd72155,17'd70850,17'd9381,17'd71783,17'd8627,17'd8627,17'd13673,17'd7498,17'd10362,17'd8455,17'd7992,17'd72057,17'd6385,17'd71963,17'd11573,17'd11430,17'd69787,17'd70649,17'd28534,17'd28534,17'd28534,17'd28305,17'd28183,17'd69692,17'd72058,17'd68825,17'd70364,17'd72156,17'd72157,17'd72158,17'd72159,17'd72160,17'd72161,17'd72064,17'd72065,17'd72162,17'd72163,17'd71792,17'd71176,17'd69608,17'd72164,17'd72165,17'd14579,17'd23292,17'd14172,17'd65042,17'd66536,17'd63376,17'd63964,17'd66073,17'd66073,17'd66072,17'd66437,17'd66928,17'd66318,17'd66318,17'd66318,17'd66318,17'd66928,17'd68519,17'd68519,17'd68519,17'd68182,17'd68182,17'd68182,17'd69797,17'd69797,17'd71976,17'd69798,17'd70581,17'd70581,17'd70581,17'd70581,17'd70581,17'd69798,17'd69523,17'd69523,17'd69705,17'd71302,17'd70482,17'd68944,17'd68520,17'd65950,17'd67435,17'd15483,17'd15483,17'd15483,17'd15999,17'd69342,17'd70963,17'd67425,17'd68836,17'd66322,17'd71798,17'd64903,17'd65038,17'd72166,17'd67550,17'd69036,17'd72167,17'd72168,17'd71980,17'd72077,17'd72078,17'd72169,17'd71414,17'd71609,17'd71981,17'd72170,17'd72171,17'd72172,17'd68837,17'd69147,17'd68837,17'd67672,17'd67673,17'd69039,17'd69039,17'd67437,17'd70477,17'd66320,17'd66320,17'd66320,17'd67296,17'd67439,17'd67439,17'd66320,17'd70773,17'd70966,17'd70162,17'd69703,17'd70482,17'd71802,17'd63652,17'd35487,17'd2906,17'd5940,17'd5371,17'd3743,17'd3743,17'd1396,17'd1666,17'd259,17'd260,17'd206,17'd206,17'd1124,17'd972,17'd424,17'd1272,17'd1382,17'd202,17'd1382,17'd1382,17'd952,17'd204,17'd205,17'd205
},
'{
17'd3904,17'd4088,17'd3903,17'd3902,17'd4087,17'd4087,17'd5202,17'd9959,17'd4736,17'd4426,17'd4426,17'd4087,17'd5202,17'd4735,17'd5645,17'd5377,17'd71986,17'd71987,17'd72173,17'd72174,17'd71423,17'd72085,17'd71423,17'd71906,17'd65714,17'd72175,17'd63979,17'd63820,17'd11887,17'd2784,17'd64400,17'd12503,17'd65067,17'd64929,17'd6739,17'd69161,17'd64537,17'd68848,17'd67815,17'd72176,17'd72177,17'd72178,17'd71090,17'd72179,17'd67450,17'd9547,17'd8662,17'd72180,17'd13576,17'd6894,17'd8043,17'd65583,17'd70070,17'd13433,17'd12783,17'd1830,17'd806,17'd2933,17'd21,17'd20,17'd18,17'd1416,17'd2597,17'd2596,17'd2596,17'd1414,17'd2596,17'd2597,17'd2597,17'd2257,17'd1414,17'd17,17'd3905,17'd18,17'd11,17'd10,17'd27,17'd980,17'd652,17'd29,17'd4091,17'd3595,17'd3254,17'd3254,17'd3756,17'd11889,17'd11211,17'd10408,17'd6904,17'd6904,17'd10409,17'd7391,17'd70688,17'd70687,17'd8048,17'd8048,17'd7560,17'd72181,17'd72182,17'd67578,17'd72183,17'd72184,17'd72185,17'd72186,17'd72187,17'd70495,17'd72188,17'd72189,17'd6783,17'd70792,17'd38222,17'd38220,17'd38096,17'd37975,17'd70086,17'd70986,17'd38219,17'd38219,17'd70086,17'd70086,17'd70891,17'd69996,17'd63421,17'd69548,17'd69548,17'd72190,17'd70294,17'd72191,17'd68433,17'd68433,17'd68433,17'd66953,17'd7916,17'd8541,17'd5085,17'd68437,17'd42795,17'd7097,17'd72192,17'd72193,17'd72194,17'd72195,17'd72196,17'd72197,17'd65861,17'd72198,17'd61695,17'd64944,17'd5836,17'd72199,17'd34683,17'd72200,17'd72201,17'd72202,17'd72203,17'd72204,17'd72205,17'd72206,17'd71639,17'd71831,17'd72207,17'd72208,17'd72209,17'd72210,17'd72211,17'd10293,17'd10293,17'd10293,17'd9588,17'd16781,17'd72212,17'd15658,17'd72213,17'd72214,17'd54450,17'd72215,17'd72216,17'd7599,17'd72217,17'd72218,17'd72219,17'd72220,17'd72221,17'd72222,17'd72223,17'd72224,17'd72225,17'd72226,17'd72227,17'd72228,17'd72229,17'd72230,17'd72231,17'd72232,17'd72233,17'd72234,17'd72235,17'd72236,17'd72237,17'd72238,17'd72239,17'd72240,17'd72241,17'd72242,17'd137,17'd128,17'd132,17'd132,17'd130,17'd1481,17'd356,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd132,17'd130,17'd130,17'd130,17'd1481,17'd133,17'd133,17'd134,17'd132,17'd7649,17'd72243,17'd72244,17'd72245,17'd72246,17'd40073,17'd25758,17'd72044,17'd72247,17'd72248,17'd72249,17'd68919,17'd71489,17'd69966,17'd72048,17'd70845,17'd72050,17'd72050,17'd72250,17'd71962,17'd72251,17'd72054,17'd72252,17'd72253,17'd72155,17'd9515,17'd19588,17'd13795,17'd9237,17'd9237,17'd13673,17'd7498,17'd72254,17'd8455,17'd7992,17'd72057,17'd6385,17'd11572,17'd11180,17'd11430,17'd69787,17'd70649,17'd28534,17'd28534,17'd28534,17'd28305,17'd10642,17'd10516,17'd72255,17'd68724,17'd70364,17'd72156,17'd72157,17'd72158,17'd72256,17'd72257,17'd72258,17'd72259,17'd72260,17'd72261,17'd72262,17'd71693,17'd72263,17'd72264,17'd72265,17'd72266,17'd72267,17'd13929,17'd18266,17'd65288,17'd65553,17'd72268,17'd72269,17'd65951,17'd63808,17'd66676,17'd66437,17'd66072,17'd66072,17'd66072,17'd66072,17'd66072,17'd66072,17'd66318,17'd66318,17'd66928,17'd66318,17'd68944,17'd68944,17'd68944,17'd68519,17'd69706,17'd69706,17'd72270,17'd71302,17'd70582,17'd70582,17'd70482,17'd70482,17'd70570,17'd70469,17'd70469,17'd70662,17'd72271,17'd68833,17'd63962,17'd62849,17'd15483,17'd15232,17'd67557,17'd69342,17'd69342,17'd70963,17'd67425,17'd68836,17'd68741,17'd70166,17'd72272,17'd65038,17'd71409,17'd71295,17'd71410,17'd72167,17'd72167,17'd72168,17'd72273,17'd72077,17'd72078,17'd72274,17'd72275,17'd71801,17'd72276,17'd72171,17'd72277,17'd68837,17'd71190,17'd68837,17'd68947,17'd71901,17'd68738,17'd69039,17'd69039,17'd67296,17'd66320,17'd70773,17'd70773,17'd70478,17'd72278,17'd67296,17'd67296,17'd70773,17'd71299,17'd70966,17'd70261,17'd69524,17'd72270,17'd65564,17'd36903,17'd9261,17'd6416,17'd4729,17'd229,17'd3743,17'd1396,17'd644,17'd643,17'd260,17'd260,17'd206,17'd643,17'd205,17'd972,17'd1244,17'd1381,17'd1382,17'd1382,17'd1382,17'd202,17'd424,17'd205,17'd1687,17'd1828
},
'{
17'd6264,17'd3904,17'd4088,17'd4244,17'd4087,17'd4087,17'd5202,17'd5202,17'd4427,17'd4426,17'd5646,17'd4426,17'd5202,17'd4735,17'd5645,17'd5645,17'd72082,17'd72279,17'd71309,17'd72280,17'd72280,17'd71518,17'd71518,17'd65715,17'd72281,17'd65714,17'd65449,17'd66693,17'd63666,17'd6424,17'd9815,17'd9815,17'd71709,17'd65066,17'd64254,17'd6894,17'd66815,17'd64119,17'd65581,17'd8515,17'd8513,17'd71426,17'd69808,17'd71617,17'd65959,17'd66210,17'd8976,17'd8975,17'd13064,17'd13576,17'd12033,17'd67574,17'd65449,17'd64254,17'd11607,17'd64125,17'd1,17'd806,17'd20,17'd20,17'd11,17'd17,17'd2597,17'd2596,17'd1414,17'd1414,17'd2596,17'd2596,17'd2597,17'd2597,17'd1414,17'd17187,17'd17,17'd18,17'd19,17'd11,17'd27,17'd27,17'd652,17'd28,17'd4248,17'd3908,17'd3433,17'd3254,17'd3434,17'd11210,17'd72282,17'd70077,17'd6904,17'd6904,17'd9970,17'd10409,17'd70688,17'd70687,17'd8198,17'd8048,17'd7560,17'd70389,17'd72283,17'd72284,17'd61290,17'd72285,17'd72286,17'd72287,17'd72288,17'd72289,17'd72290,17'd72290,17'd72291,17'd6784,17'd38222,17'd72292,17'd38220,17'd38480,17'd38096,17'd38219,17'd38219,17'd38219,17'd70986,17'd70986,17'd69996,17'd69996,17'd69548,17'd72190,17'd72293,17'd65213,17'd72294,17'd72294,17'd70702,17'd68540,17'd69263,17'd72295,17'd72295,17'd72296,17'd64813,17'd8541,17'd71108,17'd72297,17'd72195,17'd72298,17'd72298,17'd72299,17'd72300,17'd72301,17'd72302,17'd72303,17'd72304,17'd72305,17'd69731,17'd72306,17'd72307,17'd72308,17'd72309,17'd72310,17'd72311,17'd72312,17'd71547,17'd71125,17'd72313,17'd72314,17'd72315,17'd72316,17'd72317,17'd10295,17'd8856,17'd9167,17'd9167,17'd10129,17'd9589,17'd16180,17'd16418,17'd25805,17'd72318,17'd72319,17'd53175,17'd72320,17'd37979,17'd72321,17'd72322,17'd72323,17'd72324,17'd6962,17'd72325,17'd6665,17'd72326,17'd72327,17'd72225,17'd72328,17'd72329,17'd72330,17'd72331,17'd72332,17'd72029,17'd72333,17'd72334,17'd72335,17'd72336,17'd72337,17'd72338,17'd72339,17'd72340,17'd72341,17'd72342,17'd72343,17'd137,17'd139,17'd130,17'd132,17'd130,17'd4163,17'd4163,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd132,17'd130,17'd130,17'd1481,17'd133,17'd133,17'd134,17'd131,17'd11821,17'd72344,17'd72345,17'd72346,17'd72246,17'd23961,17'd19578,17'd72347,17'd72247,17'd72348,17'd72349,17'd68919,17'd72350,17'd72351,17'd72352,17'd70845,17'd72050,17'd72353,17'd72354,17'd72355,17'd72054,17'd72054,17'd72252,17'd72356,17'd10216,17'd9515,17'd19588,17'd13795,17'd9237,17'd9237,17'd13673,17'd8470,17'd7664,17'd8455,17'd7992,17'd72057,17'd6385,17'd71963,17'd11573,17'd11430,17'd69787,17'd70649,17'd28305,17'd28534,17'd28305,17'd28305,17'd10642,17'd9933,17'd31718,17'd68724,17'd69129,17'd72357,17'd72157,17'd72158,17'd72358,17'd72359,17'd72360,17'd72259,17'd72260,17'd72361,17'd71968,17'd71791,17'd72362,17'd70257,17'd70659,17'd72363,17'd72364,17'd72365,17'd22771,17'd64509,17'd64090,17'd66306,17'd72268,17'd71508,17'd63378,17'd63964,17'd66676,17'd66072,17'd66072,17'd66072,17'd66072,17'd66072,17'd66072,17'd66072,17'd66072,17'd66318,17'd66318,17'd66318,17'd66318,17'd66318,17'd66318,17'd68944,17'd68519,17'd69706,17'd69705,17'd70482,17'd70482,17'd69705,17'd70570,17'd70469,17'd70857,17'd70857,17'd69338,17'd68520,17'd63962,17'd62849,17'd16959,17'd67426,17'd67557,17'd67557,17'd14734,17'd69342,17'd67425,17'd68836,17'd70373,17'd72075,17'd65421,17'd64766,17'd71409,17'd67663,17'd72076,17'd72076,17'd72076,17'd72168,17'd72366,17'd72273,17'd72077,17'd72367,17'd72368,17'd72369,17'd72276,17'd72171,17'd72370,17'd72371,17'd71076,17'd71190,17'd68837,17'd68947,17'd71901,17'd68738,17'd69039,17'd69039,17'd67296,17'd67295,17'd70773,17'd69711,17'd70478,17'd72278,17'd67296,17'd69711,17'd71417,17'd70966,17'd70162,17'd69703,17'd70482,17'd72372,17'd60030,17'd36903,17'd8187,17'd4882,17'd3895,17'd1261,17'd1262,17'd1666,17'd643,17'd206,17'd260,17'd260,17'd206,17'd643,17'd205,17'd971,17'd1244,17'd1381,17'd202,17'd422,17'd422,17'd203,17'd204,17'd205,17'd1828,17'd1410
},
'{
17'd4887,17'd4733,17'd4088,17'd3903,17'd4427,17'd4087,17'd4087,17'd4087,17'd4736,17'd4087,17'd4426,17'd4426,17'd5201,17'd5201,17'd5201,17'd5645,17'd5791,17'd72373,17'd72374,17'd72375,17'd72376,17'd72377,17'd72378,17'd72379,17'd72380,17'd72281,17'd65712,17'd66815,17'd63978,17'd72381,17'd2781,17'd3249,17'd63257,17'd70972,17'd64798,17'd72382,17'd11885,17'd65449,17'd64396,17'd67574,17'd7220,17'd8512,17'd72383,17'd70285,17'd70975,17'd69809,17'd9127,17'd11447,17'd6737,17'd64254,17'd13576,17'd11885,17'd70070,17'd66693,17'd70178,17'd12783,17'd63118,17'd1,17'd806,17'd8814,17'd1128,17'd4089,17'd1414,17'd2596,17'd2257,17'd1416,17'd1415,17'd1414,17'd2597,17'd2597,17'd1414,17'd1415,17'd17,17'd18,17'd19,17'd19,17'd27,17'd27,17'd27,17'd27,17'd27444,17'd4248,17'd3595,17'd3254,17'd3431,17'd12335,17'd10269,17'd10093,17'd6904,17'd6600,17'd6747,17'd7227,17'd7560,17'd7560,17'd8198,17'd70687,17'd7391,17'd70077,17'd72384,17'd72385,17'd72386,17'd72387,17'd72388,17'd72389,17'd72390,17'd72391,17'd72392,17'd62122,17'd72393,17'd6784,17'd6784,17'd38095,17'd38220,17'd38220,17'd38095,17'd71103,17'd69360,17'd69549,17'd70295,17'd70295,17'd69997,17'd69997,17'd39054,17'd70082,17'd72394,17'd72394,17'd72395,17'd72395,17'd69547,17'd72396,17'd72396,17'd72397,17'd72398,17'd72399,17'd72400,17'd72401,17'd72402,17'd72403,17'd72404,17'd72404,17'd72405,17'd72406,17'd72407,17'd72408,17'd72409,17'd72410,17'd72411,17'd72412,17'd72413,17'd72414,17'd72415,17'd72416,17'd72417,17'd72418,17'd72419,17'd72420,17'd72421,17'd70614,17'd72422,17'd58549,17'd62244,17'd72423,17'd71454,17'd72424,17'd9167,17'd9167,17'd8856,17'd9315,17'd9993,17'd16295,17'd26483,17'd72425,17'd9024,17'd7768,17'd72426,17'd72427,17'd72428,17'd72217,17'd72429,17'd72430,17'd72431,17'd72432,17'd72433,17'd72434,17'd72435,17'd70734,17'd72436,17'd72436,17'd72437,17'd72438,17'd72439,17'd72440,17'd72441,17'd72333,17'd72442,17'd72443,17'd72444,17'd72445,17'd72446,17'd72447,17'd72448,17'd72449,17'd72342,17'd72242,17'd137,17'd127,17'd130,17'd132,17'd356,17'd70217,17'd70217,17'd70438,17'd1481,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd131,17'd132,17'd132,17'd130,17'd130,17'd133,17'd133,17'd134,17'd132,17'd11683,17'd72450,17'd72451,17'd72452,17'd72453,17'd72454,17'd19699,17'd72455,17'd72247,17'd72348,17'd72349,17'd68919,17'd72350,17'd70754,17'd69322,17'd71868,17'd72050,17'd72353,17'd72354,17'd72355,17'd72054,17'd72456,17'd72457,17'd72253,17'd72458,17'd70053,17'd19588,17'd13795,17'd9237,17'd9237,17'd9088,17'd7173,17'd72254,17'd8455,17'd7992,17'd72057,17'd6385,17'd11572,17'd11180,17'd11430,17'd69787,17'd70649,17'd28305,17'd28534,17'd11181,17'd11181,17'd10642,17'd9933,17'd57865,17'd70650,17'd69029,17'd72459,17'd72460,17'd72158,17'd72461,17'd72359,17'd72462,17'd72463,17'd72260,17'd72361,17'd72162,17'd71692,17'd72464,17'd72465,17'd72466,17'd72467,17'd72468,17'd28421,17'd18029,17'd64509,17'd63639,17'd63789,17'd66306,17'd71596,17'd63376,17'd63964,17'd63964,17'd66073,17'd66073,17'd66073,17'd66073,17'd66073,17'd66073,17'd66072,17'd66072,17'd66072,17'd65054,17'd65054,17'd65054,17'd65054,17'd66072,17'd66318,17'd66318,17'd68944,17'd69337,17'd69885,17'd69885,17'd69885,17'd72271,17'd70061,17'd68833,17'd68833,17'd63962,17'd66197,17'd68834,17'd17179,17'd67427,17'd62449,17'd62449,17'd62449,17'd62854,17'd65705,17'd66322,17'd68416,17'd72469,17'd65686,17'd66062,17'd67788,17'd67663,17'd72470,17'd72471,17'd72366,17'd72366,17'd72472,17'd72472,17'd72273,17'd72473,17'd72474,17'd72475,17'd72369,17'd72476,17'd72477,17'd72478,17'd69147,17'd71076,17'd71190,17'd67672,17'd67673,17'd71901,17'd68738,17'd67674,17'd66076,17'd67296,17'd66320,17'd70773,17'd69711,17'd72278,17'd72479,17'd67296,17'd70773,17'd70867,17'd70868,17'd70163,17'd69523,17'd72081,17'd64917,17'd36903,17'd12923,17'd5958,17'd3897,17'd1119,17'd1262,17'd1262,17'd970,17'd206,17'd1829,17'd206,17'd206,17'd643,17'd644,17'd972,17'd1685,17'd1381,17'd1382,17'd202,17'd422,17'd1382,17'd2256,17'd205,17'd972,17'd645,17'd458
},
'{
17'd4577,17'd4887,17'd4733,17'd4088,17'd3903,17'd4427,17'd4087,17'd4087,17'd7042,17'd4736,17'd4087,17'd4426,17'd5201,17'd5201,17'd5201,17'd4735,17'd5053,17'd72480,17'd72481,17'd72482,17'd72483,17'd72484,17'd72485,17'd72486,17'd72487,17'd72488,17'd72489,17'd68751,17'd67305,17'd66333,17'd2781,17'd1689,17'd3750,17'd70076,17'd71086,17'd72490,17'd68645,17'd65583,17'd71708,17'd71195,17'd6896,17'd7378,17'd72176,17'd69250,17'd67946,17'd68313,17'd8975,17'd11447,17'd8343,17'd13064,17'd64254,17'd13064,17'd13576,17'd64397,17'd64666,17'd70178,17'd10923,17'd63118,17'd3,17'd806,17'd1128,17'd3905,17'd1414,17'd1414,17'd22965,17'd1416,17'd1415,17'd1414,17'd2596,17'd2597,17'd1414,17'd1414,17'd17,17'd16,17'd18,17'd19,17'd27,17'd27,17'd27,17'd27,17'd20570,17'd27444,17'd3755,17'd3431,17'd2942,17'd12036,17'd11210,17'd10093,17'd9970,17'd6600,17'd6747,17'd6747,17'd7063,17'd7390,17'd8198,17'd70687,17'd10409,17'd70077,17'd68854,17'd72491,17'd72492,17'd60897,17'd72493,17'd72494,17'd72495,17'd72496,17'd72497,17'd72498,17'd72499,17'd69168,17'd69360,17'd69360,17'd38220,17'd38484,17'd38095,17'd38095,17'd71103,17'd69549,17'd70295,17'd70295,17'd69817,17'd69817,17'd39054,17'd70185,17'd63708,17'd63708,17'd72394,17'd72500,17'd72501,17'd72502,17'd72503,17'd72504,17'd72505,17'd72408,17'd72506,17'd72507,17'd72405,17'd72508,17'd72509,17'd72510,17'd72511,17'd72512,17'd72413,17'd72513,17'd72514,17'd32267,17'd72515,17'd72512,17'd72516,17'd72517,17'd72518,17'd72519,17'd72520,17'd72521,17'd71733,17'd72522,17'd71638,17'd71549,17'd58549,17'd72115,17'd62124,17'd72523,17'd72524,17'd72424,17'd9167,17'd9167,17'd10129,17'd9315,17'd16180,17'd25660,17'd9994,17'd72318,17'd72525,17'd53175,17'd72526,17'd38744,17'd72527,17'd72528,17'd72529,17'd72530,17'd72531,17'd72532,17'd72533,17'd72534,17'd72535,17'd72536,17'd72436,17'd72537,17'd72538,17'd72539,17'd72540,17'd72541,17'd72542,17'd72543,17'd72544,17'd72545,17'd72546,17'd72547,17'd72548,17'd72549,17'd72550,17'd72551,17'd71033,17'd72242,17'd72552,17'd138,17'd130,17'd130,17'd72553,17'd70744,17'd70217,17'd70438,17'd1481,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd130,17'd130,17'd133,17'd132,17'd132,17'd131,17'd5593,17'd72554,17'd72555,17'd72556,17'd72557,17'd23611,17'd19971,17'd72558,17'd72247,17'd72348,17'd72249,17'd68919,17'd71270,17'd72151,17'd72352,17'd70756,17'd72559,17'd72353,17'd72560,17'd72561,17'd72562,17'd72456,17'd72563,17'd72564,17'd72565,17'd8774,17'd19588,17'd13795,17'd9391,17'd9087,17'd9088,17'd7174,17'd7664,17'd7993,17'd7992,17'd72057,17'd6385,17'd71963,17'd11573,17'd11430,17'd69787,17'd69787,17'd28305,17'd28305,17'd11181,17'd11181,17'd10515,17'd9933,17'd57865,17'd72566,17'd69029,17'd72567,17'd72568,17'd72569,17'd72570,17'd72159,17'd71879,17'd71966,17'd72571,17'd72572,17'd72573,17'd71882,17'd72574,17'd72575,17'd72576,17'd72577,17'd72578,17'd72579,17'd13929,17'd17177,17'd63495,17'd63640,17'd63789,17'd65040,17'd65286,17'd63378,17'd67440,17'd63808,17'd63808,17'd66073,17'd66073,17'd66073,17'd66073,17'd66073,17'd66072,17'd66072,17'd65054,17'd65054,17'd65054,17'd65054,17'd65054,17'd65054,17'd66072,17'd66318,17'd66319,17'd68944,17'd68944,17'd68944,17'd70061,17'd69145,17'd68520,17'd64387,17'd66197,17'd62851,17'd65571,17'd65705,17'd69146,17'd62976,17'd62976,17'd69146,17'd68742,17'd16255,17'd65816,17'd65040,17'd65686,17'd72580,17'd67788,17'd71410,17'd72581,17'd68516,17'd72471,17'd72366,17'd72273,17'd72472,17'd72472,17'd72273,17'd72474,17'd72582,17'd72583,17'd72584,17'd72585,17'd72172,17'd69147,17'd71076,17'd72586,17'd71190,17'd67672,17'd67673,17'd71901,17'd68738,17'd67674,17'd66076,17'd66320,17'd66320,17'd69711,17'd70478,17'd72278,17'd72278,17'd66320,17'd70773,17'd70867,17'd70163,17'd69524,17'd72270,17'd65564,17'd60030,17'd11882,17'd9544,17'd4575,17'd2586,17'd625,17'd625,17'd1962,17'd259,17'd2779,17'd1829,17'd206,17'd206,17'd643,17'd644,17'd971,17'd1272,17'd202,17'd1382,17'd202,17'd1382,17'd202,17'd13940,17'd205,17'd1410,17'd274,17'd272
},
'{
17'd4577,17'd4577,17'd6584,17'd3904,17'd9960,17'd4244,17'd4087,17'd4087,17'd4736,17'd4736,17'd4427,17'd4426,17'd4426,17'd4426,17'd5201,17'd4735,17'd10532,17'd72587,17'd72588,17'd72589,17'd72590,17'd72591,17'd72592,17'd72593,17'd72485,17'd72594,17'd65717,17'd71427,17'd65583,17'd71310,17'd10668,17'd1127,17'd1689,17'd9684,17'd71085,17'd64665,17'd72595,17'd12330,17'd64254,17'd64122,17'd6739,17'd6895,17'd8513,17'd72177,17'd70975,17'd9675,17'd70977,17'd72596,17'd7053,17'd6737,17'd13576,17'd63979,17'd6740,17'd64254,17'd66693,17'd13815,17'd64667,17'd65314,17'd3749,17'd283,17'd1128,17'd18,17'd17,17'd1414,17'd22965,17'd1416,17'd1414,17'd1415,17'd2596,17'd2596,17'd1414,17'd2257,17'd1416,17'd17,17'd18,17'd19,17'd27,17'd27,17'd27,17'd27,17'd20570,17'd6745,17'd3907,17'd11208,17'd12654,17'd12036,17'd3754,17'd6598,17'd6600,17'd7389,17'd72597,17'd69437,17'd6749,17'd6906,17'd7559,17'd7390,17'd7731,17'd7562,17'd9817,17'd72598,17'd72599,17'd68315,17'd72600,17'd72601,17'd72602,17'd72603,17'd72604,17'd72605,17'd72606,17'd71626,17'd69448,17'd38219,17'd37973,17'd38222,17'd38222,17'd38222,17'd71103,17'd69549,17'd69733,17'd69733,17'd72607,17'd63421,17'd70083,17'd72608,17'd63296,17'd63296,17'd63296,17'd72609,17'd63858,17'd72610,17'd72610,17'd72611,17'd72612,17'd72613,17'd72614,17'd72510,17'd72510,17'd72509,17'd72615,17'd72616,17'd37319,17'd36334,17'd34528,17'd72617,17'd32903,17'd72618,17'd72616,17'd72619,17'd72620,17'd72621,17'd72622,17'd72623,17'd72624,17'd70417,17'd72520,17'd72625,17'd70812,17'd72314,17'd72115,17'd71234,17'd72626,17'd72627,17'd72628,17'd72424,17'd9167,17'd10293,17'd10129,17'd72629,17'd27464,17'd10436,17'd15024,17'd12541,17'd8707,17'd72630,17'd72631,17'd72632,17'd40433,17'd72633,17'd72634,17'd6962,17'd72635,17'd72533,17'd72534,17'd72636,17'd72637,17'd72638,17'd72639,17'd72640,17'd72641,17'd72642,17'd72031,17'd72643,17'd72644,17'd72645,17'd72646,17'd72647,17'd72648,17'd72649,17'd72650,17'd72651,17'd72652,17'd72653,17'd72654,17'd72655,17'd71477,17'd137,17'd130,17'd72656,17'd72657,17'd72658,17'd127,17'd70438,17'd356,17'd1481,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd132,17'd131,17'd11683,17'd72659,17'd72660,17'd72661,17'd72662,17'd19829,17'd20356,17'd72558,17'd72663,17'd72248,17'd72150,17'd68919,17'd71270,17'd71588,17'd69217,17'd70756,17'd72559,17'd71049,17'd72560,17'd72664,17'd72665,17'd72456,17'd72563,17'd72666,17'd72667,17'd72155,17'd19588,17'd13795,17'd9391,17'd9087,17'd9088,17'd7173,17'd20245,17'd7993,17'd7992,17'd72668,17'd11849,17'd11572,17'd11180,17'd11430,17'd71784,17'd69787,17'd11181,17'd11181,17'd11181,17'd11181,17'd10514,17'd8780,17'd10238,17'd69692,17'd68930,17'd72567,17'd72568,17'd72669,17'd72670,17'd72159,17'd71879,17'd72671,17'd72571,17'd72572,17'd72361,17'd72162,17'd72672,17'd72673,17'd72674,17'd72675,17'd72676,17'd23291,17'd18137,17'd27431,17'd25488,17'd63639,17'd63640,17'd63789,17'd64630,17'd65286,17'd63378,17'd63808,17'd63808,17'd63808,17'd63808,17'd63808,17'd66073,17'd66073,17'd66073,17'd64651,17'd65054,17'd65054,17'd64651,17'd64651,17'd64651,17'd65054,17'd65054,17'd66319,17'd66318,17'd68519,17'd68519,17'd68944,17'd70061,17'd68833,17'd68520,17'd63807,17'd62850,17'd17179,17'd67427,17'd62976,17'd68634,17'd68634,17'd72677,17'd15102,17'd17543,17'd72678,17'd66791,17'd65553,17'd66180,17'd65552,17'd67420,17'd67662,17'd68288,17'd68408,17'd72581,17'd72366,17'd72679,17'd72367,17'd72367,17'd72367,17'd72680,17'd72583,17'd72681,17'd72682,17'd72683,17'd72478,17'd69147,17'd71076,17'd72684,17'd72685,17'd68187,17'd67673,17'd71901,17'd68738,17'd71416,17'd66076,17'd66320,17'd66320,17'd69800,17'd71191,17'd71191,17'd71191,17'd65055,17'd64789,17'd70059,17'd70164,17'd69797,17'd72686,17'd71420,17'd36903,17'd8187,17'd4882,17'd3423,17'd4712,17'd3898,17'd2249,17'd1240,17'd207,17'd640,17'd72687,17'd206,17'd643,17'd644,17'd803,17'd971,17'd1098,17'd1381,17'd1382,17'd43331,17'd1526,17'd203,17'd42648,17'd205,17'd1410,17'd273,17'd1406
},
'{
17'd6260,17'd4577,17'd4577,17'd6584,17'd4088,17'd3903,17'd4244,17'd4087,17'd4426,17'd4427,17'd4427,17'd4087,17'd4426,17'd4087,17'd5202,17'd4735,17'd5053,17'd5643,17'd72688,17'd72689,17'd72690,17'd72591,17'd72691,17'd72692,17'd72693,17'd71906,17'd66561,17'd71710,17'd69050,17'd6739,17'd70872,17'd9815,17'd4247,17'd63116,17'd72694,17'd64797,17'd64538,17'd12330,17'd6739,17'd64122,17'd63979,17'd6895,17'd8512,17'd72383,17'd9675,17'd66210,17'd9546,17'd72090,17'd6896,17'd7053,17'd13064,17'd71310,17'd6740,17'd6739,17'd66815,17'd67305,17'd66942,17'd70972,17'd63117,17'd1412,17'd11,17'd1128,17'd16,17'd1414,17'd2257,17'd2257,17'd1414,17'd1415,17'd1415,17'd1415,17'd1414,17'd2257,17'd1414,17'd1416,17'd17,17'd18,17'd19,17'd27,17'd27,17'd26,17'd20570,17'd7060,17'd9554,17'd11208,17'd12036,17'd2942,17'd3754,17'd18037,17'd7556,17'd6600,17'd6600,17'd6748,17'd6749,17'd6749,17'd7559,17'd7390,17'd71092,17'd71092,17'd10672,17'd6279,17'd72695,17'd72696,17'd72697,17'd65968,17'd72698,17'd72699,17'd4773,17'd72700,17'd41644,17'd70889,17'd38222,17'd71435,17'd72701,17'd37972,17'd6784,17'd38222,17'd70594,17'd70696,17'd72702,17'd72703,17'd70790,17'd70790,17'd70083,17'd63296,17'd72704,17'd72705,17'd72706,17'd72707,17'd72708,17'd72709,17'd72710,17'd72711,17'd72712,17'd72713,17'd72714,17'd72715,17'd72715,17'd72715,17'd72414,17'd72616,17'd35781,17'd34813,17'd34528,17'd36615,17'd37319,17'd72716,17'd72007,17'd67596,17'd72717,17'd72718,17'd72719,17'd72720,17'd72721,17'd71830,17'd72624,17'd70615,17'd71640,17'd72722,17'd72209,17'd72523,17'd72723,17'd72724,17'd8857,17'd8855,17'd8856,17'd10129,17'd72725,17'd27837,17'd9853,17'd12072,17'd72016,17'd50938,17'd33560,17'd72726,17'd72727,17'd72728,17'd72729,17'd72730,17'd72731,17'd72732,17'd72433,17'd72733,17'd72734,17'd72735,17'd72736,17'd72737,17'd72738,17'd70823,17'd72739,17'd72740,17'd72741,17'd72742,17'd72645,17'd72743,17'd72744,17'd72745,17'd72746,17'd72747,17'd72748,17'd72749,17'd72750,17'd72751,17'd72752,17'd72753,17'd71477,17'd72754,17'd71477,17'd72755,17'd72756,17'd72757,17'd70538,17'd127,17'd70438,17'd1481,17'd130,17'd128,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd132,17'd357,17'd11821,17'd72758,17'd72759,17'd72760,17'd72761,17'd72762,17'd19970,17'd72763,17'd72663,17'd72764,17'd72765,17'd72766,17'd71270,17'd71588,17'd69217,17'd71868,17'd72767,17'd71049,17'd72768,17'd72664,17'd72665,17'd72054,17'd72769,17'd72252,17'd72253,17'd72155,17'd19476,17'd9086,17'd9391,17'd9392,17'd9088,17'd7174,17'd72770,17'd7172,17'd7992,17'd72668,17'd68172,17'd71963,17'd11573,17'd11430,17'd71784,17'd69787,17'd11181,17'd11181,17'd11181,17'd11181,17'd10514,17'd7668,17'd10238,17'd69692,17'd72771,17'd72567,17'd72568,17'd72669,17'd72670,17'd72159,17'd71964,17'd72772,17'd72773,17'd72774,17'd72572,17'd72573,17'd72775,17'd72776,17'd69792,17'd70465,17'd72777,17'd72778,17'd72779,17'd17909,17'd72780,17'd65555,17'd63639,17'd63640,17'd65688,17'd64630,17'd66788,17'd63378,17'd67440,17'd67440,17'd67440,17'd63808,17'd63808,17'd66073,17'd66073,17'd64651,17'd64651,17'd64651,17'd64651,17'd64651,17'd64651,17'd64651,17'd65054,17'd65054,17'd66318,17'd66318,17'd66318,17'd68833,17'd64387,17'd63962,17'd63372,17'd66927,17'd67426,17'd62449,17'd62976,17'd68952,17'd72781,17'd66539,17'd17911,17'd15231,17'd72782,17'd65556,17'd63789,17'd65289,17'd65552,17'd67550,17'd67662,17'd68408,17'd68288,17'd68408,17'd72581,17'd72783,17'd72679,17'd72367,17'd72367,17'd72582,17'd72583,17'd72681,17'd72784,17'd72682,17'd72785,17'd72478,17'd71076,17'd71076,17'd71190,17'd72786,17'd69425,17'd67673,17'd67673,17'd68738,17'd71416,17'd66076,17'd66199,17'd66320,17'd66077,17'd71191,17'd71191,17'd65056,17'd64789,17'd67920,17'd68293,17'd69523,17'd72081,17'd72372,17'd71803,17'd12923,17'd6581,17'd4085,17'd1119,17'd3898,17'd3072,17'd2249,17'd1679,17'd258,17'd640,17'd269,17'd643,17'd643,17'd644,17'd971,17'd1685,17'd1381,17'd202,17'd1382,17'd1526,17'd1382,17'd43059,17'd32250,17'd1687,17'd458,17'd1268,17'd72787
},
'{
17'd4886,17'd7711,17'd4577,17'd27591,17'd6584,17'd4088,17'd4244,17'd3902,17'd4427,17'd4736,17'd69718,17'd9959,17'd5202,17'd5201,17'd5201,17'd5201,17'd5197,17'd5374,17'd72788,17'd72789,17'd72790,17'd71809,17'd65581,17'd65581,17'd64396,17'd72791,17'd72380,17'd72281,17'd65715,17'd72792,17'd72793,17'd66090,17'd1967,17'd1415,17'd64668,17'd72794,17'd72795,17'd72796,17'd12033,17'd66693,17'd70487,17'd7052,17'd7886,17'd7888,17'd8514,17'd8514,17'd7718,17'd68645,17'd68645,17'd6895,17'd6737,17'd64254,17'd71615,17'd13064,17'd68645,17'd12191,17'd65583,17'd66693,17'd63387,17'd1412,17'd21,17'd20,17'd17,17'd17187,17'd4247,17'd4247,17'd1414,17'd1414,17'd1415,17'd1415,17'd1414,17'd1414,17'd1127,17'd15,17'd1127,17'd1414,17'd979,17'd808,17'd980,17'd5516,17'd26,17'd7061,17'd6902,17'd4431,17'd3755,17'd3595,17'd3595,17'd4091,17'd6902,17'd7225,17'd7225,17'd7388,17'd6747,17'd7063,17'd6907,17'd6907,17'd7063,17'd7227,17'd69988,17'd72797,17'd72798,17'd72799,17'd67818,17'd72800,17'd72801,17'd72802,17'd72803,17'd72804,17'd53885,17'd72805,17'd39814,17'd6644,17'd37184,17'd37184,17'd37972,17'd6784,17'd71818,17'd71818,17'd72806,17'd72807,17'd72808,17'd72809,17'd63296,17'd72810,17'd72811,17'd72812,17'd72813,17'd72813,17'd72814,17'd72815,17'd72816,17'd72817,17'd72818,17'd72819,17'd72820,17'd72821,17'd72822,17'd72823,17'd72824,17'd72715,17'd72825,17'd72826,17'd72827,17'd72828,17'd68213,17'd72829,17'd72830,17'd72831,17'd72832,17'd72833,17'd72834,17'd72834,17'd72835,17'd70614,17'd70316,17'd71735,17'd72836,17'd72837,17'd72423,17'd72210,17'd72724,17'd72838,17'd72424,17'd9315,17'd9588,17'd72839,17'd72839,17'd16295,17'd9994,17'd72840,17'd50938,17'd33560,17'd72841,17'd72842,17'd40738,17'd72843,17'd72844,17'd72845,17'd72846,17'd72432,17'd72847,17'd72848,17'd72849,17'd72850,17'd72851,17'd72852,17'd72853,17'd72854,17'd72855,17'd72856,17'd72857,17'd72858,17'd72859,17'd72444,17'd72860,17'd72861,17'd72862,17'd72863,17'd72864,17'd72865,17'd72866,17'd72867,17'd72868,17'd141,17'd141,17'd72655,17'd72869,17'd72870,17'd72871,17'd72872,17'd72873,17'd70537,17'd137,17'd70538,17'd72874,17'd136,17'd130,17'd132,17'd131,17'd131,17'd131,17'd131,17'd132,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd357,17'd70349,17'd72875,17'd72876,17'd72877,17'd72878,17'd72879,17'd72880,17'd72881,17'd72882,17'd72883,17'd72884,17'd69590,17'd68923,17'd72885,17'd69217,17'd71775,17'd72050,17'd71871,17'd72152,17'd72886,17'd72153,17'd72887,17'd72769,17'd72252,17'd72888,17'd72889,17'd9388,17'd9390,17'd10231,17'd10232,17'd9089,17'd7665,17'd7666,17'd7175,17'd8147,17'd72057,17'd7169,17'd11035,17'd11036,17'd11430,17'd71784,17'd69787,17'd32876,17'd32876,17'd11431,17'd11431,17'd10642,17'd9933,17'd9934,17'd31718,17'd68825,17'd72890,17'd72891,17'd72669,17'd72892,17'd72893,17'd72894,17'd72360,17'd72895,17'd72896,17'd72897,17'd72898,17'd71593,17'd72899,17'd72900,17'd69333,17'd72577,17'd72901,17'd72902,17'd17072,17'd72903,17'd64768,17'd65555,17'd63639,17'd63789,17'd65040,17'd64630,17'd66788,17'd68299,17'd67440,17'd67440,17'd67440,17'd65951,17'd69712,17'd69712,17'd64655,17'd69712,17'd67049,17'd66676,17'd66676,17'd66677,17'd66677,17'd68060,17'd68060,17'd72904,17'd66437,17'd64919,17'd65702,17'd65057,17'd64531,17'd65571,17'd67427,17'd62976,17'd68634,17'd68634,17'd14174,17'd66539,17'd18267,17'd14857,17'd66181,17'd72072,17'd63640,17'd66062,17'd71294,17'd72905,17'd67662,17'd68408,17'd68288,17'd68288,17'd72906,17'd72783,17'd72783,17'd72680,17'd72907,17'd72582,17'd72582,17'd72681,17'd72908,17'd72585,17'd72785,17'd72909,17'd69147,17'd71190,17'd71190,17'd72910,17'd69425,17'd69425,17'd69425,17'd69039,17'd67437,17'd67296,17'd67674,17'd66076,17'd66076,17'd67674,17'd66320,17'd65056,17'd67436,17'd67920,17'd70059,17'd71902,17'd71613,17'd70380,17'd65439,17'd58864,17'd8187,17'd4423,17'd445,17'd1263,17'd1962,17'd953,17'd607,17'd41316,17'd261,17'd207,17'd642,17'd970,17'd644,17'd425,17'd972,17'd14315,17'd72911,17'd4731,17'd4731,17'd1382,17'd43059,17'd424,17'd1111,17'd274,17'd72912,17'd1274,17'd72913
},
'{
17'd4886,17'd4886,17'd6583,17'd4577,17'd4887,17'd4245,17'd4428,17'd4244,17'd4427,17'd4736,17'd69718,17'd9959,17'd5202,17'd5201,17'd5201,17'd5201,17'd5197,17'd5374,17'd7540,17'd72914,17'd71987,17'd66684,17'd71809,17'd71809,17'd68848,17'd64795,17'd72915,17'd72792,17'd72916,17'd72916,17'd72487,17'd72917,17'd64400,17'd1414,17'd12929,17'd70972,17'd64798,17'd72918,17'd12033,17'd12033,17'd64537,17'd66815,17'd6896,17'd7220,17'd7888,17'd7716,17'd7718,17'd8344,17'd68645,17'd6896,17'd6895,17'd6739,17'd64397,17'd64254,17'd8043,17'd67815,17'd69249,17'd67305,17'd6433,17'd67453,17'd1128,17'd1128,17'd1277,17'd1415,17'd1127,17'd1689,17'd1414,17'd1414,17'd17,17'd17,17'd1415,17'd1414,17'd1689,17'd1967,17'd1689,17'd1127,17'd1277,17'd979,17'd27,17'd3906,17'd27,17'd286,17'd6902,17'd18037,17'd4091,17'd3595,17'd3595,17'd3755,17'd18037,17'd6902,17'd7728,17'd7728,17'd7557,17'd7063,17'd7063,17'd6907,17'd7390,17'd7227,17'd69988,17'd68646,17'd72919,17'd72920,17'd72921,17'd72922,17'd72923,17'd72924,17'd72925,17'd72926,17'd60788,17'd72927,17'd6487,17'd40274,17'd70697,17'd37593,17'd37972,17'd72928,17'd72929,17'd72929,17'd72928,17'd72928,17'd72930,17'd72931,17'd72932,17'd63296,17'd72933,17'd72812,17'd72813,17'd72813,17'd72707,17'd72934,17'd72934,17'd72935,17'd72936,17'd72937,17'd72938,17'd72939,17'd72940,17'd72941,17'd72942,17'd72943,17'd72944,17'd72945,17'd72946,17'd72947,17'd72419,17'd71923,17'd72948,17'd72948,17'd72949,17'd72950,17'd72951,17'd72951,17'd72952,17'd70614,17'd70812,17'd71832,17'd61988,17'd72423,17'd72210,17'd72628,17'd27329,17'd72838,17'd8855,17'd9020,17'd9589,17'd9993,17'd16045,17'd16296,17'd72953,17'd72954,17'd8553,17'd72955,17'd72956,17'd72957,17'd72958,17'd72959,17'd72960,17'd72961,17'd72962,17'd72963,17'd72848,17'd72964,17'd72965,17'd72966,17'd72967,17'd72968,17'd72969,17'd72439,17'd72970,17'd72971,17'd72744,17'd72972,17'd72973,17'd72974,17'd72974,17'd72975,17'd72976,17'd72977,17'd72978,17'd72979,17'd72980,17'd72981,17'd72982,17'd141,17'd72552,17'd72983,17'd72984,17'd72985,17'd72986,17'd72987,17'd71669,17'd72655,17'd71477,17'd126,17'd72988,17'd141,17'd136,17'd132,17'd131,17'd5593,17'd5593,17'd131,17'd132,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd1481,17'd130,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd2698,17'd72989,17'd72990,17'd72991,17'd72992,17'd72993,17'd22724,17'd21444,17'd72994,17'd72882,17'd72995,17'd72884,17'd69590,17'd68923,17'd72996,17'd69217,17'd71775,17'd72050,17'd71871,17'd72152,17'd72886,17'd71962,17'd72053,17'd72769,17'd72252,17'd16117,17'd72889,17'd9653,17'd11032,17'd10231,17'd10233,17'd9088,17'd7665,17'd7666,17'd7175,17'd8147,17'd72997,17'd7169,17'd70951,17'd68823,17'd11180,17'd11430,17'd69787,17'd32876,17'd32876,17'd11181,17'd11181,17'd10642,17'd27815,17'd9934,17'd31718,17'd68825,17'd72890,17'd72998,17'd72569,17'd72461,17'd72893,17'd72999,17'd72462,17'd71966,17'd73000,17'd72897,17'd72571,17'd73001,17'd73002,17'd72575,17'd73003,17'd73004,17'd73005,17'd73006,17'd17540,17'd13929,17'd25091,17'd64769,17'd65555,17'd63788,17'd63942,17'd65688,17'd64630,17'd64767,17'd65286,17'd66788,17'd66788,17'd71508,17'd63510,17'd65951,17'd69712,17'd69712,17'd64655,17'd63964,17'd66676,17'd65570,17'd66677,17'd66677,17'd66677,17'd66072,17'd66435,17'd65702,17'd65308,17'd64390,17'd17415,17'd62449,17'd62976,17'd68952,17'd72781,17'd14174,17'd66539,17'd18267,17'd17178,17'd15998,17'd63788,17'd65165,17'd67037,17'd65163,17'd68409,17'd67662,17'd68408,17'd73007,17'd73007,17'd73008,17'd72906,17'd72783,17'd72783,17'd72680,17'd72680,17'd72582,17'd72583,17'd72908,17'd72585,17'd72785,17'd72785,17'd72909,17'd69147,17'd71190,17'd71190,17'd73009,17'd73010,17'd69425,17'd69425,17'd67437,17'd67437,17'd67296,17'd67296,17'd66076,17'd66076,17'd67674,17'd66320,17'd64789,17'd71300,17'd67921,17'd68517,17'd70482,17'd71303,17'd73011,17'd59125,17'd9261,17'd6581,17'd4085,17'd1261,17'd1680,17'd1962,17'd1240,17'd1539,17'd261,17'd261,17'd258,17'd271,17'd970,17'd970,17'd425,17'd971,17'd1244,17'd72911,17'd4731,17'd4731,17'd202,17'd1272,17'd605,17'd803,17'd21161,17'd457,17'd1684,17'd73012
},
'{
17'd6419,17'd5196,17'd5196,17'd7711,17'd4887,17'd4733,17'd4088,17'd4428,17'd4244,17'd4244,17'd4736,17'd4427,17'd4087,17'd4087,17'd4087,17'd5202,17'd5645,17'd5197,17'd5374,17'd73013,17'd73014,17'd71807,17'd73015,17'd65579,17'd64537,17'd64253,17'd71989,17'd72380,17'd72281,17'd73016,17'd72281,17'd71615,17'd70874,17'd3750,17'd2781,17'd65314,17'd71908,17'd67575,17'd65583,17'd7886,17'd67305,17'd64120,17'd7547,17'd7053,17'd7886,17'd7718,17'd7888,17'd7888,17'd8191,17'd7052,17'd7053,17'd7221,17'd13576,17'd64397,17'd67574,17'd7886,17'd68645,17'd67574,17'd10922,17'd6267,17'd1830,17'd12,17'd3748,17'd17,17'd14,17'd1127,17'd22965,17'd1416,17'd17,17'd16,17'd1415,17'd1414,17'd1689,17'd1689,17'd1414,17'd1415,17'd289,17'd28,17'd286,17'd980,17'd27,17'd286,17'd6902,17'd18037,17'd5971,17'd3910,17'd5208,17'd5208,17'd5971,17'd6437,17'd7728,17'd8988,17'd7557,17'd6747,17'd6905,17'd7063,17'd73017,17'd7560,17'd7389,17'd6440,17'd12037,17'd73018,17'd73019,17'd73020,17'd73021,17'd73022,17'd73023,17'd73024,17'd60413,17'd73025,17'd73026,17'd41023,17'd6788,17'd51774,17'd6644,17'd72929,17'd73027,17'd73028,17'd70791,17'd6644,17'd73029,17'd72808,17'd72809,17'd63296,17'd72933,17'd73030,17'd63020,17'd73031,17'd73032,17'd73032,17'd73033,17'd62490,17'd73034,17'd73035,17'd73036,17'd73036,17'd73037,17'd72942,17'd72943,17'd73038,17'd73038,17'd73039,17'd72417,17'd72310,17'd71637,17'd70011,17'd73040,17'd69918,17'd71637,17'd73041,17'd73042,17'd71450,17'd70810,17'd71232,17'd73043,17'd72208,17'd73044,17'd73045,17'd71348,17'd26023,17'd72838,17'd72838,17'd8857,17'd9020,17'd9851,17'd9852,17'd9853,17'd11096,17'd73046,17'd73047,17'd53175,17'd73048,17'd73049,17'd73050,17'd73051,17'd73052,17'd73053,17'd73054,17'd73055,17'd73056,17'd73057,17'd72850,17'd73058,17'd72967,17'd73059,17'd72969,17'd73060,17'd73061,17'd73062,17'd73063,17'd73064,17'd73065,17'd72973,17'd72861,17'd73066,17'd73067,17'd73068,17'd73069,17'd73070,17'd73071,17'd73072,17'd73073,17'd141,17'd72982,17'd73074,17'd72986,17'd73075,17'd73076,17'd72986,17'd73077,17'd73078,17'd73079,17'd70537,17'd70537,17'd126,17'd137,17'd136,17'd132,17'd131,17'd131,17'd131,17'd131,17'd132,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd1481,17'd1481,17'd132,17'd132,17'd133,17'd133,17'd130,17'd130,17'd128,17'd5898,17'd73080,17'd72990,17'd72991,17'd73081,17'd73082,17'd54591,17'd20983,17'd73083,17'd73084,17'd72995,17'd73085,17'd68813,17'd68923,17'd73086,17'd69218,17'd71776,17'd73087,17'd71871,17'd72152,17'd73088,17'd72152,17'd71682,17'd73089,17'd72457,17'd16117,17'd15599,17'd9929,17'd11032,17'd10231,17'd10234,17'd9088,17'd9089,17'd7666,17'd7175,17'd8147,17'd72997,17'd7169,17'd6551,17'd68823,17'd11573,17'd11430,17'd11315,17'd70649,17'd70649,17'd11181,17'd11181,17'd10642,17'd27815,17'd9934,17'd31718,17'd68929,17'd73090,17'd73091,17'd73092,17'd72570,17'd72256,17'd72359,17'd71965,17'd72671,17'd73093,17'd73094,17'd72897,17'd73001,17'd73095,17'd73096,17'd73097,17'd73098,17'd73099,17'd73100,17'd72902,17'd22770,17'd23292,17'd24157,17'd64768,17'd65420,17'd63788,17'd63942,17'd70166,17'd65040,17'd71596,17'd64630,17'd65286,17'd65286,17'd63376,17'd63510,17'd63510,17'd63378,17'd63378,17'd63378,17'd63808,17'd63808,17'd66073,17'd66073,17'd66073,17'd63963,17'd63375,17'd65308,17'd64390,17'd73101,17'd69146,17'd14309,17'd67164,17'd72781,17'd73102,17'd66182,17'd17542,17'd65290,17'd72072,17'd64090,17'd66180,17'd66062,17'd71409,17'd71896,17'd72167,17'd67662,17'd68288,17'd68407,17'd73103,17'd72906,17'd72906,17'd73104,17'd73104,17'd72680,17'd72583,17'd73105,17'd72908,17'd72683,17'd72683,17'd72785,17'd72909,17'd69147,17'd69147,17'd71190,17'd71190,17'd68947,17'd73106,17'd67673,17'd67673,17'd67296,17'd67296,17'd71077,17'd67560,17'd71077,17'd67560,17'd65831,17'd65055,17'd65307,17'd67920,17'd68292,17'd69144,17'd72686,17'd65564,17'd66547,17'd58864,17'd8187,17'd4882,17'd3895,17'd1262,17'd1380,17'd953,17'd607,17'd209,17'd262,17'd256,17'd207,17'd271,17'd259,17'd425,17'd205,17'd14066,17'd72911,17'd73107,17'd4731,17'd4731,17'd1244,17'd1244,17'd972,17'd273,17'd189,17'd1274,17'd18387,17'd18387
},
'{
17'd4885,17'd4885,17'd5196,17'd5196,17'd7711,17'd4887,17'd4733,17'd3904,17'd4428,17'd3903,17'd4244,17'd4427,17'd4427,17'd4427,17'd4087,17'd4087,17'd5201,17'd5645,17'd5374,17'd5959,17'd73108,17'd72083,17'd66684,17'd65579,17'd70070,17'd64120,17'd72084,17'd73016,17'd72487,17'd65715,17'd65714,17'd73109,17'd65067,17'd12652,17'd3250,17'd12929,17'd12783,17'd11070,17'd66815,17'd7886,17'd8043,17'd64120,17'd64254,17'd6738,17'd7052,17'd7886,17'd7888,17'd7219,17'd6895,17'd7547,17'd6896,17'd7550,17'd7221,17'd64397,17'd64397,17'd7052,17'd12033,17'd11885,17'd10665,17'd6269,17'd64668,17'd63116,17'd5969,17'd18,17'd0,17'd2,17'd1416,17'd1416,17'd17,17'd16,17'd1415,17'd1414,17'd1127,17'd4247,17'd1415,17'd1415,17'd468,17'd289,17'd287,17'd28,17'd27,17'd6744,17'd73110,17'd10269,17'd6278,17'd5657,17'd5657,17'd5657,17'd5656,17'd6598,17'd9555,17'd9276,17'd7557,17'd7557,17'd73111,17'd6905,17'd69810,17'd7390,17'd7558,17'd73112,17'd5975,17'd73113,17'd73114,17'd73115,17'd73116,17'd73117,17'd73118,17'd73119,17'd73120,17'd73121,17'd73122,17'd73026,17'd40877,17'd51870,17'd73123,17'd73028,17'd73028,17'd52207,17'd60679,17'd73124,17'd73125,17'd73029,17'd73126,17'd72932,17'd73127,17'd73030,17'd72707,17'd72707,17'd73032,17'd73128,17'd61329,17'd73129,17'd73130,17'd73131,17'd73132,17'd73133,17'd73134,17'd73135,17'd73136,17'd72624,17'd73137,17'd72522,17'd72622,17'd72952,17'd73138,17'd73139,17'd73140,17'd73141,17'd73142,17'd73042,17'd71548,17'd73143,17'd73144,17'd73145,17'd59417,17'd73044,17'd73045,17'd73146,17'd27603,17'd27603,17'd8857,17'd8857,17'd8857,17'd9168,17'd9316,17'd73147,17'd73148,17'd72214,17'd73149,17'd54449,17'd48308,17'd73150,17'd73151,17'd73152,17'd73153,17'd73154,17'd40281,17'd73155,17'd73156,17'd73157,17'd73158,17'd73159,17'd73160,17'd73161,17'd73162,17'd73163,17'd73164,17'd73165,17'd73166,17'd73167,17'd73168,17'd73169,17'd73170,17'd73171,17'd73172,17'd73173,17'd73174,17'd73175,17'd73176,17'd73177,17'd70831,17'd72757,17'd71477,17'd72988,17'd73178,17'd72449,17'd73179,17'd73180,17'd73181,17'd73077,17'd73182,17'd73183,17'd73184,17'd70537,17'd126,17'd70438,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd130,17'd128,17'd5898,17'd73080,17'd72875,17'd73185,17'd73186,17'd73187,17'd73188,17'd54407,17'd73189,17'd73190,17'd73191,17'd73192,17'd73193,17'd68923,17'd73194,17'd70149,17'd71775,17'd71049,17'd71962,17'd73195,17'd73088,17'd72152,17'd71778,17'd73196,17'd72457,17'd16117,17'd15600,17'd9387,17'd9389,17'd10231,17'd10234,17'd9088,17'd9089,17'd7666,17'd7175,17'd8146,17'd72997,17'd7169,17'd6385,17'd68823,17'd11573,17'd11430,17'd11315,17'd70649,17'd70649,17'd11181,17'd11181,17'd10642,17'd27815,17'd9934,17'd31718,17'd33993,17'd73197,17'd72567,17'd73198,17'd73199,17'd72358,17'd72256,17'd72257,17'd72360,17'd73093,17'd73094,17'd73094,17'd72898,17'd73001,17'd71055,17'd69790,17'd69138,17'd73200,17'd73201,17'd73006,17'd13684,17'd28421,17'd22598,17'd14580,17'd64768,17'd65420,17'd63788,17'd63942,17'd63942,17'd65040,17'd64507,17'd64767,17'd64630,17'd63247,17'd66789,17'd66078,17'd71975,17'd63247,17'd63247,17'd71975,17'd71975,17'd63108,17'd63108,17'd63375,17'd66078,17'd62852,17'd73202,17'd15734,17'd69146,17'd68952,17'd67173,17'd72781,17'd73102,17'd73203,17'd73204,17'd14975,17'd63640,17'd65165,17'd64368,17'd64902,17'd65163,17'd72076,17'd73205,17'd73206,17'd68288,17'd73008,17'd73207,17'd73208,17'd73209,17'd73209,17'd73104,17'd72680,17'd72583,17'd72584,17'd72908,17'd72585,17'd73210,17'd73210,17'd73211,17'd72478,17'd72478,17'd68837,17'd68837,17'd68947,17'd73212,17'd73212,17'd67673,17'd67673,17'd67674,17'd67674,17'd67560,17'd67560,17'd71077,17'd67560,17'd65055,17'd65307,17'd67920,17'd68292,17'd67923,17'd68518,17'd70380,17'd63652,17'd59125,17'd7705,17'd8186,17'd3391,17'd1261,17'd1263,17'd953,17'd427,17'd41316,17'd41161,17'd262,17'd257,17'd271,17'd259,17'd1112,17'd425,17'd972,17'd971,17'd1381,17'd73107,17'd4731,17'd1382,17'd1244,17'd971,17'd645,17'd409,17'd257,17'd73213,17'd18387,17'd17789
},
'{
17'd2,17'd2,17'd14,17'd1967,17'd1689,17'd3250,17'd4887,17'd4733,17'd4245,17'd4428,17'd4892,17'd4244,17'd3903,17'd3903,17'd4244,17'd4087,17'd5202,17'd5376,17'd5374,17'd5374,17'd73214,17'd73215,17'd63974,17'd68848,17'd64537,17'd70070,17'd64396,17'd65312,17'd65449,17'd67574,17'd71990,17'd67305,17'd64123,17'd71085,17'd6265,17'd1689,17'd73216,17'd69723,17'd64397,17'd65583,17'd8191,17'd67305,17'd63978,17'd6735,17'd6738,17'd7547,17'd7886,17'd7378,17'd6895,17'd6738,17'd7547,17'd7053,17'd8192,17'd6739,17'd71195,17'd13064,17'd6894,17'd6894,17'd69161,17'd13064,17'd65068,17'd64125,17'd3,17'd806,17'd11,17'd3905,17'd1416,17'd1416,17'd809,17'd981,17'd1415,17'd1415,17'd1415,17'd22965,17'd17,17'd17,17'd468,17'd289,17'd18037,17'd18037,17'd4430,17'd6437,17'd6598,17'd11889,17'd12507,17'd13068,17'd13068,17'd13068,17'd13067,17'd5804,17'd11211,17'd9555,17'd7556,17'd7557,17'd73111,17'd70288,17'd69986,17'd73217,17'd6907,17'd11345,17'd12786,17'd13437,17'd73218,17'd73219,17'd73220,17'd73221,17'd73222,17'd73223,17'd73224,17'd54352,17'd73225,17'd73122,17'd73226,17'd73227,17'd73228,17'd60940,17'd60810,17'd52207,17'd73229,17'd73230,17'd73230,17'd73231,17'd73232,17'd73233,17'd73234,17'd73235,17'd72707,17'd72707,17'd73031,17'd73128,17'd61987,17'd61987,17'd73236,17'd61595,17'd73237,17'd73132,17'd73135,17'd73238,17'd73239,17'd71639,17'd73240,17'd72952,17'd72835,17'd73041,17'd73241,17'd73242,17'd73242,17'd73243,17'd73244,17'd73245,17'd73246,17'd73247,17'd73248,17'd72114,17'd73249,17'd73250,17'd73251,17'd33393,17'd13222,17'd13222,17'd9168,17'd9168,17'd9168,17'd9316,17'd73147,17'd73148,17'd72214,17'd72525,17'd73252,17'd73253,17'd73254,17'd73255,17'd73256,17'd73257,17'd73258,17'd73259,17'd73260,17'd73261,17'd73262,17'd73263,17'd73264,17'd73265,17'd73266,17'd73267,17'd73268,17'd73269,17'd73270,17'd73271,17'd73272,17'd73273,17'd73274,17'd73275,17'd73276,17'd73277,17'd73278,17'd73279,17'd73280,17'd73281,17'd73282,17'd72866,17'd72983,17'd73283,17'd73284,17'd73285,17'd73286,17'd73287,17'd73288,17'd73289,17'd73290,17'd73291,17'd73292,17'd73072,17'd73293,17'd70742,17'd70437,17'd127,17'd130,17'd130,17'd130,17'd130,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd131,17'd133,17'd133,17'd132,17'd132,17'd720,17'd2698,17'd15202,17'd73294,17'd73185,17'd73295,17'd73296,17'd73297,17'd20517,17'd73298,17'd73299,17'd73300,17'd73301,17'd73193,17'd70048,17'd73194,17'd70149,17'd71776,17'd73302,17'd71962,17'd73195,17'd73088,17'd72886,17'd72052,17'd73089,17'd72457,17'd16950,17'd72888,17'd14044,17'd9519,17'd10378,17'd10234,17'd9088,17'd9089,17'd7666,17'd7175,17'd8146,17'd72997,17'd7167,17'd6385,17'd68823,17'd11573,17'd11430,17'd11315,17'd70649,17'd70649,17'd11181,17'd27932,17'd10642,17'd27815,17'd10380,17'd31718,17'd33993,17'd69410,17'd73303,17'd73304,17'd73305,17'd73199,17'd72256,17'd72257,17'd73306,17'd73307,17'd73308,17'd73309,17'd73310,17'd73001,17'd71055,17'd73311,17'd73312,17'd73313,17'd15994,17'd73314,17'd26954,17'd23291,17'd28421,17'd22598,17'd14580,17'd64768,17'd63495,17'd65420,17'd63640,17'd65553,17'd66306,17'd72268,17'd64630,17'd63247,17'd63247,17'd63247,17'd73315,17'd73315,17'd66790,17'd66790,17'd66790,17'd62973,17'd62973,17'd62852,17'd73316,17'd73202,17'd16255,17'd68634,17'd13808,17'd13418,17'd72781,17'd65690,17'd73203,17'd64905,17'd64631,17'd63639,17'd64227,17'd68057,17'd65163,17'd67787,17'd67549,17'd73206,17'd73317,17'd73103,17'd73103,17'd73208,17'd73208,17'd73208,17'd73318,17'd73318,17'd73104,17'd73319,17'd73320,17'd72908,17'd72683,17'd73211,17'd73321,17'd73321,17'd73322,17'd73323,17'd72172,17'd68837,17'd68947,17'd68947,17'd73212,17'd73212,17'd71901,17'd67673,17'd67674,17'd71077,17'd67560,17'd73324,17'd67560,17'd66075,17'd64653,17'd64241,17'd64529,17'd66804,17'd68519,17'd72271,17'd70380,17'd65439,17'd38460,17'd8186,17'd4729,17'd229,17'd625,17'd626,17'd427,17'd209,17'd408,17'd408,17'd262,17'd257,17'd271,17'd271,17'd643,17'd425,17'd204,17'd1244,17'd72911,17'd73107,17'd1245,17'd1381,17'd14315,17'd972,17'd1963,17'd21161,17'd1964,17'd1404,17'd17789,17'd73325
},
'{
17'd0,17'd0,17'd15,17'd14,17'd1967,17'd1689,17'd7711,17'd4887,17'd4245,17'd6420,17'd4428,17'd4428,17'd3903,17'd3903,17'd4244,17'd4087,17'd5202,17'd5377,17'd5960,17'd5374,17'd7540,17'd72914,17'd71306,17'd63975,17'd64396,17'd65449,17'd64537,17'd63816,17'd64396,17'd11885,17'd71906,17'd65583,17'd73326,17'd64123,17'd70874,17'd2781,17'd73327,17'd13065,17'd63978,17'd65449,17'd68645,17'd12033,17'd63978,17'd13184,17'd6592,17'd6894,17'd8191,17'd8191,17'd7547,17'd7221,17'd7547,17'd7547,17'd7549,17'd8343,17'd13815,17'd71310,17'd6735,17'd6593,17'd11885,17'd67574,17'd64256,17'd70076,17'd1,17'd806,17'd11,17'd1128,17'd3905,17'd1416,17'd30,17'd809,17'd1415,17'd17187,17'd17,17'd1416,17'd1416,17'd17,17'd468,17'd809,17'd3907,17'd9554,17'd5971,17'd5803,17'd12931,17'd5808,17'd5383,17'd12787,17'd13437,17'd12787,17'd32729,17'd5808,17'd6110,17'd11211,17'd6904,17'd7557,17'd8047,17'd73111,17'd73328,17'd73217,17'd9277,17'd69438,17'd6109,17'd5382,17'd66694,17'd72284,17'd73329,17'd73330,17'd73331,17'd73332,17'd73333,17'd73334,17'd63706,17'd61590,17'd62889,17'd73335,17'd73336,17'd73228,17'd73123,17'd52207,17'd6948,17'd73337,17'd73338,17'd73230,17'd73231,17'd73339,17'd73340,17'd73341,17'd72813,17'd73342,17'd73342,17'd73250,17'd73343,17'd73343,17'd73343,17'd73343,17'd73344,17'd73345,17'd73346,17'd73347,17'd73348,17'd73144,17'd71450,17'd73349,17'd73142,17'd73142,17'd73350,17'd73351,17'd73352,17'd73353,17'd73354,17'd73355,17'd73356,17'd73357,17'd72422,17'd72315,17'd73358,17'd73359,17'd33393,17'd7105,17'd8224,17'd8224,17'd9168,17'd9448,17'd9316,17'd73360,17'd73361,17'd73362,17'd72525,17'd50599,17'd49115,17'd46711,17'd73363,17'd73364,17'd73365,17'd73366,17'd73367,17'd73368,17'd73369,17'd73370,17'd73371,17'd73372,17'd73373,17'd73374,17'd73375,17'd73376,17'd73269,17'd73377,17'd73378,17'd73379,17'd72546,17'd73380,17'd72648,17'd73381,17'd73382,17'd73383,17'd73384,17'd73385,17'd73386,17'd72240,17'd73387,17'd72986,17'd73183,17'd73284,17'd73388,17'd73389,17'd73390,17'd73391,17'd73392,17'd73393,17'd73394,17'd73395,17'd73396,17'd73397,17'd72869,17'd70742,17'd70437,17'd127,17'd130,17'd130,17'd130,17'd130,17'd136,17'd136,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd131,17'd131,17'd131,17'd133,17'd132,17'd132,17'd720,17'd135,17'd17139,17'd73398,17'd73399,17'd73400,17'd73401,17'd56526,17'd73402,17'd22075,17'd73403,17'd73404,17'd73405,17'd73193,17'd70048,17'd69322,17'd69323,17'd69683,17'd71049,17'd71962,17'd73195,17'd73088,17'd72886,17'd72153,17'd73406,17'd72457,17'd16950,17'd72888,17'd9386,17'd9388,17'd9390,17'd10233,17'd9088,17'd9089,17'd7666,17'd7666,17'd8146,17'd72997,17'd7167,17'd6386,17'd68823,17'd11573,17'd11430,17'd11315,17'd69787,17'd69787,17'd27932,17'd27932,17'd10515,17'd10515,17'd27815,17'd69692,17'd33993,17'd69410,17'd73407,17'd73408,17'd73409,17'd73305,17'd73410,17'd72359,17'd73411,17'd73412,17'd73308,17'd73413,17'd73414,17'd73415,17'd73416,17'd70953,17'd73417,17'd73418,17'd73419,17'd65680,17'd73420,17'd26954,17'd13805,17'd23291,17'd22598,17'd24157,17'd25091,17'd63495,17'd63639,17'd63640,17'd65553,17'd66306,17'd64507,17'd64630,17'd64630,17'd64630,17'd64630,17'd65688,17'd65040,17'd66536,17'd66536,17'd65816,17'd65816,17'd65816,17'd15231,17'd17659,17'd14174,17'd13808,17'd73421,17'd65422,17'd73422,17'd73423,17'd64370,17'd65554,17'd64227,17'd68057,17'd64902,17'd65163,17'd73424,17'd73425,17'd68288,17'd73103,17'd73208,17'd73208,17'd73103,17'd73208,17'd73208,17'd73208,17'd73318,17'd73426,17'd73319,17'd73320,17'd72908,17'd72683,17'd73211,17'd73211,17'd73321,17'd73321,17'd73322,17'd73323,17'd72172,17'd72172,17'd68947,17'd68947,17'd73212,17'd73212,17'd71901,17'd71901,17'd67674,17'd71077,17'd73324,17'd73324,17'd66075,17'd64921,17'd65306,17'd64529,17'd66804,17'd66928,17'd72271,17'd73427,17'd66547,17'd64648,17'd8507,17'd5194,17'd3895,17'd1401,17'd626,17'd627,17'd1539,17'd1242,17'd408,17'd40563,17'd262,17'd256,17'd258,17'd426,17'd606,17'd425,17'd204,17'd1272,17'd1381,17'd73107,17'd1381,17'd1244,17'd1685,17'd644,17'd10073,17'd268,17'd596,17'd1404,17'd27824,17'd73325
},
'{
17'd12,17'd12,17'd0,17'd0,17'd14,17'd1689,17'd3250,17'd2422,17'd4246,17'd14743,17'd6420,17'd6420,17'd4088,17'd4088,17'd3903,17'd4087,17'd5202,17'd5202,17'd5376,17'd5197,17'd5374,17'd70486,17'd73428,17'd71307,17'd64253,17'd64120,17'd65449,17'd64396,17'd64253,17'd70070,17'd12191,17'd12191,17'd12330,17'd12500,17'd63820,17'd13186,17'd6096,17'd10801,17'd65067,17'd71195,17'd67305,17'd12033,17'd63979,17'd63980,17'd67306,17'd6736,17'd68645,17'd8043,17'd73429,17'd12329,17'd7721,17'd10921,17'd6737,17'd8343,17'd6593,17'd63980,17'd63821,17'd6735,17'd11885,17'd65583,17'd67574,17'd63980,17'd73430,17'd806,17'd11,17'd1128,17'd3905,17'd1416,17'd30,17'd30,17'd1415,17'd17187,17'd17,17'd3905,17'd4089,17'd17,17'd29,17'd809,17'd3255,17'd11210,17'd11889,17'd5809,17'd5383,17'd32562,17'd53229,17'd30197,17'd69541,17'd69541,17'd53229,17'd32562,17'd5659,17'd12337,17'd10408,17'd9970,17'd7557,17'd73111,17'd73328,17'd69986,17'd7560,17'd7731,17'd11890,17'd13579,17'd73431,17'd73432,17'd73115,17'd64802,17'd73433,17'd73434,17'd73435,17'd73436,17'd73437,17'd73438,17'd73439,17'd61455,17'd73440,17'd70987,17'd73441,17'd60810,17'd6948,17'd40122,17'd73442,17'd73443,17'd73444,17'd73445,17'd73446,17'd73447,17'd73448,17'd73449,17'd73449,17'd73450,17'd73451,17'd73451,17'd73452,17'd61860,17'd73344,17'd73453,17'd73454,17'd73455,17'd73456,17'd73457,17'd73458,17'd73459,17'd73349,17'd73460,17'd73351,17'd73461,17'd73352,17'd73462,17'd73463,17'd73464,17'd73465,17'd60813,17'd57797,17'd73466,17'd73467,17'd26023,17'd33393,17'd8224,17'd12823,17'd7266,17'd9170,17'd9316,17'd9591,17'd73361,17'd73468,17'd73469,17'd50599,17'd49115,17'd36927,17'd73470,17'd41180,17'd73471,17'd73472,17'd73473,17'd73474,17'd73475,17'd73476,17'd73477,17'd73478,17'd73479,17'd73480,17'd73481,17'd73376,17'd73482,17'd73483,17'd73484,17'd73485,17'd73486,17'd73487,17'd73488,17'd73489,17'd73382,17'd73490,17'd73491,17'd73492,17'd73493,17'd73494,17'd73495,17'd73496,17'd73497,17'd73498,17'd73388,17'd73499,17'd73500,17'd73501,17'd73502,17'd73503,17'd73504,17'd73505,17'd73506,17'd73290,17'd73389,17'd73507,17'd70831,17'd72658,17'd70438,17'd130,17'd130,17'd130,17'd136,17'd136,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd131,17'd131,17'd133,17'd133,17'd132,17'd132,17'd356,17'd134,17'd17139,17'd73508,17'd73509,17'd73510,17'd73511,17'd59106,17'd73512,17'd73513,17'd73514,17'd73515,17'd73516,17'd73517,17'd70048,17'd73194,17'd70149,17'd71273,17'd71870,17'd71962,17'd73195,17'd73088,17'd73195,17'd72153,17'd73406,17'd72457,17'd73518,17'd73519,17'd15220,17'd9653,17'd11033,17'd10232,17'd9392,17'd9521,17'd7666,17'd7666,17'd6848,17'd72997,17'd7167,17'd6386,17'd11035,17'd11573,17'd11430,17'd11315,17'd69787,17'd69787,17'd27932,17'd27932,17'd27932,17'd10515,17'd10515,17'd10515,17'd68510,17'd69325,17'd73090,17'd73303,17'd73520,17'd73521,17'd73199,17'd72256,17'd73522,17'd73523,17'd73524,17'd73525,17'd73414,17'd72773,17'd73526,17'd71391,17'd70055,17'd73527,17'd68732,17'd66909,17'd15995,17'd73420,17'd27085,17'd73528,17'd23291,17'd22598,17'd18748,17'd17177,17'd64509,17'd65288,17'd65042,17'd72072,17'd63789,17'd65040,17'd66306,17'd66306,17'd65040,17'd65040,17'd65556,17'd65556,17'd65689,17'd66915,17'd15231,17'd15231,17'd18267,17'd14174,17'd66183,17'd65422,17'd65422,17'd13054,17'd73529,17'd65043,17'd65041,17'd67037,17'd64902,17'd65163,17'd65037,17'd73530,17'd73531,17'd73007,17'd68407,17'd73532,17'd73532,17'd73533,17'd73208,17'd73208,17'd73318,17'd73318,17'd73534,17'd73534,17'd73535,17'd73536,17'd72683,17'd73321,17'd73321,17'd73322,17'd73322,17'd73322,17'd73322,17'd73322,17'd72478,17'd72172,17'd73212,17'd73212,17'd73212,17'd73212,17'd71982,17'd71901,17'd71415,17'd71416,17'd73324,17'd73324,17'd73537,17'd63657,17'd63965,17'd65703,17'd70259,17'd68519,17'd70270,17'd66547,17'd59125,17'd7705,17'd6095,17'd3425,17'd1119,17'd446,17'd623,17'd428,17'd1097,17'd595,17'd2255,17'd595,17'd262,17'd256,17'd640,17'd3746,17'd205,17'd1537,17'd204,17'd1272,17'd202,17'd202,17'd1244,17'd1244,17'd971,17'd803,17'd935,17'd2115,17'd69346,17'd26728,17'd20009,17'd17789
},
'{
17'd12,17'd12,17'd1,17'd1,17'd15,17'd1127,17'd1688,17'd2422,17'd4887,17'd14743,17'd6420,17'd6420,17'd4088,17'd3904,17'd3903,17'd3902,17'd4087,17'd5202,17'd5377,17'd5645,17'd5509,17'd5374,17'd73538,17'd73539,17'd64253,17'd63976,17'd65449,17'd67305,17'd64795,17'd64253,17'd68645,17'd12191,17'd12330,17'd70387,17'd13576,17'd71196,17'd6260,17'd73540,17'd73541,17'd63980,17'd65449,17'd67574,17'd6735,17'd63820,17'd71714,17'd6431,17'd11885,17'd68645,17'd12501,17'd12034,17'd10921,17'd7051,17'd6735,17'd6592,17'd6897,17'd13184,17'd65189,17'd13815,17'd11885,17'd67816,17'd12191,17'd13815,17'd13434,17'd73542,17'd2423,17'd1128,17'd18,17'd1416,17'd290,17'd290,17'd1415,17'd1277,17'd18,17'd18,17'd4089,17'd4089,17'd288,17'd654,17'd2941,17'd73543,17'd12786,17'd5384,17'd4899,17'd30197,17'd6116,17'd5815,17'd5815,17'd5815,17'd4901,17'd30197,17'd32087,17'd5659,17'd11345,17'd10409,17'd9970,17'd7557,17'd71521,17'd6905,17'd7227,17'd7391,17'd7562,17'd12200,17'd73544,17'd13306,17'd73545,17'd73546,17'd73547,17'd73548,17'd73549,17'd73550,17'd73551,17'd73552,17'd73553,17'd73554,17'd73555,17'd73440,17'd70987,17'd73123,17'd51869,17'd38603,17'd51775,17'd73556,17'd73557,17'd73558,17'd73559,17'd73560,17'd73561,17'd73562,17'd73563,17'd73450,17'd73564,17'd73564,17'd73452,17'd60324,17'd73565,17'd73565,17'd73566,17'd73567,17'd73568,17'd73569,17'd73570,17'd73243,17'd73244,17'd73352,17'd73571,17'd73571,17'd73350,17'd73572,17'd73356,17'd73573,17'd72422,17'd72208,17'd73358,17'd73251,17'd25397,17'd33393,17'd13222,17'd13222,17'd7266,17'd9170,17'd9317,17'd9591,17'd14641,17'd30206,17'd73469,17'd73574,17'd53175,17'd7274,17'd73575,17'd73576,17'd73577,17'd73578,17'd73579,17'd73580,17'd73581,17'd73582,17'd73583,17'd73584,17'd73585,17'd73586,17'd73587,17'd73588,17'd73589,17'd73590,17'd73591,17'd73592,17'd73593,17'd73488,17'd73488,17'd73594,17'd73489,17'd73595,17'd72862,17'd73596,17'd73597,17'd73598,17'd73599,17'd73600,17'd73601,17'd73602,17'd73603,17'd73604,17'd73605,17'd73501,17'd73606,17'd73607,17'd73608,17'd73609,17'd73610,17'd73505,17'd73076,17'd73290,17'd73611,17'd73612,17'd70538,17'd1481,17'd132,17'd132,17'd130,17'd136,17'd136,17'd130,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd131,17'd131,17'd131,17'd133,17'd132,17'd132,17'd1481,17'd1759,17'd15202,17'd73613,17'd19427,17'd73614,17'd28300,17'd57585,17'd20366,17'd53659,17'd73615,17'd73616,17'd73617,17'd73517,17'd70048,17'd69322,17'd69323,17'd71273,17'd71870,17'd71962,17'd73195,17'd73088,17'd73195,17'd72355,17'd73406,17'd72563,17'd73518,17'd73519,17'd15220,17'd9929,17'd14162,17'd10232,17'd9392,17'd9521,17'd7666,17'd7666,17'd6848,17'd72997,17'd7167,17'd6550,17'd11035,17'd11573,17'd11430,17'd11315,17'd69787,17'd69787,17'd27932,17'd27932,17'd27932,17'd27932,17'd10642,17'd10642,17'd68510,17'd69325,17'd73090,17'd73407,17'd73618,17'd73619,17'd73305,17'd73410,17'd72257,17'd73620,17'd73621,17'd73525,17'd73622,17'd73623,17'd73624,17'd73625,17'd73626,17'd73627,17'd73628,17'd73629,17'd73630,17'd64763,17'd73631,17'd73006,17'd73528,17'd23291,17'd17072,17'd18029,17'd18266,17'd14432,17'd64508,17'd65287,17'd63788,17'd63788,17'd63789,17'd65553,17'd63789,17'd63788,17'd15482,17'd15482,17'd65290,17'd17414,17'd17414,17'd17542,17'd73632,17'd73422,17'd13289,17'd13289,17'd13054,17'd18030,17'd73633,17'd15230,17'd63940,17'd64628,17'd65163,17'd73424,17'd73530,17'd73634,17'd73007,17'd73635,17'd73636,17'd73637,17'd73638,17'd73533,17'd73639,17'd73208,17'd73640,17'd73318,17'd73534,17'd73641,17'd73320,17'd73642,17'd73643,17'd73321,17'd73322,17'd73322,17'd73322,17'd73322,17'd73322,17'd73322,17'd72909,17'd72785,17'd72477,17'd72172,17'd73212,17'd73212,17'd71982,17'd71901,17'd71415,17'd71416,17'd73324,17'd73324,17'd67800,17'd63657,17'd65570,17'd66677,17'd70259,17'd70662,17'd73011,17'd70272,17'd58864,17'd8187,17'd3896,17'd3246,17'd625,17'd626,17'd782,17'd3100,17'd2255,17'd2255,17'd2255,17'd595,17'd262,17'd256,17'd640,17'd2779,17'd205,17'd1537,17'd424,17'd1272,17'd202,17'd202,17'd1244,17'd971,17'd645,17'd10073,17'd967,17'd69615,17'd69346,17'd965,17'd20009,17'd73644
},
'{
17'd18,17'd19,17'd1,17'd0,17'd15,17'd15,17'd1689,17'd2422,17'd2784,17'd2935,17'd4245,17'd6420,17'd4088,17'd3904,17'd3903,17'd3902,17'd4087,17'd4087,17'd9959,17'd5202,17'd5197,17'd6263,17'd7212,17'd71614,17'd64663,17'd63976,17'd70070,17'd66815,17'd65712,17'd63975,17'd65712,17'd8191,17'd8043,17'd7547,17'd12033,17'd64397,17'd70777,17'd6096,17'd73645,17'd73646,17'd71310,17'd65449,17'd13064,17'd63979,17'd63822,17'd9550,17'd6894,17'd67305,17'd12329,17'd73429,17'd64399,17'd6590,17'd10922,17'd66942,17'd7051,17'd70587,17'd63980,17'd66447,17'd67574,17'd67574,17'd65449,17'd6740,17'd10088,17'd73647,17'd3,17'd2423,17'd18,17'd16,17'd809,17'd30,17'd17,17'd16,17'd19,17'd18,17'd20404,17'd4089,17'd289,17'd809,17'd3754,17'd5210,17'd5383,17'd6284,17'd5063,17'd26128,17'd73648,17'd73649,17'd26976,17'd25651,17'd11893,17'd29446,17'd6115,17'd32087,17'd12337,17'd11345,17'd10409,17'd69724,17'd9276,17'd8048,17'd70288,17'd6905,17'd9277,17'd70880,17'd73650,17'd73651,17'd73652,17'd73653,17'd73654,17'd73655,17'd73656,17'd73657,17'd73658,17'd73659,17'd73660,17'd73661,17'd73662,17'd73663,17'd73664,17'd71105,17'd73665,17'd73665,17'd73666,17'd73667,17'd73668,17'd73669,17'd73670,17'd73671,17'd73672,17'd73561,17'd73673,17'd73563,17'd73674,17'd73674,17'd73675,17'd73676,17'd73677,17'd73678,17'd73679,17'd57667,17'd73680,17'd73681,17'd73682,17'd73683,17'd73684,17'd73684,17'd73352,17'd73244,17'd73570,17'd73685,17'd73464,17'd73043,17'd72722,17'd73686,17'd73687,17'd26023,17'd7105,17'd8224,17'd12823,17'd29457,17'd9170,17'd9852,17'd13614,17'd11632,17'd73688,17'd28803,17'd32115,17'd33395,17'd48308,17'd73689,17'd40431,17'd73690,17'd73691,17'd73692,17'd73693,17'd73694,17'd73695,17'd73696,17'd73697,17'd73698,17'd73699,17'd73700,17'd73701,17'd73702,17'd73377,17'd73703,17'd73592,17'd73704,17'd73705,17'd73706,17'd73706,17'd73383,17'd73707,17'd73708,17'd73709,17'd73710,17'd73711,17'd73712,17'd73713,17'd73714,17'd73715,17'd73716,17'd73717,17'd73609,17'd73718,17'd73719,17'd73720,17'd73607,17'd72449,17'd73721,17'd73180,17'd73722,17'd73723,17'd73724,17'd73497,17'd70831,17'd70538,17'd1481,17'd132,17'd132,17'd130,17'd130,17'd130,17'd132,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd131,17'd131,17'd133,17'd133,17'd132,17'd132,17'd4163,17'd130,17'd2861,17'd73725,17'd73726,17'd73727,17'd73728,17'd73729,17'd20670,17'd73730,17'd73731,17'd73732,17'd73733,17'd73734,17'd70360,17'd69403,17'd70149,17'd71273,17'd71870,17'd72152,17'd73088,17'd73088,17'd73195,17'd72355,17'd73735,17'd72457,17'd73736,17'd73736,17'd15471,17'd9929,17'd9389,17'd10775,17'd9087,17'd9521,17'd7666,17'd7175,17'd8146,17'd8147,17'd7167,17'd7168,17'd11035,17'd68823,17'd68927,17'd69691,17'd70649,17'd70649,17'd27932,17'd10897,17'd27932,17'd27932,17'd27815,17'd10515,17'd28183,17'd29158,17'd73197,17'd73197,17'd73737,17'd73303,17'd73198,17'd73738,17'd71878,17'd73739,17'd72895,17'd73623,17'd73622,17'd73740,17'd73624,17'd73741,17'd71391,17'd73742,17'd69232,17'd73743,17'd73744,17'd14053,17'd73745,17'd73746,17'd73747,17'd73748,17'd17412,17'd13416,17'd20553,17'd18506,17'd18138,17'd73633,17'd15733,17'd65042,17'd72072,17'd15482,17'd15482,17'd15482,17'd65290,17'd73749,17'd73749,17'd73749,17'd14173,17'd13686,17'd73750,17'd73750,17'd13417,17'd73751,17'd18030,17'd17177,17'd73752,17'd73753,17'd66914,17'd65683,17'd67420,17'd67419,17'd67548,17'd68832,17'd68179,17'd73754,17'd73755,17'd73754,17'd73756,17'd73756,17'd73639,17'd73318,17'd73426,17'd73757,17'd73641,17'd73758,17'd73759,17'd73760,17'd73761,17'd73762,17'd73763,17'd73322,17'd73763,17'd73322,17'd73321,17'd73764,17'd72785,17'd72477,17'd72477,17'd72476,17'd73212,17'd73212,17'd72276,17'd72276,17'd71981,17'd71703,17'd68739,17'd66074,17'd69531,17'd65306,17'd64529,17'd68060,17'd69708,17'd73765,17'd65439,17'd59125,17'd64525,17'd4883,17'd3099,17'd228,17'd2249,17'd627,17'd429,17'd1094,17'd211,17'd2420,17'd2255,17'd255,17'd802,17'd974,17'd7539,17'd644,17'd972,17'd972,17'd424,17'd1272,17'd1244,17'd1244,17'd971,17'd971,17'd274,17'd21161,17'd49713,17'd69536,17'd1683,17'd181,17'd805,17'd181
},
'{
17'd18,17'd18,17'd1,17'd0,17'd15,17'd15,17'd1967,17'd1688,17'd2422,17'd2784,17'd4733,17'd4245,17'd4088,17'd3904,17'd9960,17'd4244,17'd4244,17'd4427,17'd4427,17'd5202,17'd5645,17'd6263,17'd5377,17'd71706,17'd73766,17'd64253,17'd64396,17'd65449,17'd12191,17'd68848,17'd63975,17'd8043,17'd7052,17'd7547,17'd67815,17'd65583,17'd65067,17'd13186,17'd73327,17'd73767,17'd12928,17'd64397,17'd13576,17'd63979,17'd63822,17'd13816,17'd6740,17'd6739,17'd72796,17'd73429,17'd11735,17'd11607,17'd6270,17'd10922,17'd6590,17'd10665,17'd63980,17'd66447,17'd71195,17'd13576,17'd64254,17'd63979,17'd9550,17'd73768,17'd4884,17'd3,17'd1277,17'd1277,17'd809,17'd30,17'd17,17'd16,17'd19,17'd18,17'd20404,17'd3905,17'd289,17'd809,17'd3754,17'd5658,17'd4899,17'd5063,17'd26128,17'd11741,17'd25116,17'd25116,17'd7232,17'd7232,17'd73649,17'd11893,17'd31415,17'd73769,17'd5659,17'd12337,17'd11345,17'd10409,17'd9685,17'd70686,17'd7729,17'd7729,17'd7390,17'd71092,17'd73770,17'd66336,17'd54787,17'd73771,17'd73772,17'd73773,17'd73548,17'd73774,17'd73775,17'd73776,17'd73777,17'd73778,17'd73779,17'd73780,17'd73781,17'd43752,17'd60678,17'd73782,17'd60938,17'd60938,17'd73667,17'd73783,17'd73784,17'd73785,17'd73786,17'd73672,17'd73787,17'd73788,17'd73789,17'd73790,17'd73790,17'd73675,17'd73676,17'd73677,17'd73679,17'd73679,17'd57667,17'd57933,17'd58908,17'd73791,17'd73792,17'd73684,17'd73793,17'd73570,17'd73570,17'd73794,17'd72013,17'd59417,17'd62124,17'd73795,17'd26023,17'd33393,17'd8224,17'd7267,17'd7764,17'd12824,17'd9852,17'd9319,17'd11632,17'd29458,17'd29051,17'd8083,17'd48936,17'd7274,17'd73796,17'd73797,17'd73798,17'd73799,17'd73800,17'd73801,17'd73802,17'd73803,17'd73804,17'd73805,17'd73806,17'd73807,17'd73808,17'd73809,17'd73810,17'd73811,17'd73812,17'd73813,17'd73814,17'd73815,17'd73816,17'd73817,17'd73818,17'd73819,17'd73820,17'd73821,17'd73822,17'd73823,17'd73824,17'd73825,17'd73826,17'd73827,17'd73828,17'd73602,17'd73827,17'd73829,17'd73830,17'd73831,17'd73832,17'd73393,17'd73394,17'd73833,17'd73834,17'd73835,17'd73834,17'd73836,17'd73497,17'd73388,17'd72754,17'd133,17'd131,17'd131,17'd132,17'd130,17'd130,17'd132,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd131,17'd131,17'd131,17'd133,17'd132,17'd132,17'd356,17'd132,17'd15202,17'd73837,17'd73838,17'd73839,17'd73840,17'd73841,17'd60385,17'd22726,17'd73842,17'd73843,17'd73844,17'd73845,17'd70048,17'd73846,17'd73847,17'd71273,17'd71870,17'd71962,17'd73195,17'd73088,17'd73195,17'd72153,17'd73735,17'd72457,17'd73736,17'd73736,17'd15471,17'd9387,17'd9519,17'd10511,17'd9087,17'd9392,17'd73848,17'd7666,17'd6848,17'd8147,17'd7167,17'd6550,17'd11035,17'd68621,17'd68927,17'd69691,17'd69787,17'd70649,17'd27932,17'd10897,17'd27932,17'd27932,17'd10515,17'd10515,17'd28183,17'd28057,17'd69325,17'd73197,17'd73197,17'd73737,17'd73408,17'd73198,17'd73849,17'd73850,17'd72258,17'd73740,17'd73623,17'd73740,17'd73851,17'd73852,17'd73853,17'd71170,17'd69516,17'd69136,17'd73743,17'd73744,17'd66530,17'd73854,17'd73855,17'd73856,17'd12767,17'd17540,17'd12478,17'd64092,17'd13288,17'd73857,17'd18138,17'd14432,17'd64508,17'd64508,17'd64508,17'd65043,17'd65043,17'd73529,17'd18030,17'd18030,17'd17910,17'd13417,17'd73858,17'd73859,17'd63641,17'd13685,17'd14580,17'd73860,17'd73861,17'd73862,17'd65551,17'd73863,17'd67419,17'd73864,17'd68832,17'd68179,17'd73865,17'd73865,17'd73636,17'd73754,17'd73756,17'd73866,17'd73867,17'd73318,17'd73757,17'd73868,17'd73869,17'd73759,17'd73870,17'd73761,17'd73762,17'd73762,17'd73322,17'd73322,17'd73322,17'd73321,17'd73321,17'd73643,17'd72683,17'd72585,17'd73871,17'd73871,17'd72477,17'd73212,17'd71801,17'd71801,17'd71981,17'd71609,17'd68839,17'd69243,17'd69531,17'd65703,17'd67423,17'd66318,17'd69338,17'd66801,17'd59125,17'd58865,17'd5789,17'd3423,17'd228,17'd446,17'd627,17'd609,17'd20008,17'd1095,17'd2420,17'd2420,17'd2115,17'd2115,17'd974,17'd262,17'd269,17'd644,17'd1687,17'd972,17'd424,17'd1272,17'd1244,17'd971,17'd972,17'd803,17'd73872,17'd2588,17'd1403,17'd69153,17'd1683,17'd253,17'd461,17'd461
},
'{
17'd0,17'd0,17'd1,17'd0,17'd15,17'd1830,17'd15,17'd1689,17'd3250,17'd3250,17'd2784,17'd2935,17'd4245,17'd4245,17'd3904,17'd4088,17'd4428,17'd4244,17'd4427,17'd4427,17'd5201,17'd4734,17'd5645,17'd7212,17'd71614,17'd64663,17'd64253,17'd64537,17'd68645,17'd65713,17'd63975,17'd70070,17'd73873,17'd72090,17'd71713,17'd71713,17'd64254,17'd71196,17'd70277,17'd73874,17'd71908,17'd65313,17'd64399,17'd64399,17'd65313,17'd63668,17'd70178,17'd66942,17'd67305,17'd13064,17'd7376,17'd6433,17'd9419,17'd7376,17'd11205,17'd70587,17'd11205,17'd11070,17'd65188,17'd12928,17'd63979,17'd12928,17'd67306,17'd10264,17'd63669,17'd1412,17'd14442,17'd9422,17'd1415,17'd1414,17'd17,17'd1416,17'd18,17'd18,17'd18,17'd3905,17'd289,17'd809,17'd3754,17'd13950,17'd53229,17'd6116,17'd11741,17'd25651,17'd25116,17'd73875,17'd9283,17'd7232,17'd7395,17'd27826,17'd28320,17'd26236,17'd26733,17'd5809,17'd11737,17'd70077,17'd9555,17'd8197,17'd70288,17'd7729,17'd69986,17'd8989,17'd7228,17'd73770,17'd73876,17'd64540,17'd73877,17'd73878,17'd73879,17'd73880,17'd73881,17'd73882,17'd73883,17'd73884,17'd73885,17'd73886,17'd5862,17'd6016,17'd43604,17'd61456,17'd61456,17'd73887,17'd73888,17'd73667,17'd51870,17'd73443,17'd73889,17'd73786,17'd73890,17'd73561,17'd73787,17'd73789,17'd73789,17'd73790,17'd73891,17'd73891,17'd73892,17'd73892,17'd73892,17'd57412,17'd60558,17'd73893,17'd73894,17'd73895,17'd73896,17'd73455,17'd73455,17'd73897,17'd72315,17'd73466,17'd73146,17'd27603,17'd7105,17'd7267,17'd9021,17'd13613,17'd9171,17'd9591,17'd9319,17'd14641,17'd73898,17'd73899,17'd50850,17'd52634,17'd73900,17'd73796,17'd73901,17'd73902,17'd73903,17'd73904,17'd73905,17'd73906,17'd73907,17'd73908,17'd73909,17'd73910,17'd73911,17'd73912,17'd73913,17'd73914,17'd73915,17'd73916,17'd73917,17'd73918,17'd73919,17'd73920,17'd73921,17'd73922,17'd73923,17'd73924,17'd73924,17'd73925,17'd73492,17'd73926,17'd73927,17'd73928,17'd73723,17'd73929,17'd73930,17'd73931,17'd73932,17'd73933,17'd73934,17'd73935,17'd73936,17'd73937,17'd73506,17'd73394,17'd73938,17'd73834,17'd73075,17'd73939,17'd73072,17'd72655,17'd20762,17'd128,17'd132,17'd131,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd1481,17'd132,17'd131,17'd131,17'd131,17'd133,17'd132,17'd132,17'd356,17'd128,17'd2861,17'd73940,17'd73941,17'd73942,17'd73943,17'd73944,17'd27810,17'd73945,17'd73946,17'd73947,17'd73948,17'd73949,17'd73950,17'd73846,17'd73951,17'd73952,17'd71870,17'd71962,17'd72355,17'd73088,17'd73195,17'd71778,17'd73953,17'd72563,17'd73736,17'd73519,17'd15471,17'd14044,17'd10895,17'd10230,17'd9392,17'd9392,17'd10234,17'd10235,17'd6848,17'd8147,17'd7169,17'd6550,17'd10512,17'd68621,17'd73954,17'd69128,17'd69787,17'd69787,17'd69787,17'd71784,17'd10897,17'd27932,17'd10641,17'd10641,17'd10515,17'd28183,17'd29158,17'd34792,17'd69325,17'd73197,17'd69326,17'd72567,17'd73955,17'd73956,17'd73739,17'd72063,17'd73093,17'd72895,17'd73851,17'd73957,17'd73958,17'd71278,17'd70154,17'd73959,17'd73960,17'd73961,17'd73962,17'd14577,17'd73963,17'd73964,17'd73965,17'd12630,17'd73966,17'd12171,17'd12768,17'd73967,17'd18751,17'd27087,17'd18752,17'd18507,17'd73968,17'd73969,17'd73969,17'd65044,17'd13173,17'd13173,17'd73970,17'd73970,17'd73971,17'd73972,17'd72903,17'd24157,17'd70855,17'd69977,17'd73862,17'd73973,17'd66913,17'd67160,17'd67786,17'd67915,17'd73974,17'd73975,17'd73865,17'd73865,17'd73754,17'd73754,17'd73976,17'd73866,17'd73318,17'd73426,17'd73977,17'd73978,17'd73979,17'd73980,17'd73981,17'd73761,17'd73762,17'd73762,17'd73321,17'd73321,17'd73764,17'd73321,17'd73982,17'd73983,17'd72683,17'd73642,17'd73984,17'd73984,17'd72370,17'd72276,17'd71981,17'd71703,17'd73985,17'd71514,17'd69887,17'd69531,17'd64109,17'd65570,17'd66928,17'd69145,17'd73427,17'd73986,17'd58865,17'd6094,17'd3897,17'd5195,17'd1402,17'd2587,17'd1122,17'd622,17'd2420,17'd182,17'd181,17'd182,17'd1123,17'd73987,17'd974,17'd268,17'd272,17'd643,17'd1124,17'd1687,17'd971,17'd1685,17'd971,17'd972,17'd1828,17'd273,17'd18390,17'd254,17'd69536,17'd69154,17'd1683,17'd461,17'd254,17'd460
},
'{
17'd0,17'd1,17'd1,17'd0,17'd1830,17'd1830,17'd15,17'd14,17'd1689,17'd2781,17'd3250,17'd2935,17'd4245,17'd4245,17'd3904,17'd3904,17'd4428,17'd4892,17'd4244,17'd4427,17'd4087,17'd4735,17'd5197,17'd5645,17'd71706,17'd73988,17'd63976,17'd65449,17'd65713,17'd67816,17'd65713,17'd64795,17'd73109,17'd72090,17'd8344,17'd71713,17'd11885,17'd65067,17'd70680,17'd73989,17'd63387,17'd63668,17'd11205,17'd64124,17'd70178,17'd63668,17'd71908,17'd6594,17'd13064,17'd13815,17'd7376,17'd6733,17'd6268,17'd9270,17'd9270,17'd11735,17'd6590,17'd11607,17'd71197,17'd13185,17'd13816,17'd63980,17'd13433,17'd63821,17'd73990,17'd63117,17'd14442,17'd14442,17'd1415,17'd1415,17'd17,17'd22965,17'd3905,17'd18,17'd19,17'd16,17'd289,17'd809,17'd3755,17'd13950,17'd53229,17'd5815,17'd73648,17'd73649,17'd25116,17'd73991,17'd73875,17'd7232,17'd9282,17'd6605,17'd28320,17'd26236,17'd73992,17'd34004,17'd6110,17'd70077,17'd9555,17'd8047,17'd70288,17'd7729,17'd69987,17'd7559,17'd6906,17'd7731,17'd73993,17'd73994,17'd73995,17'd73996,17'd73997,17'd73998,17'd73999,17'd74000,17'd74001,17'd74002,17'd74003,17'd73885,17'd54712,17'd62744,17'd74004,17'd74005,17'd74006,17'd73664,17'd60808,17'd74007,17'd74008,17'd51870,17'd73443,17'd74009,17'd73785,17'd73559,17'd74010,17'd74011,17'd74011,17'd74012,17'd74012,17'd73790,17'd73790,17'd73790,17'd73790,17'd73891,17'd73892,17'd60558,17'd73893,17'd59038,17'd74013,17'd74014,17'd74015,17'd57666,17'd73466,17'd73251,17'd33393,17'd12372,17'd7267,17'd8388,17'd7926,17'd14490,17'd9172,17'd14641,17'd74016,17'd74017,17'd31932,17'd74018,17'd52555,17'd7113,17'd73796,17'd73901,17'd74019,17'd74020,17'd74021,17'd74022,17'd74023,17'd74024,17'd74025,17'd74026,17'd74027,17'd74028,17'd74029,17'd74030,17'd74031,17'd74032,17'd74033,17'd74034,17'd74035,17'd74036,17'd74037,17'd74038,17'd74039,17'd74040,17'd74041,17'd74042,17'd74043,17'd74044,17'd74045,17'd74046,17'd74047,17'd74048,17'd74049,17'd74050,17'd74051,17'd74052,17'd74053,17'd74054,17'd73606,17'd73393,17'd74055,17'd73506,17'd74056,17'd74057,17'd73938,17'd73834,17'd73836,17'd73507,17'd73388,17'd72552,17'd136,17'd134,17'd132,17'd131,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd1481,17'd130,17'd132,17'd131,17'd131,17'd133,17'd132,17'd132,17'd356,17'd128,17'd2861,17'd74058,17'd74059,17'd73942,17'd73943,17'd74060,17'd27810,17'd74061,17'd22384,17'd74062,17'd74063,17'd74064,17'd74065,17'd73846,17'd74066,17'd74067,17'd71870,17'd72052,17'd72153,17'd73088,17'd73195,17'd72251,17'd73953,17'd72769,17'd73736,17'd74068,17'd15471,17'd15220,17'd9388,17'd11032,17'd9087,17'd9392,17'd10234,17'd10235,17'd6848,17'd8147,17'd7167,17'd7168,17'd6850,17'd68621,17'd73954,17'd69128,17'd69787,17'd69787,17'd69787,17'd69787,17'd10897,17'd27932,17'd11576,17'd10641,17'd10515,17'd10515,17'd28183,17'd34792,17'd69325,17'd74069,17'd69129,17'd74070,17'd74071,17'd72569,17'd73850,17'd74072,17'd72063,17'd72063,17'd72360,17'd74073,17'd74074,17'd71501,17'd71390,17'd70253,17'd74075,17'd74076,17'd74077,17'd67154,17'd14577,17'd74078,17'd74079,17'd74080,17'd74081,17'd74082,17'd74083,17'd74084,17'd62426,17'd62561,17'd74085,17'd74085,17'd12910,17'd63232,17'd63232,17'd74086,17'd74087,17'd74088,17'd74089,17'd74090,17'd13929,17'd26331,17'd74091,17'd69794,17'd65162,17'd66786,17'd66786,17'd66786,17'd67418,17'd74092,17'd67785,17'd74093,17'd73975,17'd73975,17'd74094,17'd73865,17'd74095,17'd73756,17'd73866,17'd74096,17'd73534,17'd73868,17'd74097,17'd74098,17'd74099,17'd73981,17'd73761,17'd73761,17'd73762,17'd73762,17'd73762,17'd73321,17'd73321,17'd73643,17'd73983,17'd74100,17'd73642,17'd72908,17'd74101,17'd73984,17'd72171,17'd72276,17'd71981,17'd73985,17'd71514,17'd69887,17'd69241,17'd66321,17'd65570,17'd66437,17'd70061,17'd69339,17'd66802,17'd74102,17'd6890,17'd4883,17'd4712,17'd3072,17'd2587,17'd234,17'd622,17'd611,17'd182,17'd639,17'd182,17'd1683,17'd1403,17'd73987,17'd262,17'd271,17'd644,17'd643,17'd1124,17'd1828,17'd971,17'd972,17'd972,17'd644,17'd273,17'd189,17'd188,17'd1123,17'd1548,17'd74103,17'd1826,17'd461,17'd254,17'd460
},
'{
17'd1,17'd1412,17'd1,17'd1,17'd1,17'd1,17'd0,17'd14,17'd1127,17'd1689,17'd3250,17'd2422,17'd3101,17'd3101,17'd2593,17'd2782,17'd6420,17'd4892,17'd4892,17'd4244,17'd4427,17'd4087,17'd4735,17'd4734,17'd69718,17'd71421,17'd63817,17'd71195,17'd64120,17'd67305,17'd12191,17'd63976,17'd74104,17'd74105,17'd70976,17'd74106,17'd68645,17'd13815,17'd74107,17'd73989,17'd10668,17'd69255,17'd64667,17'd70178,17'd70178,17'd65313,17'd14441,17'd63520,17'd14186,17'd14186,17'd10799,17'd7714,17'd6269,17'd64667,17'd64799,17'd6268,17'd7885,17'd9683,17'd6273,17'd69255,17'd67817,17'd71714,17'd63978,17'd13433,17'd6268,17'd14867,17'd14742,17'd15,17'd17187,17'd16,17'd18,17'd26344,17'd3905,17'd18,17'd1277,17'd16,17'd289,17'd289,17'd4431,17'd12336,17'd74108,17'd29446,17'd29447,17'd28433,17'd25116,17'd25116,17'd25116,17'd26976,17'd74109,17'd74110,17'd5063,17'd73769,17'd5221,17'd5808,17'd6110,17'd11211,17'd6903,17'd8047,17'd70288,17'd73111,17'd6748,17'd6905,17'd7559,17'd7560,17'd7562,17'd74111,17'd74112,17'd74113,17'd74114,17'd74115,17'd74116,17'd74117,17'd74118,17'd74119,17'd4935,17'd73884,17'd74120,17'd54811,17'd74121,17'd73780,17'd73555,17'd74005,17'd6326,17'd52711,17'd74122,17'd74123,17'd74124,17'd74125,17'd74126,17'd73785,17'd74127,17'd74128,17'd74129,17'd74011,17'd74130,17'd74012,17'd74012,17'd74012,17'd74131,17'd74131,17'd74132,17'd74133,17'd74134,17'd57412,17'd73678,17'd74135,17'd74136,17'd74137,17'd74138,17'd74139,17'd74139,17'd9021,17'd74140,17'd7926,17'd74141,17'd74016,17'd74142,17'd74143,17'd74144,17'd74145,17'd74146,17'd54272,17'd7435,17'd74147,17'd74148,17'd74149,17'd74150,17'd74151,17'd74152,17'd74153,17'd74154,17'd74155,17'd74156,17'd74157,17'd74158,17'd74159,17'd74160,17'd74161,17'd74162,17'd74163,17'd74164,17'd74165,17'd74166,17'd74167,17'd74168,17'd74169,17'd74169,17'd74170,17'd74171,17'd74172,17'd74173,17'd74174,17'd74175,17'd74176,17'd74177,17'd74178,17'd74179,17'd73075,17'd74180,17'd74181,17'd74182,17'd74183,17'd74184,17'd74055,17'd74185,17'd73833,17'd74186,17'd74187,17'd73834,17'd72985,17'd74188,17'd72983,17'd74189,17'd20762,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd1481,17'd130,17'd132,17'd132,17'd131,17'd133,17'd132,17'd132,17'd4163,17'd128,17'd3168,17'd6691,17'd74190,17'd74191,17'd74192,17'd74193,17'd74194,17'd56410,17'd62306,17'd74195,17'd74196,17'd74197,17'd74198,17'd73846,17'd74066,17'd74199,17'd71870,17'd72052,17'd74200,17'd73088,17'd73088,17'd72251,17'd73735,17'd73196,17'd73736,17'd74068,17'd15334,17'd10773,17'd9929,17'd9389,17'd9783,17'd74201,17'd10234,17'd10235,17'd6848,17'd8146,17'd7167,17'd7169,17'd6217,17'd10512,17'd68621,17'd11573,17'd11315,17'd69787,17'd32719,17'd32719,17'd10897,17'd27932,17'd11576,17'd10641,17'd27815,17'd27815,17'd27933,17'd28057,17'd68622,17'd74202,17'd74069,17'd73090,17'd73303,17'd73198,17'd72670,17'd73850,17'd74203,17'd74072,17'd74072,17'd74073,17'd74204,17'd74205,17'd71500,17'd70154,17'd73959,17'd74075,17'd68284,17'd74206,17'd14169,17'd74207,17'd31554,17'd24316,17'd74208,17'd74209,17'd74210,17'd63948,17'd62313,17'd23293,17'd22772,17'd74211,17'd74212,17'd74213,17'd74214,17'd74215,17'd74216,17'd74217,17'd74218,17'd27816,17'd71795,17'd70661,17'd65284,17'd74219,17'd66785,17'd66785,17'd67283,17'd67033,17'd67785,17'd68054,17'd73975,17'd73975,17'd74220,17'd74220,17'd74095,17'd74095,17'd73756,17'd73756,17'd73866,17'd74221,17'd73868,17'd74097,17'd73979,17'd73980,17'd74222,17'd74223,17'd74224,17'd74225,17'd73762,17'd73762,17'd73761,17'd73761,17'd73643,17'd73760,17'd74100,17'd74226,17'd72784,17'd72584,17'd74101,17'd74227,17'd72080,17'd72080,17'd74228,17'd71799,17'd70376,17'd68290,17'd67422,17'd63964,17'd66072,17'd68945,17'd69421,17'd66802,17'd74229,17'd10395,17'd14060,17'd5357,17'd3072,17'd3248,17'd447,17'd793,17'd611,17'd964,17'd592,17'd213,17'd180,17'd1548,17'd1404,17'd2255,17'd268,17'd271,17'd643,17'd643,17'd1687,17'd1551,17'd1828,17'd1124,17'd643,17'd644,17'd273,17'd267,17'd456,17'd18387,17'd15492,17'd401,17'd1826,17'd461,17'd254,17'd2255
},
'{
17'd1412,17'd1412,17'd1412,17'd1,17'd1,17'd1,17'd1,17'd2,17'd1127,17'd1127,17'd1688,17'd2422,17'd2935,17'd3101,17'd2593,17'd2782,17'd4245,17'd6420,17'd4892,17'd4892,17'd3903,17'd4427,17'd5201,17'd4735,17'd5202,17'd71304,17'd65838,17'd63977,17'd64120,17'd70070,17'd67816,17'd67816,17'd74230,17'd65714,17'd74231,17'd74231,17'd8043,17'd7547,17'd12928,17'd71312,17'd63116,17'd68083,17'd9552,17'd64667,17'd64666,17'd70178,17'd63520,17'd9552,17'd74232,17'd8822,17'd67306,17'd10799,17'd70587,17'd64667,17'd6433,17'd6268,17'd9419,17'd10662,17'd6589,17'd74233,17'd74234,17'd71714,17'd71708,17'd66693,17'd6269,17'd6273,17'd63259,17'd63116,17'd16,17'd1277,17'd18,17'd4089,17'd4089,17'd16,17'd1277,17'd16,17'd289,17'd289,17'd4431,17'd5804,17'd5059,17'd26014,17'd5666,17'd4902,17'd4099,17'd4264,17'd73649,17'd27826,17'd74110,17'd26472,17'd74235,17'd11611,17'd5659,17'd12507,17'd6110,17'd11211,17'd6903,17'd7728,17'd7557,17'd7557,17'd6747,17'd7063,17'd7063,17'd8198,17'd71521,17'd10408,17'd74236,17'd74237,17'd74238,17'd74114,17'd74239,17'd74240,17'd74241,17'd74242,17'd74243,17'd74244,17'd74245,17'd60907,17'd74246,17'd63018,17'd73780,17'd74004,17'd43351,17'd48644,17'd42936,17'd6648,17'd59809,17'd59414,17'd74247,17'd74248,17'd74249,17'd74250,17'd74251,17'd74252,17'd74129,17'd74130,17'd74130,17'd73787,17'd74253,17'd74131,17'd74131,17'd74131,17'd74254,17'd74131,17'd74255,17'd74256,17'd74257,17'd74139,17'd74139,17'd9021,17'd9021,17'd13613,17'd7926,17'd7594,17'd74258,17'd31428,17'd31932,17'd74259,17'd74018,17'd74260,17'd53531,17'd74261,17'd74262,17'd74263,17'd74264,17'd74265,17'd74266,17'd74267,17'd74268,17'd74269,17'd74270,17'd74271,17'd74272,17'd74273,17'd74274,17'd74275,17'd74276,17'd74277,17'd74278,17'd74279,17'd74165,17'd74280,17'd74281,17'd74282,17'd74283,17'd74284,17'd74284,17'd74285,17'd74286,17'd74287,17'd74288,17'd74289,17'd74290,17'd74291,17'd74292,17'd74293,17'd74294,17'd73500,17'd74295,17'd74296,17'd74054,17'd73606,17'd73179,17'd72866,17'd73604,17'd73389,17'd74187,17'd74297,17'd74298,17'd72984,17'd74299,17'd74300,17'd1481,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd1481,17'd130,17'd132,17'd132,17'd131,17'd133,17'd132,17'd132,17'd356,17'd128,17'd3168,17'd6691,17'd74301,17'd74302,17'd74192,17'd74303,17'd74304,17'd59107,17'd57862,17'd74305,17'd74306,17'd74307,17'd74308,17'd74309,17'd74066,17'd74310,17'd74311,17'd72052,17'd74200,17'd73195,17'd73088,17'd71778,17'd74312,17'd73196,17'd73518,17'd74313,17'd15334,17'd10773,17'd9929,17'd10895,17'd13029,17'd74314,17'd10235,17'd7010,17'd7175,17'd8146,17'd7167,17'd7991,17'd6850,17'd10379,17'd73954,17'd69691,17'd69787,17'd69787,17'd32876,17'd32876,17'd10897,17'd27932,17'd10641,17'd10641,17'd10515,17'd27815,17'd27933,17'd28183,17'd68510,17'd68622,17'd69325,17'd74069,17'd73090,17'd73303,17'd74315,17'd73849,17'd74316,17'd73522,17'd73739,17'd74072,17'd74317,17'd74318,17'd71688,17'd71390,17'd70253,17'd69231,17'd68938,17'd74319,17'd74320,17'd74321,17'd31719,17'd29029,17'd23119,17'd32877,17'd74322,17'd74323,17'd63948,17'd62185,17'd62185,17'd74324,17'd74325,17'd74325,17'd74326,17'd74327,17'd62052,17'd74328,17'd15345,17'd65161,17'd74329,17'd66178,17'd66532,17'd66784,17'd69140,17'd74330,17'd74331,17'd74332,17'd68406,17'd68406,17'd68406,17'd68406,17'd73975,17'd74220,17'd74095,17'd74095,17'd73756,17'd74333,17'd74221,17'd74334,17'd73869,17'd74335,17'd73980,17'd74099,17'd74223,17'd74223,17'd74225,17'd74225,17'd73762,17'd73761,17'd73761,17'd73981,17'd73760,17'd74336,17'd74226,17'd73536,17'd72681,17'd72681,17'd74101,17'd74337,17'd72079,17'd74338,17'd71899,17'd74339,17'd67919,17'd67421,17'd66788,17'd63964,17'd66317,17'd69421,17'd66925,17'd74102,17'd10395,17'd6891,17'd37708,17'd4400,17'd1402,17'd2587,17'd234,17'd633,17'd212,17'd592,17'd213,17'd250,17'd17422,17'd17185,17'd73644,17'd801,17'd646,17'd260,17'd1538,17'd643,17'd14597,17'd1551,17'd1124,17'd1829,17'd206,17'd272,17'd935,17'd264,17'd965,17'd18271,17'd15492,17'd17422,17'd1826,17'd17551,17'd595,17'd2115
},
'{
17'd3,17'd283,17'd3,17'd3,17'd3,17'd283,17'd3,17'd12,17'd2,17'd1127,17'd1688,17'd1688,17'd2422,17'd3252,17'd2935,17'd2784,17'd4246,17'd4245,17'd4428,17'd4428,17'd3903,17'd3903,17'd4087,17'd4426,17'd5201,17'd9959,17'd74340,17'd65187,17'd64396,17'd64537,17'd65581,17'd12191,17'd74341,17'd74341,17'd72175,17'd74105,17'd68645,17'd8043,17'd13576,17'd69723,17'd63117,17'd62981,17'd14867,17'd63668,17'd64798,17'd64666,17'd9683,17'd6273,17'd74342,17'd6734,17'd13815,17'd63979,17'd10799,17'd10403,17'd10662,17'd10662,17'd6103,17'd6103,17'd6589,17'd73990,17'd74343,17'd73541,17'd71708,17'd71195,17'd63821,17'd8823,17'd63521,17'd63118,17'd1277,17'd19,17'd20404,17'd3905,17'd13,17'd2,17'd16,17'd17187,17'd29,17'd289,17'd4248,17'd5804,17'd32562,17'd69541,17'd30198,17'd5666,17'd73648,17'd73649,17'd27826,17'd29447,17'd26128,17'd74344,17'd4900,17'd69622,17'd12786,17'd6109,17'd11889,17'd6598,17'd6902,17'd9275,17'd7556,17'd9276,17'd7227,17'd7227,17'd69724,17'd8048,17'd70388,17'd7557,17'd11345,17'd74345,17'd72284,17'd74346,17'd74347,17'd74348,17'd74349,17'd74350,17'd74351,17'd74352,17'd74353,17'd74354,17'd63156,17'd60936,17'd74355,17'd54100,17'd74356,17'd74357,17'd43073,17'd43206,17'd44522,17'd41925,17'd40879,17'd74358,17'd74359,17'd74360,17'd74249,17'd74361,17'd74362,17'd74129,17'd74130,17'd74130,17'd74363,17'd74363,17'd74253,17'd74364,17'd74364,17'd73562,17'd74365,17'd10702,17'd9021,17'd9021,17'd9021,17'd7764,17'd7593,17'd7926,17'd11240,17'd30357,17'd31428,17'd31932,17'd74366,17'd74260,17'd54272,17'd52633,17'd74367,17'd74368,17'd74369,17'd74370,17'd74371,17'd74372,17'd74373,17'd74374,17'd74375,17'd74376,17'd74377,17'd74378,17'd74273,17'd74379,17'd74380,17'd74381,17'd74382,17'd74383,17'd74279,17'd74384,17'd74385,17'd74386,17'd74387,17'd74388,17'd74389,17'd74390,17'd74391,17'd74392,17'd74393,17'd74394,17'd74395,17'd74396,17'd74397,17'd74398,17'd74399,17'd74400,17'd74400,17'd74400,17'd74401,17'd74402,17'd74403,17'd73713,17'd74298,17'd74404,17'd73290,17'd72551,17'd74405,17'd74406,17'd74056,17'd74407,17'd72242,17'd71154,17'd133,17'd11541,17'd131,17'd132,17'd132,17'd130,17'd132,17'd132,17'd132,17'd132,17'd1481,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd1481,17'd1481,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd1481,17'd356,17'd2698,17'd2865,17'd74408,17'd74409,17'd74410,17'd74411,17'd74412,17'd20513,17'd74413,17'd74414,17'd74415,17'd74416,17'd74417,17'd74418,17'd74419,17'd74420,17'd74421,17'd72052,17'd74200,17'd73195,17'd74422,17'd74423,17'd73196,17'd73196,17'd73518,17'd74313,17'd15334,17'd10773,17'd9387,17'd9388,17'd9655,17'd9783,17'd10235,17'd7010,17'd7175,17'd6848,17'd7167,17'd7825,17'd6216,17'd6850,17'd68621,17'd68927,17'd11430,17'd69787,17'd32719,17'd32876,17'd10897,17'd27932,17'd10641,17'd10641,17'd27932,17'd27932,17'd27933,17'd27933,17'd27933,17'd28183,17'd28057,17'd34792,17'd69410,17'd74424,17'd74425,17'd74426,17'd73199,17'd72256,17'd72257,17'd71879,17'd71879,17'd74318,17'd74427,17'd74428,17'd70154,17'd69329,17'd69032,17'd74076,17'd74429,17'd15097,17'd12474,17'd29029,17'd23467,17'd74430,17'd5489,17'd63499,17'd74431,17'd4547,17'd32244,17'd74432,17'd74433,17'd74432,17'd74434,17'd74435,17'd19594,17'd74436,17'd74437,17'd74438,17'd70854,17'd74439,17'd74440,17'd74441,17'd74442,17'd74442,17'd74443,17'd74444,17'd68178,17'd68178,17'd74445,17'd74445,17'd74446,17'd74446,17'd74095,17'd74095,17'd73756,17'd74333,17'd74447,17'd74448,17'd74335,17'd74449,17'd74450,17'd74223,17'd74225,17'd74225,17'd74225,17'd74225,17'd73761,17'd73643,17'd73643,17'd73760,17'd74451,17'd74226,17'd73320,17'd73535,17'd72681,17'd72784,17'd74337,17'd74452,17'd74453,17'd74454,17'd74339,17'd74455,17'd70771,17'd66788,17'd65951,17'd67049,17'd69238,17'd69339,17'd66802,17'd58864,17'd14312,17'd4575,17'd4712,17'd1825,17'd447,17'd234,17'd244,17'd212,17'd40102,17'd251,17'd1543,17'd589,17'd17552,17'd17422,17'd27824,17'd967,17'd646,17'd207,17'd206,17'd643,17'd1411,17'd74456,17'd1273,17'd72687,17'd206,17'd272,17'd268,17'd1274,17'd17789,17'd17422,17'd17552,17'd15492,17'd639,17'd253,17'd460,17'd2115
},
'{
17'd3,17'd3,17'd3,17'd3,17'd3,17'd283,17'd283,17'd3,17'd0,17'd466,17'd4247,17'd1689,17'd3250,17'd2422,17'd2935,17'd2784,17'd4887,17'd4733,17'd4088,17'd4428,17'd3903,17'd3903,17'd4427,17'd4426,17'd4426,17'd9959,17'd71304,17'd74457,17'd63977,17'd64120,17'd65449,17'd66815,17'd74105,17'd74458,17'd65447,17'd74459,17'd11885,17'd12191,17'd11885,17'd67306,17'd74460,17'd14742,17'd64125,17'd64930,17'd11070,17'd70178,17'd6268,17'd10662,17'd74234,17'd73646,17'd10799,17'd63821,17'd13816,17'd9132,17'd8194,17'd6101,17'd10662,17'd8669,17'd6589,17'd6589,17'd74343,17'd70873,17'd64122,17'd64929,17'd63820,17'd10401,17'd10662,17'd64125,17'd3749,17'd16,17'd3905,17'd19,17'd2,17'd2,17'd16,17'd16,17'd29,17'd29,17'd653,17'd3910,17'd5807,17'd4898,17'd53229,17'd12508,17'd69541,17'd6116,17'd6116,17'd5665,17'd6115,17'd74461,17'd69622,17'd12656,17'd67454,17'd11889,17'd10269,17'd6598,17'd6902,17'd6902,17'd9555,17'd9685,17'd69724,17'd69724,17'd70686,17'd8197,17'd74462,17'd70388,17'd7390,17'd6280,17'd51861,17'd74463,17'd74464,17'd74465,17'd74466,17'd74467,17'd74468,17'd74469,17'd74470,17'd74471,17'd74472,17'd63156,17'd74473,17'd74355,17'd62744,17'd54101,17'd74474,17'd74475,17'd6160,17'd42938,17'd51104,17'd54030,17'd58175,17'd74476,17'd74477,17'd74249,17'd74478,17'd74479,17'd74480,17'd74480,17'd74481,17'd31749,17'd31749,17'd31426,17'd31426,17'd31273,17'd74482,17'd34025,17'd13613,17'd13613,17'd13613,17'd7926,17'd13614,17'd12221,17'd74483,17'd30206,17'd31932,17'd74259,17'd74146,17'd54272,17'd52633,17'd74261,17'd74484,17'd74485,17'd74486,17'd74487,17'd74488,17'd74489,17'd74490,17'd74491,17'd74492,17'd74493,17'd74494,17'd74495,17'd74496,17'd74497,17'd74498,17'd74499,17'd73271,17'd72336,17'd74500,17'd74166,17'd74501,17'd74502,17'd74503,17'd74504,17'd74390,17'd74505,17'd74506,17'd74507,17'd74508,17'd74509,17'd74510,17'd74511,17'd74512,17'd74513,17'd74514,17'd74515,17'd74516,17'd74517,17'd74518,17'd74519,17'd73393,17'd73289,17'd73610,17'd74520,17'd73286,17'd74521,17'd74522,17'd74523,17'd74188,17'd73388,17'd72552,17'd356,17'd11541,17'd131,17'd131,17'd132,17'd132,17'd130,17'd132,17'd132,17'd132,17'd132,17'd1481,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd1481,17'd130,17'd132,17'd132,17'd131,17'd133,17'd132,17'd133,17'd1481,17'd356,17'd2698,17'd13534,17'd74524,17'd74525,17'd74526,17'd74527,17'd74528,17'd20673,17'd21125,17'd74529,17'd74530,17'd74531,17'd74532,17'd14556,17'd74533,17'd74534,17'd74535,17'd72052,17'd72052,17'd73195,17'd74536,17'd74537,17'd72769,17'd73196,17'd16733,17'd74313,17'd15334,17'd10773,17'd9387,17'd9388,17'd9085,17'd9656,17'd11848,17'd7010,17'd10235,17'd7175,17'd7169,17'd7825,17'd6216,17'd7176,17'd10379,17'd68927,17'd11430,17'd71784,17'd69787,17'd32719,17'd27932,17'd10897,17'd10897,17'd10641,17'd27932,17'd27932,17'd27932,17'd27933,17'd27933,17'd28183,17'd28057,17'd27934,17'd69325,17'd73090,17'd74538,17'd73520,17'd74539,17'd74540,17'd72358,17'd72159,17'd73850,17'd72892,17'd74541,17'd74542,17'd71499,17'd69971,17'd74543,17'd74075,17'd74544,17'd74545,17'd16739,17'd31892,17'd24155,17'd11860,17'd10519,17'd74546,17'd74547,17'd74548,17'd74209,17'd19355,17'd74549,17'd74550,17'd21315,17'd74551,17'd74552,17'd74553,17'd74554,17'd70466,17'd74555,17'd74556,17'd74557,17'd74558,17'd74559,17'd74560,17'd74560,17'd74444,17'd74561,17'd74561,17'd74445,17'd74446,17'd74446,17'd74095,17'd74095,17'd73756,17'd73866,17'd74221,17'd74334,17'd74562,17'd74449,17'd74563,17'd74223,17'd74223,17'd74450,17'd74225,17'd74225,17'd74564,17'd73762,17'd73643,17'd73760,17'd74336,17'd74565,17'd74097,17'd73535,17'd73535,17'd72784,17'd74101,17'd74337,17'd74566,17'd74567,17'd74568,17'd67791,17'd65164,17'd66663,17'd67440,17'd67049,17'd64919,17'd69339,17'd66925,17'd74229,17'd64525,17'd6582,17'd5357,17'd1824,17'd1264,17'd1122,17'd799,17'd611,17'd636,17'd249,17'd433,17'd589,17'd400,17'd74569,17'd15354,17'd460,17'd263,17'd207,17'd426,17'd206,17'd643,17'd270,17'd1407,17'd269,17'd640,17'd206,17'd642,17'd257,17'd804,17'd252,17'd17075,17'd74570,17'd15626,17'd181,17'd254,17'd801,17'd2255
},
'{
17'd3,17'd3,17'd3,17'd3,17'd979,17'd979,17'd979,17'd979,17'd18,17'd17,17'd466,17'd1127,17'd1689,17'd3250,17'd4887,17'd4246,17'd2782,17'd2593,17'd3751,17'd3901,17'd3901,17'd3751,17'd4244,17'd4891,17'd4891,17'd4087,17'd4736,17'd65710,17'd64927,17'd63977,17'd64929,17'd64929,17'd13576,17'd64254,17'd74571,17'd74571,17'd74572,17'd74572,17'd65714,17'd6739,17'd63821,17'd74573,17'd71425,17'd13302,17'd14441,17'd11607,17'd74574,17'd74574,17'd14441,17'd70076,17'd9683,17'd9683,17'd6267,17'd6104,17'd8669,17'd6102,17'd6102,17'd6589,17'd6106,17'd6103,17'd6267,17'd11736,17'd74575,17'd65313,17'd13185,17'd74232,17'd8983,17'd9552,17'd10668,17'd3249,17'd1830,17'd0,17'd18,17'd3905,17'd3905,17'd18,17'd18,17'd652,17'd29,17'd4431,17'd5971,17'd5804,17'd12931,17'd12507,17'd5808,17'd5383,17'd12038,17'd5222,17'd5521,17'd5659,17'd5976,17'd11345,17'd70077,17'd6903,17'd6903,17'd6744,17'd6903,17'd6903,17'd6902,17'd9275,17'd8988,17'd70686,17'd8197,17'd74462,17'd70288,17'd71521,17'd69810,17'd71092,17'd12200,17'd3913,17'd74576,17'd74577,17'd74578,17'd74579,17'd74580,17'd74581,17'd74582,17'd74583,17'd74584,17'd74585,17'd74586,17'd74587,17'd61454,17'd74121,17'd74588,17'd53959,17'd74356,17'd74357,17'd6160,17'd53889,17'd53090,17'd54181,17'd54545,17'd54716,17'd74360,17'd37977,17'd74479,17'd31750,17'd8227,17'd74481,17'd8390,17'd74589,17'd74589,17'd74589,17'd7432,17'd35220,17'd35220,17'd34026,17'd7594,17'd30357,17'd29906,17'd28671,17'd74590,17'd74591,17'd74592,17'd74593,17'd7597,17'd54364,17'd48934,17'd74594,17'd74595,17'd74596,17'd74597,17'd74598,17'd74599,17'd74600,17'd74601,17'd74602,17'd74603,17'd74604,17'd74605,17'd74606,17'd74607,17'd74608,17'd74609,17'd74610,17'd74611,17'd74612,17'd74613,17'd74501,17'd74614,17'd74615,17'd74616,17'd74617,17'd74618,17'd74619,17'd74620,17'd74621,17'd74622,17'd74623,17'd74624,17'd74625,17'd74626,17'd74627,17'd74515,17'd74628,17'd73393,17'd74629,17'd74629,17'd72652,17'd74630,17'd74631,17'd74632,17'd73723,17'd73076,17'd73075,17'd72866,17'd73497,17'd73073,17'd126,17'd356,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd1481,17'd1481,17'd356,17'd128,17'd132,17'd74633,17'd74634,17'd74635,17'd74636,17'd74637,17'd74528,17'd20821,17'd21441,17'd22058,17'd74638,17'd74639,17'd15833,17'd15321,17'd74533,17'd74533,17'd74640,17'd74641,17'd72052,17'd71962,17'd74642,17'd74643,17'd74644,17'd74645,17'd16608,17'd15599,17'd15333,17'd72889,17'd9386,17'd9653,17'd10229,17'd9389,17'd11176,17'd6849,17'd6550,17'd6847,17'd7169,17'd7169,17'd6215,17'd7176,17'd6851,17'd10236,17'd9932,17'd11430,17'd69787,17'd69787,17'd28306,17'd27932,17'd10897,17'd10897,17'd10897,17'd10897,17'd27932,17'd27932,17'd10642,17'd10515,17'd27933,17'd27933,17'd31551,17'd31889,17'd74646,17'd74647,17'd74538,17'd74425,17'd74539,17'd73521,17'd74648,17'd73199,17'd73410,17'd74649,17'd72059,17'd74650,17'd69602,17'd69328,17'd74075,17'd74651,17'd74652,17'd14304,17'd13283,17'd12473,17'd12008,17'd31892,17'd74653,17'd74654,17'd74655,17'd74656,17'd74657,17'd74658,17'd74659,17'd74660,17'd74660,17'd74661,17'd70369,17'd67658,17'd70369,17'd71398,17'd69236,17'd74662,17'd74663,17'd74664,17'd74665,17'd74561,17'd68178,17'd74445,17'd74666,17'd74666,17'd74667,17'd73756,17'd73976,17'd73866,17'd74668,17'd74447,17'd74669,17'd74670,17'd74099,17'd73981,17'd73761,17'd74222,17'd73981,17'd73981,17'd73321,17'd73322,17'd73763,17'd73321,17'd73870,17'd74562,17'd74671,17'd74671,17'd74097,17'd73536,17'd74101,17'd74672,17'd72170,17'd74566,17'd71295,17'd72166,17'd69419,17'd69336,17'd63808,17'd65054,17'd69338,17'd69526,17'd73427,17'd73986,17'd10395,17'd14060,17'd5357,17'd1824,17'd2587,17'd234,17'd451,17'd784,17'd635,17'd28656,17'd786,17'd790,17'd74673,17'd74674,17'd15492,17'd27824,17'd263,17'd1406,17'd640,17'd2779,17'd260,17'd207,17'd257,17'd1267,17'd74675,17'd41005,17'd426,17'd208,17'd2255,17'd182,17'd74676,17'd74677,17'd74678,17'd20271,17'd2255,17'd974,17'd266,17'd74679
},
'{
17'd3,17'd3,17'd3,17'd3,17'd979,17'd979,17'd979,17'd979,17'd18,17'd3905,17'd466,17'd1127,17'd1689,17'd2781,17'd4887,17'd4246,17'd2784,17'd2782,17'd2593,17'd3751,17'd3751,17'd3751,17'd3903,17'd4244,17'd3902,17'd3902,17'd4427,17'd7042,17'd74680,17'd74681,17'd65066,17'd64929,17'd71195,17'd64254,17'd74682,17'd74683,17'd74684,17'd74685,17'd74459,17'd73109,17'd13433,17'd65189,17'd70777,17'd70680,17'd63387,17'd14441,17'd74686,17'd74574,17'd6433,17'd12783,17'd9552,17'd10662,17'd6102,17'd6102,17'd6106,17'd6102,17'd6101,17'd6102,17'd10662,17'd8194,17'd6433,17'd70076,17'd63667,17'd11453,17'd71714,17'd69723,17'd10402,17'd8823,17'd64668,17'd64400,17'd14742,17'd14,17'd16,17'd3905,17'd20404,17'd1128,17'd18,17'd18,17'd29,17'd29,17'd4430,17'd4430,17'd4431,17'd5971,17'd6278,17'd11889,17'd6110,17'd6110,17'd12931,17'd12931,17'd27445,17'd11211,17'd9555,17'd9275,17'd7061,17'd7061,17'd6903,17'd6903,17'd6902,17'd6902,17'd8988,17'd70686,17'd8197,17'd74462,17'd7729,17'd7729,17'd7559,17'd7227,17'd68756,17'd13068,17'd25902,17'd13952,17'd74687,17'd74688,17'd74689,17'd74690,17'd74691,17'd74692,17'd74693,17'd74694,17'd74695,17'd74696,17'd74697,17'd74698,17'd74699,17'd74700,17'd74701,17'd74702,17'd54101,17'd53960,17'd74703,17'd74704,17'd53306,17'd58175,17'd58545,17'd74705,17'd74706,17'd74707,17'd74708,17'd36618,17'd36618,17'd74709,17'd74709,17'd74710,17'd74710,17'd8550,17'd74711,17'd7595,17'd28802,17'd8082,17'd74712,17'd7928,17'd32274,17'd74713,17'd74593,17'd7597,17'd74714,17'd74715,17'd74716,17'd74717,17'd74718,17'd74719,17'd74720,17'd74721,17'd74722,17'd74723,17'd74724,17'd74725,17'd74726,17'd74727,17'd74728,17'd74729,17'd74730,17'd74731,17'd74732,17'd74733,17'd74734,17'd74735,17'd74736,17'd74502,17'd74737,17'd74738,17'd74739,17'd74740,17'd74741,17'd74742,17'd74743,17'd74744,17'd74745,17'd74746,17'd74747,17'd74748,17'd74749,17'd74750,17'd73606,17'd74751,17'd74752,17'd74753,17'd73075,17'd74754,17'd74755,17'd74632,17'd73835,17'd73834,17'd73724,17'd72984,17'd74756,17'd73612,17'd70217,17'd720,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd1481,17'd1481,17'd128,17'd132,17'd131,17'd74633,17'd74757,17'd74758,17'd74759,17'd74760,17'd74761,17'd29586,17'd74762,17'd74763,17'd74638,17'd74764,17'd13025,17'd15588,17'd74066,17'd73951,17'd74765,17'd74766,17'd73302,17'd72152,17'd74642,17'd74767,17'd74768,17'd74769,17'd16608,17'd16117,17'd74770,17'd74770,17'd9386,17'd9653,17'd10228,17'd10229,17'd10775,17'd11568,17'd6550,17'd6550,17'd7169,17'd7169,17'd6215,17'd6216,17'd6705,17'd10236,17'd9932,17'd11430,17'd69787,17'd69787,17'd28306,17'd28306,17'd10897,17'd10897,17'd10897,17'd10897,17'd11430,17'd10641,17'd10515,17'd10515,17'd27933,17'd27933,17'd31551,17'd29158,17'd31889,17'd74646,17'd74538,17'd74538,17'd73520,17'd73619,17'd73521,17'd73305,17'd74771,17'd73738,17'd72569,17'd72157,17'd72460,17'd70153,17'd74772,17'd74773,17'd74774,17'd74775,17'd74776,17'd74652,17'd74777,17'd74778,17'd74779,17'd74779,17'd74780,17'd74781,17'd68051,17'd74782,17'd74783,17'd74783,17'd74784,17'd68940,17'd68940,17'd74785,17'd74785,17'd74786,17'd71060,17'd74787,17'd74788,17'd74789,17'd74790,17'd74791,17'd74792,17'd74793,17'd74666,17'd74666,17'd74095,17'd73756,17'd73866,17'd73866,17'd74447,17'd74669,17'd74794,17'd74795,17'd74796,17'd74222,17'd74222,17'd74222,17'd73981,17'd73981,17'd73321,17'd73322,17'd73763,17'd73321,17'd73870,17'd73869,17'd74797,17'd74221,17'd74798,17'd72784,17'd72584,17'd72079,17'd71800,17'd74799,17'd71294,17'd69037,17'd70374,17'd66788,17'd64651,17'd68833,17'd69526,17'd66547,17'd65944,17'd58865,17'd48187,17'd37708,17'd11049,17'd4398,17'd1122,17'd1257,17'd784,17'd635,17'd28656,17'd786,17'd766,17'd19864,17'd18868,17'd400,17'd24333,17'd456,17'd263,17'd1406,17'd640,17'd260,17'd260,17'd207,17'd256,17'd263,17'd256,17'd258,17'd208,17'd31100,17'd211,17'd252,17'd16860,17'd74800,17'd74801,17'd253,17'd408,17'd41005,17'd1407,17'd1405
},
'{
17'd12,17'd3,17'd3,17'd283,17'd283,17'd283,17'd979,17'd19,17'd3,17'd12,17'd2,17'd1127,17'd1689,17'd2781,17'd2592,17'd2784,17'd2592,17'd2784,17'd2784,17'd2593,17'd2593,17'd2593,17'd4088,17'd4428,17'd4244,17'd3902,17'd3902,17'd3903,17'd6892,17'd74802,17'd66211,17'd66447,17'd70487,17'd71195,17'd63979,17'd65189,17'd74803,17'd74684,17'd74804,17'd74804,17'd6740,17'd10799,17'd67693,17'd74805,17'd63257,17'd63387,17'd74806,17'd74807,17'd6103,17'd6267,17'd74233,17'd6101,17'd6100,17'd14187,17'd5965,17'd5965,17'd73990,17'd73990,17'd10662,17'd8194,17'd6433,17'd64930,17'd70972,17'd63667,17'd13816,17'd71197,17'd6433,17'd9415,17'd9552,17'd63260,17'd14742,17'd15,17'd16,17'd18,17'd20404,17'd1128,17'd18,17'd19,17'd288,17'd29,17'd28,17'd6744,17'd4431,17'd5971,17'd5971,17'd6746,17'd11889,17'd6110,17'd11737,17'd11889,17'd5803,17'd6598,17'd9555,17'd74808,17'd7728,17'd7061,17'd7556,17'd7225,17'd6902,17'd6902,17'd9275,17'd8988,17'd8197,17'd74462,17'd7729,17'd7729,17'd70288,17'd7063,17'd74809,17'd74810,17'd67069,17'd66817,17'd74811,17'd74812,17'd74813,17'd74814,17'd74815,17'd74816,17'd74817,17'd74818,17'd74819,17'd74820,17'd74821,17'd74822,17'd74823,17'd63018,17'd74824,17'd74825,17'd74826,17'd54028,17'd74827,17'd74828,17'd6160,17'd50193,17'd54031,17'd59161,17'd74829,17'd74830,17'd74831,17'd74831,17'd36925,17'd74832,17'd74832,17'd8390,17'd34026,17'd74833,17'd32114,17'd32426,17'd31428,17'd74712,17'd7767,17'd51422,17'd74146,17'd7597,17'd74834,17'd74835,17'd74836,17'd74837,17'd74838,17'd74839,17'd74840,17'd74841,17'd74842,17'd74843,17'd74844,17'd74845,17'd74846,17'd74847,17'd74848,17'd74849,17'd74850,17'd74851,17'd74852,17'd74853,17'd74854,17'd74855,17'd74856,17'd74857,17'd74858,17'd74859,17'd74741,17'd74860,17'd74861,17'd74861,17'd74862,17'd74863,17'd74864,17'd74865,17'd74866,17'd74867,17'd74868,17'd74869,17'd74870,17'd74871,17'd74872,17'd74751,17'd74873,17'd74874,17'd73721,17'd73610,17'd74523,17'd74875,17'd74876,17'd74877,17'd74878,17'd73072,17'd73612,17'd355,17'd356,17'd132,17'd132,17'd132,17'd132,17'd134,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd1481,17'd1481,17'd134,17'd132,17'd131,17'd73080,17'd74879,17'd74880,17'd74881,17'd74882,17'd74883,17'd32708,17'd74884,17'd74885,17'd74886,17'd74887,17'd15719,17'd13547,17'd74888,17'd73951,17'd74889,17'd74890,17'd73302,17'd74891,17'd74642,17'd74892,17'd74893,17'd74644,17'd16608,17'd74894,17'd74770,17'd9081,17'd15220,17'd9653,17'd10228,17'd10228,17'd11032,17'd68822,17'd6550,17'd6386,17'd6847,17'd7169,17'd6214,17'd6215,17'd6850,17'd10512,17'd11036,17'd11180,17'd11430,17'd69787,17'd27932,17'd27932,17'd10897,17'd10897,17'd10897,17'd10897,17'd10777,17'd10777,17'd27815,17'd27815,17'd27933,17'd27933,17'd27933,17'd28183,17'd31551,17'd29158,17'd74646,17'd74646,17'd74647,17'd73618,17'd73520,17'd73619,17'd73619,17'd74315,17'd73955,17'd73955,17'd73092,17'd72568,17'd72568,17'd70252,17'd74895,17'd74896,17'd74897,17'd74898,17'd74899,17'd74900,17'd74900,17'd74901,17'd74901,17'd74900,17'd74902,17'd74903,17'd74904,17'd74905,17'd73628,17'd74906,17'd74907,17'd72674,17'd74908,17'd72069,17'd74909,17'd74910,17'd74911,17'd74790,17'd74791,17'd74791,17'd74912,17'd74913,17'd74914,17'd74915,17'd74916,17'd74916,17'd74917,17'd74447,17'd74918,17'd74919,17'd74795,17'd74920,17'd74796,17'd74222,17'd74222,17'd73981,17'd74921,17'd73210,17'd73210,17'd73211,17'd73210,17'd74451,17'd74565,17'd74798,17'd73868,17'd74922,17'd73978,17'd74923,17'd74924,17'd74925,17'd74926,17'd70863,17'd69142,17'd69334,17'd70265,17'd63510,17'd66435,17'd64650,17'd66193,17'd73986,17'd7878,17'd6094,17'd37708,17'd4558,17'd4398,17'd628,17'd799,17'd430,17'd441,17'd28656,17'd32882,17'd18633,17'd74927,17'd74928,17'd74929,17'd770,17'd279,17'd1274,17'd1266,17'd74675,17'd257,17'd646,17'd268,17'd2778,17'd459,17'd459,17'd256,17'd257,17'd41316,17'd1093,17'd182,17'd24000,17'd74930,17'd16861,17'd20868,17'd975,17'd262,17'd258,17'd1269,17'd1552
},
'{
17'd12,17'd3,17'd3,17'd283,17'd283,17'd283,17'd19,17'd19,17'd283,17'd3,17'd2,17'd466,17'd1127,17'd1689,17'd2781,17'd3250,17'd3250,17'd3250,17'd2422,17'd2935,17'd2935,17'd2593,17'd3904,17'd4428,17'd3903,17'd3902,17'd3902,17'd3903,17'd3903,17'd6892,17'd69892,17'd74931,17'd64121,17'd64121,17'd71310,17'd12928,17'd74932,17'd74932,17'd74933,17'd74934,17'd6736,17'd6740,17'd13184,17'd71197,17'd12652,17'd9684,17'd10090,17'd74935,17'd6589,17'd6589,17'd74233,17'd6274,17'd5964,17'd14187,17'd67577,17'd6100,17'd5964,17'd63521,17'd6102,17'd6103,17'd10662,17'd6433,17'd11453,17'd67451,17'd69723,17'd13185,17'd64930,17'd63520,17'd8194,17'd69255,17'd12929,17'd3749,17'd16,17'd18,17'd1128,17'd1128,17'd19,17'd19,17'd288,17'd288,17'd28,17'd28,17'd18037,17'd18037,17'd18037,17'd6598,17'd10269,17'd10269,17'd72282,17'd10269,17'd6598,17'd18037,17'd6902,17'd9275,17'd4429,17'd1833,17'd7728,17'd7556,17'd6902,17'd6902,17'd6902,17'd9275,17'd8988,17'd8197,17'd70288,17'd7729,17'd70288,17'd8048,17'd7561,17'd74936,17'd67454,17'd53874,17'd65846,17'd74937,17'd74938,17'd73020,17'd74939,17'd74940,17'd74941,17'd74942,17'd74943,17'd74944,17'd74945,17'd74946,17'd74947,17'd74697,17'd54904,17'd74948,17'd74121,17'd74949,17'd74950,17'd62744,17'd74827,17'd59950,17'd53821,17'd53889,17'd54180,17'd50847,17'd59036,17'd74477,17'd74951,17'd74952,17'd36925,17'd74708,17'd7595,17'd8705,17'd74953,17'd74954,17'd74955,17'd74956,17'd74957,17'd74958,17'd74959,17'd74960,17'd54548,17'd74961,17'd74962,17'd74963,17'd74964,17'd74841,17'd74965,17'd74966,17'd74967,17'd74968,17'd74969,17'd74970,17'd74971,17'd74972,17'd74973,17'd74974,17'd74975,17'd74976,17'd74977,17'd74978,17'd74979,17'd74980,17'd74981,17'd74982,17'd74859,17'd74983,17'd74862,17'd74861,17'd74861,17'd74984,17'd74985,17'd74986,17'd74987,17'd74988,17'd74989,17'd74990,17'd74991,17'd74992,17'd74993,17'd74994,17'd73288,17'd74995,17'd74996,17'd74997,17'd73506,17'd73724,17'd74057,17'd74998,17'd74877,17'd73929,17'd73072,17'd70831,17'd70833,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd1481,17'd1481,17'd134,17'd132,17'd131,17'd72989,17'd74999,17'd75000,17'd75001,17'd75002,17'd75003,17'd75004,17'd60261,17'd75005,17'd75006,17'd75007,17'd15980,17'd13546,17'd75008,17'd73951,17'd75009,17'd75010,17'd75011,17'd74891,17'd75012,17'd74892,17'd75013,17'd74769,17'd74894,17'd16608,17'd72889,17'd9081,17'd9386,17'd9387,17'd10228,17'd10774,17'd9519,17'd11176,17'd68172,17'd6550,17'd6847,17'd7169,17'd6214,17'd6215,17'd7176,17'd10512,17'd11036,17'd11180,17'd11430,17'd71784,17'd27932,17'd27932,17'd27932,17'd10897,17'd10897,17'd10897,17'd10777,17'd10777,17'd27815,17'd27815,17'd27933,17'd27933,17'd27933,17'd27933,17'd30933,17'd30933,17'd30934,17'd31715,17'd75014,17'd75015,17'd74647,17'd75016,17'd75016,17'd75016,17'd75017,17'd75018,17'd75019,17'd72459,17'd72459,17'd72567,17'd75020,17'd75020,17'd71498,17'd70364,17'd69878,17'd69878,17'd75021,17'd75021,17'd75021,17'd69878,17'd68932,17'd75022,17'd75023,17'd68937,17'd74904,17'd75024,17'd75025,17'd69700,17'd75026,17'd75027,17'd75028,17'd74910,17'd74911,17'd75029,17'd74790,17'd74791,17'd75030,17'd74913,17'd74914,17'd74915,17'd74916,17'd74917,17'd75031,17'd74669,17'd75032,17'd75032,17'd74920,17'd74920,17'd75033,17'd74796,17'd73981,17'd73981,17'd73210,17'd73210,17'd74451,17'd74451,17'd73979,17'd74098,17'd75034,17'd74798,17'd74922,17'd74922,17'd75035,17'd75036,17'd75037,17'd74926,17'd71188,17'd75038,17'd69334,17'd64506,17'd71508,17'd63375,17'd69527,17'd67432,17'd65944,17'd70169,17'd6890,17'd13933,17'd6085,17'd4399,17'd628,17'd235,17'd611,17'd27948,17'd39034,17'd434,17'd435,17'd75039,17'd74928,17'd75039,17'd20001,17'd20569,17'd75040,17'd1271,17'd459,17'd74679,17'd266,17'd257,17'd1242,17'd595,17'd265,17'd265,17'd256,17'd1242,17'd1093,17'd593,17'd24000,17'd649,17'd75041,17'd17186,17'd20271,17'd404,17'd1097,17'd207,17'd1269,17'd1552
},
'{
17'd12,17'd12,17'd3,17'd3,17'd1,17'd1,17'd3,17'd3,17'd283,17'd3,17'd12,17'd2,17'd1127,17'd1689,17'd1689,17'd1689,17'd1689,17'd1689,17'd1688,17'd2422,17'd2935,17'd2935,17'd4245,17'd6420,17'd4428,17'd4892,17'd4892,17'd4428,17'd4428,17'd4245,17'd68191,17'd69347,17'd12502,17'd75042,17'd66447,17'd63980,17'd71714,17'd69723,17'd13185,17'd13184,17'd6593,17'd6739,17'd6894,17'd13815,17'd70972,17'd11608,17'd63259,17'd67452,17'd5967,17'd5966,17'd5967,17'd75043,17'd5968,17'd75044,17'd9274,17'd5968,17'd75045,17'd75046,17'd6100,17'd6589,17'd10662,17'd6103,17'd6433,17'd70076,17'd63518,17'd71908,17'd12783,17'd70076,17'd8194,17'd6102,17'd63117,17'd3749,17'd16,17'd18,17'd1128,17'd1128,17'd19,17'd19,17'd19,17'd19,17'd27,17'd27,17'd28,17'd28,17'd288,17'd18037,17'd18037,17'd18037,17'd18037,17'd73110,17'd6902,17'd287,17'd27,17'd286,17'd1833,17'd70686,17'd7556,17'd7556,17'd6903,17'd6903,17'd6902,17'd6902,17'd7728,17'd8047,17'd74462,17'd74462,17'd70288,17'd8048,17'd7227,17'd7561,17'd69988,17'd75047,17'd2945,17'd2267,17'd1707,17'd74938,17'd74346,17'd75048,17'd74239,17'd75049,17'd75050,17'd75051,17'd75052,17'd75053,17'd74818,17'd74946,17'd75054,17'd75055,17'd70706,17'd5856,17'd5706,17'd5706,17'd74699,17'd75056,17'd60807,17'd75057,17'd5863,17'd6018,17'd53614,17'd6648,17'd51103,17'd40735,17'd75058,17'd38608,17'd75059,17'd75060,17'd75061,17'd38226,17'd75062,17'd75063,17'd75064,17'd75065,17'd75066,17'd75067,17'd75068,17'd75069,17'd75070,17'd75071,17'd75072,17'd75073,17'd75074,17'd75075,17'd75076,17'd75077,17'd75078,17'd75079,17'd75080,17'd75081,17'd74975,17'd75082,17'd75083,17'd75084,17'd75085,17'd75086,17'd75087,17'd75088,17'd75089,17'd75090,17'd75091,17'd75092,17'd75093,17'd75094,17'd75094,17'd75095,17'd75096,17'd75097,17'd75098,17'd75099,17'd75100,17'd75101,17'd75102,17'd75103,17'd73935,17'd73392,17'd75104,17'd75105,17'd75106,17'd73721,17'd73290,17'd75107,17'd72551,17'd75108,17'd75109,17'd75110,17'd75111,17'd126,17'd356,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd131,17'd72989,17'd75112,17'd75113,17'd75114,17'd75115,17'd75116,17'd75117,17'd75118,17'd75005,17'd75119,17'd75120,17'd16114,17'd14703,17'd75121,17'd75122,17'd75123,17'd75124,17'd75125,17'd75126,17'd75127,17'd75128,17'd75013,17'd75129,17'd16733,17'd73518,17'd72888,17'd74770,17'd9781,17'd9518,17'd10774,17'd10774,17'd10229,17'd10775,17'd68172,17'd6550,17'd6847,17'd7169,17'd6846,17'd6214,17'd7667,17'd6850,17'd10236,17'd9932,17'd11430,17'd11430,17'd27932,17'd27932,17'd27932,17'd10897,17'd10897,17'd10897,17'd10897,17'd27931,17'd10897,17'd10897,17'd27932,17'd27932,17'd28306,17'd28306,17'd27933,17'd29592,17'd30933,17'd30933,17'd30934,17'd31715,17'd31889,17'd74646,17'd74646,17'd75015,17'd75015,17'd74424,17'd73407,17'd73407,17'd73407,17'd73737,17'd69326,17'd69326,17'd75130,17'd69225,17'd69225,17'd69225,17'd75130,17'd69225,17'd69225,17'd69225,17'd69225,17'd69225,17'd69131,17'd75131,17'd69231,17'd75132,17'd75025,17'd75133,17'd70658,17'd75134,17'd75135,17'd74910,17'd75136,17'd75137,17'd75138,17'd75139,17'd75140,17'd75141,17'd75142,17'd74915,17'd74917,17'd75031,17'd74918,17'd74670,17'd74920,17'd74920,17'd75143,17'd75143,17'd75144,17'd74563,17'd74449,17'd73760,17'd73210,17'd72683,17'd74451,17'd74565,17'd75034,17'd75145,17'd75146,17'd74922,17'd75147,17'd75035,17'd75036,17'd75148,17'd75149,17'd71073,17'd69237,17'd65038,17'd66535,17'd71508,17'd65183,17'd66197,17'd68411,17'd66926,17'd58865,17'd6890,17'd14060,17'd37708,17'd52918,17'd628,17'd798,17'd1379,17'd27948,17'd1541,17'd767,17'd52107,17'd616,17'd617,17'd75150,17'd29442,17'd75151,17'd75152,17'd75153,17'd75154,17'd1271,17'd459,17'd266,17'd1126,17'd456,17'd2115,17'd265,17'd265,17'd255,17'd2255,17'd1682,17'd462,17'd17298,17'd15873,17'd75155,17'd589,17'd461,17'd801,17'd262,17'd968,17'd74456,17'd1552
},
'{
17'd12,17'd12,17'd12,17'd3,17'd1,17'd1,17'd283,17'd283,17'd283,17'd3,17'd3,17'd12,17'd2,17'd1127,17'd1689,17'd1689,17'd1127,17'd1127,17'd1689,17'd1831,17'd3252,17'd2935,17'd4733,17'd4245,17'd4088,17'd4428,17'd4428,17'd4088,17'd4245,17'd6420,17'd6424,17'd12193,17'd74575,17'd12502,17'd65066,17'd65067,17'd12928,17'd71714,17'd69723,17'd65189,17'd6740,17'd69161,17'd7052,17'd7052,17'd71316,17'd11736,17'd12929,17'd14069,17'd75156,17'd75046,17'd5967,17'd75157,17'd9274,17'd11446,17'd5801,17'd75158,17'd5800,17'd6275,17'd75159,17'd6100,17'd6589,17'd6103,17'd10662,17'd64930,17'd63519,17'd70076,17'd9967,17'd70076,17'd6273,17'd10662,17'd74233,17'd63116,17'd14442,17'd16,17'd18,17'd1128,17'd19,17'd19,17'd19,17'd19,17'd27,17'd27,17'd28,17'd28,17'd288,17'd288,17'd288,17'd288,17'd288,17'd70879,17'd2424,17'd287,17'd27,17'd27,17'd1833,17'd4429,17'd8988,17'd7556,17'd9555,17'd6903,17'd6902,17'd6902,17'd7728,17'd7728,17'd8047,17'd74462,17'd71521,17'd70288,17'd8048,17'd7227,17'd7391,17'd70588,17'd72282,17'd3105,17'd1283,17'd2787,17'd75160,17'd74238,17'd75161,17'd75162,17'd75163,17'd75164,17'd75165,17'd75166,17'd75167,17'd75168,17'd75169,17'd75170,17'd75171,17'd75172,17'd75173,17'd75174,17'd75174,17'd75175,17'd75176,17'd75177,17'd75178,17'd75179,17'd61590,17'd53959,17'd43351,17'd75180,17'd52629,17'd51103,17'd50847,17'd50765,17'd54908,17'd54182,17'd75181,17'd54543,17'd58905,17'd58783,17'd75182,17'd75183,17'd75184,17'd75185,17'd75186,17'd75187,17'd75188,17'd75189,17'd75190,17'd75191,17'd75192,17'd75193,17'd75194,17'd75195,17'd75196,17'd75197,17'd75198,17'd75199,17'd75200,17'd75201,17'd75202,17'd75203,17'd75204,17'd75205,17'd75206,17'd75207,17'd75208,17'd75209,17'd75094,17'd75210,17'd75211,17'd75212,17'd75213,17'd75214,17'd75215,17'd75216,17'd75217,17'd75218,17'd75219,17'd73933,17'd75220,17'd75221,17'd75222,17'd75106,17'd74520,17'd73496,17'd73496,17'd73939,17'd73939,17'd75110,17'd72654,17'd71669,17'd126,17'd20762,17'd133,17'd1197,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd131,17'd53482,17'd75223,17'd75224,17'd75225,17'd75226,17'd75227,17'd75228,17'd75229,17'd35328,17'd75230,17'd75231,17'd75232,17'd15586,17'd75233,17'd75234,17'd75235,17'd75010,17'd75236,17'd75237,17'd75238,17'd75239,17'd75013,17'd75240,17'd74644,17'd73736,17'd16950,17'd72889,17'd9652,17'd9518,17'd10774,17'd10774,17'd10228,17'd12002,17'd11850,17'd68172,17'd6386,17'd7169,17'd6846,17'd6703,17'd6214,17'd7176,17'd8000,17'd11036,17'd9932,17'd11430,17'd10897,17'd10897,17'd27932,17'd27932,17'd10897,17'd10897,17'd10897,17'd27931,17'd10897,17'd10897,17'd10897,17'd27932,17'd28306,17'd28306,17'd27933,17'd29592,17'd30933,17'd31551,17'd31551,17'd31715,17'd31889,17'd31889,17'd74646,17'd74646,17'd35340,17'd34922,17'd34922,17'd75241,17'd75241,17'd75241,17'd73090,17'd73090,17'd74424,17'd73407,17'd73407,17'd75130,17'd75130,17'd75130,17'd75130,17'd69130,17'd69411,17'd69512,17'd69227,17'd75131,17'd69136,17'd75024,17'd75242,17'd75133,17'd70658,17'd75134,17'd75243,17'd75244,17'd75245,17'd75246,17'd75247,17'd75248,17'd75141,17'd74914,17'd75249,17'd75250,17'd75251,17'd74918,17'd74795,17'd74795,17'd74920,17'd75033,17'd75144,17'd75144,17'd75144,17'd74563,17'd74449,17'd73870,17'd72683,17'd74451,17'd74565,17'd75034,17'd74333,17'd74333,17'd75146,17'd73867,17'd75147,17'd75252,17'd75148,17'd75149,17'd72166,17'd65552,17'd65419,17'd66063,17'd71508,17'd63375,17'd66197,17'd68295,17'd67433,17'd67048,17'd6890,17'd13933,17'd37821,17'd5497,17'd628,17'd235,17'd1379,17'd23643,17'd51335,17'd18515,17'd75253,17'd618,17'd75254,17'd217,17'd75255,17'd75256,17'd23489,17'd252,17'd15240,17'd1270,17'd1274,17'd459,17'd1274,17'd456,17'd254,17'd804,17'd1270,17'd265,17'd2255,17'd1682,17'd612,17'd68749,17'd16635,17'd75257,17'd75258,17'd591,17'd20008,17'd1097,17'd256,17'd1268,17'd75259,17'd1552
},
'{
17'd12,17'd12,17'd0,17'd0,17'd0,17'd1,17'd283,17'd283,17'd283,17'd283,17'd3,17'd12,17'd2,17'd2,17'd1127,17'd1127,17'd466,17'd466,17'd1127,17'd1688,17'd2422,17'd2784,17'd6584,17'd4733,17'd3904,17'd4428,17'd4428,17'd4428,17'd4245,17'd4245,17'd2935,17'd75260,17'd12332,17'd72694,17'd71085,17'd71085,17'd63980,17'd63821,17'd63822,17'd65189,17'd71615,17'd11885,17'd8043,17'd8043,17'd6894,17'd63980,17'd10801,17'd63117,17'd75261,17'd9274,17'd5968,17'd75158,17'd75262,17'd5653,17'd75263,17'd75263,17'd75263,17'd75262,17'd75158,17'd5968,17'd6596,17'd8042,17'd5965,17'd6589,17'd63387,17'd63519,17'd11736,17'd9967,17'd10923,17'd73990,17'd5964,17'd62981,17'd1277,17'd16,17'd18,17'd18,17'd1128,17'd11,17'd19,17'd19,17'd27,17'd27,17'd11,17'd11,17'd19,17'd19,17'd19,17'd19,17'd19,17'd19,17'd979,17'd979,17'd286,17'd27,17'd286,17'd7061,17'd7388,17'd7557,17'd7556,17'd7556,17'd6902,17'd6902,17'd7061,17'd7728,17'd8047,17'd8047,17'd74462,17'd70288,17'd70288,17'd7557,17'd8048,17'd70687,17'd8988,17'd9554,17'd14447,17'd75264,17'd75265,17'd75266,17'd75267,17'd75268,17'd75269,17'd75270,17'd75271,17'd75272,17'd75273,17'd75274,17'd75275,17'd75276,17'd75169,17'd75277,17'd75277,17'd75278,17'd75278,17'd75279,17'd75280,17'd75281,17'd75282,17'd75283,17'd75284,17'd75285,17'd75286,17'd75287,17'd75288,17'd75289,17'd75290,17'd75291,17'd75292,17'd75293,17'd75294,17'd75295,17'd75296,17'd75297,17'd75298,17'd75299,17'd75300,17'd75301,17'd75302,17'd75303,17'd75304,17'd75305,17'd75306,17'd75307,17'd75308,17'd75309,17'd75310,17'd75311,17'd75312,17'd75313,17'd75314,17'd75315,17'd75316,17'd75317,17'd75318,17'd75319,17'd75320,17'd75321,17'd75091,17'd75322,17'd75323,17'd75324,17'd75325,17'd75326,17'd75327,17'd75328,17'd75329,17'd75330,17'd75331,17'd75332,17'd75333,17'd75334,17'd75335,17'd74751,17'd75336,17'd74754,17'd74520,17'd75337,17'd73075,17'd75338,17'd75108,17'd75110,17'd72654,17'd71765,17'd75339,17'd75340,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd131,17'd17139,17'd72038,17'd75341,17'd75342,17'd75343,17'd75344,17'd75345,17'd75346,17'd75347,17'd75348,17'd75349,17'd75350,17'd75351,17'd17035,17'd75352,17'd75235,17'd75010,17'd75353,17'd75354,17'd75240,17'd75355,17'd75356,17'd75357,17'd74769,17'd73736,17'd74894,17'd15599,17'd9652,17'd9781,17'd9781,17'd10228,17'd75358,17'd12621,17'd12003,17'd11849,17'd6386,17'd6386,17'd7169,17'd7167,17'd6214,17'd7667,17'd8932,17'd68621,17'd9932,17'd9932,17'd10777,17'd10777,17'd10897,17'd27932,17'd27932,17'd10897,17'd10897,17'd27931,17'd10513,17'd10513,17'd10897,17'd10897,17'd10897,17'd10897,17'd27932,17'd27932,17'd27933,17'd28183,17'd28183,17'd29158,17'd29158,17'd34792,17'd34792,17'd35340,17'd30488,17'd30488,17'd30488,17'd37559,17'd34922,17'd34922,17'd73090,17'd73197,17'd69511,17'd69029,17'd69129,17'd68932,17'd68932,17'd70651,17'd70651,17'd75022,17'd69228,17'd69230,17'd75359,17'd69136,17'd69415,17'd75242,17'd69792,17'd70159,17'd70658,17'd75134,17'd75243,17'd75360,17'd75361,17'd75362,17'd75247,17'd75363,17'd75364,17'd75365,17'd75366,17'd75367,17'd75368,17'd75369,17'd75143,17'd75370,17'd75371,17'd75371,17'd74223,17'd74223,17'd74099,17'd74099,17'd73980,17'd74336,17'd73642,17'd74226,17'd75034,17'd74333,17'd75372,17'd75373,17'd75374,17'd75147,17'd75036,17'd75148,17'd75375,17'd67664,17'd64902,17'd66180,17'd66064,17'd72268,17'd63375,17'd63243,17'd63372,17'd67433,17'd67048,17'd14858,17'd13933,17'd37821,17'd1824,17'd4059,17'd630,17'd36748,17'd23814,17'd38863,17'd35208,17'd16263,17'd30945,17'd75376,17'd39036,17'd438,17'd16263,17'd75377,17'd23489,17'd24333,17'd15240,17'd254,17'd1274,17'd1274,17'd27824,17'd17789,17'd17789,17'd15240,17'd1684,17'd1684,17'd965,17'd182,17'd68847,17'd75378,17'd75379,17'd75380,17'd15872,17'd634,17'd429,17'd1097,17'd257,17'd1269,17'd75259,17'd1273
},
'{
17'd3,17'd12,17'd0,17'd0,17'd0,17'd1,17'd283,17'd650,17'd283,17'd283,17'd3,17'd3,17'd0,17'd2,17'd1127,17'd1127,17'd2595,17'd466,17'd1127,17'd1688,17'd3250,17'd2592,17'd27591,17'd6584,17'd3904,17'd4088,17'd4892,17'd4428,17'd4245,17'd4245,17'd2935,17'd2784,17'd6265,17'd11608,17'd63667,17'd71085,17'd65189,17'd12928,17'd12928,17'd12928,17'd64122,17'd70070,17'd8043,17'd68645,17'd67574,17'd6740,17'd71714,17'd73540,17'd63118,17'd75157,17'd5801,17'd5799,17'd75263,17'd3748,17'd5651,17'd5651,17'd808,17'd6108,17'd75263,17'd5799,17'd6266,17'd6428,17'd6428,17'd6434,17'd6102,17'd63386,17'd9684,17'd10923,17'd64668,17'd14867,17'd5964,17'd6107,17'd14442,17'd16,17'd18,17'd18,17'd1128,17'd11,17'd19,17'd19,17'd27,17'd27,17'd11,17'd11,17'd19,17'd19,17'd19,17'd19,17'd19,17'd19,17'd19,17'd979,17'd286,17'd286,17'd286,17'd7060,17'd7555,17'd7557,17'd9276,17'd7556,17'd6902,17'd6902,17'd7061,17'd7061,17'd8988,17'd7555,17'd8047,17'd75381,17'd71521,17'd73111,17'd73111,17'd75381,17'd75381,17'd71091,17'd75382,17'd75383,17'd75384,17'd75385,17'd75386,17'd75387,17'd75388,17'd75389,17'd75390,17'd75391,17'd75392,17'd75393,17'd75394,17'd75395,17'd75396,17'd75397,17'd75398,17'd75398,17'd75399,17'd75400,17'd75401,17'd75401,17'd75402,17'd75403,17'd75404,17'd75405,17'd75406,17'd75407,17'd75408,17'd75408,17'd75409,17'd75410,17'd75411,17'd75412,17'd75413,17'd75414,17'd75415,17'd75416,17'd75417,17'd75418,17'd75419,17'd75420,17'd75421,17'd75422,17'd75423,17'd75424,17'd75425,17'd75426,17'd75427,17'd75428,17'd75429,17'd75430,17'd75431,17'd75432,17'd75433,17'd75434,17'd75435,17'd75436,17'd75437,17'd75438,17'd75439,17'd74983,17'd75440,17'd75441,17'd75442,17'd75443,17'd75326,17'd75328,17'd75444,17'd75444,17'd75445,17'd75446,17'd75447,17'd75448,17'd75449,17'd75450,17'd73713,17'd75222,17'd73506,17'd73833,17'd73394,17'd73724,17'd75451,17'd74051,17'd75452,17'd75453,17'd73184,17'd70437,17'd52246,17'd11541,17'd132,17'd134,17'd128,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd131,17'd5593,17'd75454,17'd75455,17'd75456,17'd75457,17'd75458,17'd75459,17'd75460,17'd75461,17'd75462,17'd75463,17'd50584,17'd75464,17'd75465,17'd75466,17'd75235,17'd75467,17'd75468,17'd75469,17'd74893,17'd75470,17'd75356,17'd75356,17'd74768,17'd73736,17'd16950,17'd15600,17'd9781,17'd10774,17'd9651,17'd10228,17'd75358,17'd75358,17'd12302,17'd11849,17'd6385,17'd6385,17'd7169,17'd7167,17'd6213,17'd6214,17'd7176,17'd68621,17'd9932,17'd9932,17'd10777,17'd10777,17'd10897,17'd27932,17'd27932,17'd10897,17'd10897,17'd27931,17'd10513,17'd10513,17'd27931,17'd27931,17'd10897,17'd10897,17'd27932,17'd27932,17'd27933,17'd27933,17'd27933,17'd28183,17'd29158,17'd29158,17'd34792,17'd34792,17'd30639,17'd30639,17'd30639,17'd37431,17'd35340,17'd74646,17'd73197,17'd75471,17'd69225,17'd69411,17'd69512,17'd70651,17'd75022,17'd75021,17'd75021,17'd75023,17'd75472,17'd69032,17'd69232,17'd75473,17'd69699,17'd73097,17'd69792,17'd70159,17'd69608,17'd75474,17'd75135,17'd75244,17'd75361,17'd75475,17'd75363,17'd75364,17'd75365,17'd75476,17'd75477,17'd75478,17'd75479,17'd75143,17'd75370,17'd75480,17'd75371,17'd75371,17'd74223,17'd75144,17'd74796,17'd74099,17'd73980,17'd74335,17'd74565,17'd75034,17'd74333,17'd73756,17'd75481,17'd75373,17'd75374,17'd75482,17'd75483,17'd72168,17'd67420,17'd69141,17'd64089,17'd64227,17'd66306,17'd66789,17'd63243,17'd64386,17'd63104,17'd67434,17'd75484,17'd48187,17'd37708,17'd4558,17'd38071,17'd38856,17'd36748,17'd24496,17'd1378,17'd33696,17'd29753,17'd75255,17'd39036,17'd32884,17'd39036,17'd586,17'd767,17'd75485,17'd612,17'd639,17'd1123,17'd804,17'd456,17'd254,17'd73644,17'd402,17'd15626,17'd252,17'd15240,17'd965,17'd186,17'd462,17'd75486,17'd39629,17'd75487,17'd75488,17'd250,17'd610,17'd1539,17'd41005,17'd968,17'd275,17'd1411,17'd72687
},
'{
17'd12,17'd12,17'd0,17'd2,17'd2,17'd1,17'd1412,17'd1,17'd283,17'd283,17'd1275,17'd806,17'd3,17'd12,17'd2,17'd466,17'd466,17'd2,17'd14,17'd1127,17'd1688,17'd2422,17'd4887,17'd27591,17'd3904,17'd3904,17'd4088,17'd4088,17'd2934,17'd2934,17'd2935,17'd3252,17'd1688,17'd9815,17'd70874,17'd71085,17'd75489,17'd11886,17'd13433,17'd13815,17'd63978,17'd71708,17'd67574,17'd8043,17'd12191,17'd12033,17'd13815,17'd9967,17'd9553,17'd9422,17'd75490,17'd75158,17'd5653,17'd16389,17'd25,17'd9,17'd25,17'd16389,17'd5652,17'd5651,17'd6276,17'd5800,17'd11730,17'd6428,17'd6434,17'd63258,17'd10668,17'd64125,17'd64125,17'd64125,17'd75156,17'd6275,17'd75491,17'd1277,17'd3905,17'd18,17'd11,17'd1128,17'd18,17'd19,17'd286,17'd285,17'd286,17'd286,17'd10,17'd11,17'd11,17'd11,17'd10,17'd10,17'd10,17'd10,17'd1833,17'd1833,17'd7061,17'd7060,17'd20570,17'd20570,17'd7728,17'd7728,17'd9275,17'd9275,17'd6902,17'd7060,17'd7060,17'd7385,17'd8047,17'd8197,17'd75381,17'd75381,17'd74462,17'd75492,17'd51860,17'd8197,17'd75493,17'd14077,17'd75494,17'd75495,17'd75496,17'd75497,17'd75498,17'd75499,17'd1297,17'd1015,17'd75500,17'd75501,17'd75502,17'd75503,17'd75504,17'd75505,17'd75506,17'd75507,17'd75508,17'd75509,17'd75510,17'd75511,17'd75512,17'd75398,17'd75513,17'd75514,17'd75515,17'd75515,17'd75516,17'd75517,17'd75400,17'd75518,17'd75519,17'd75520,17'd75521,17'd75522,17'd75523,17'd75524,17'd75525,17'd75526,17'd75527,17'd75528,17'd75529,17'd75530,17'd75531,17'd75309,17'd75532,17'd75533,17'd75534,17'd75535,17'd75536,17'd75537,17'd75538,17'd75538,17'd75539,17'd75540,17'd75541,17'd75542,17'd75543,17'd74615,17'd75544,17'd75545,17'd75441,17'd75546,17'd75547,17'd75548,17'd75549,17'd75550,17'd75551,17'd75552,17'd75553,17'd75554,17'd75555,17'd75556,17'd73831,17'd75557,17'd75558,17'd74754,17'd73290,17'd75559,17'd73836,17'd75560,17'd73836,17'd73178,17'd72987,17'd73388,17'd67858,17'd134,17'd11541,17'd131,17'd131,17'd130,17'd136,17'd136,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd133,17'd131,17'd74633,17'd75561,17'd75562,17'd75563,17'd29732,17'd30025,17'd75564,17'd75565,17'd75566,17'd75567,17'd75568,17'd75569,17'd75570,17'd75571,17'd75572,17'd75573,17'd75353,17'd75574,17'd75575,17'd75575,17'd74893,17'd75357,17'd75576,17'd73736,17'd15600,17'd16117,17'd10773,17'd10229,17'd9652,17'd10229,17'd12758,17'd12621,17'd75577,17'd11851,17'd6386,17'd6386,17'd7169,17'd7169,17'd7991,17'd7168,17'd7667,17'd6850,17'd10236,17'd11036,17'd9932,17'd9932,17'd10777,17'd10641,17'd27932,17'd27932,17'd10897,17'd10897,17'd10513,17'd10513,17'd10777,17'd10777,17'd10777,17'd10777,17'd10897,17'd10897,17'd9933,17'd27815,17'd27815,17'd10515,17'd28183,17'd28183,17'd28057,17'd27934,17'd29158,17'd34792,17'd35340,17'd74646,17'd73090,17'd74424,17'd69225,17'd69225,17'd69969,17'd69969,17'd69969,17'd75020,17'd69327,17'd69327,17'd69328,17'd69328,17'd75578,17'd75579,17'd75579,17'd75580,17'd75581,17'd75582,17'd75025,17'd75583,17'd72674,17'd74908,17'd75134,17'd75584,17'd75585,17'd75139,17'd75586,17'd75141,17'd75587,17'd75588,17'd75589,17'd75590,17'd75591,17'd75592,17'd75371,17'd74223,17'd75371,17'd75371,17'd74796,17'd74796,17'd74796,17'd74670,17'd74794,17'd74669,17'd74917,17'd75593,17'd73754,17'd73754,17'd75372,17'd75373,17'd73317,17'd72906,17'd72167,17'd67420,17'd69141,17'd67552,17'd67037,17'd63941,17'd71596,17'd62972,17'd63372,17'd66194,17'd66070,17'd44850,17'd14060,17'd37708,17'd5497,17'd4398,17'd1121,17'd3071,17'd36323,17'd22435,17'd75594,17'd51582,17'd19240,17'd75595,17'd75596,17'd32884,17'd31103,17'd15874,17'd75597,17'd75151,17'd15626,17'd639,17'd26728,17'd804,17'd804,17'd50187,17'd402,17'd1826,17'd24333,17'd180,17'd17789,17'd18271,17'd1826,17'd24000,17'd75598,17'd75599,17'd75600,17'd15873,17'd933,17'd3100,17'd1539,17'd261,17'd968,17'd275,17'd1551,17'd3747
},
'{
17'd12,17'd3,17'd0,17'd2,17'd2,17'd0,17'd1,17'd1,17'd283,17'd283,17'd1275,17'd806,17'd3,17'd12,17'd2,17'd2,17'd466,17'd2,17'd14,17'd14,17'd1688,17'd2422,17'd4887,17'd27591,17'd6264,17'd3904,17'd3904,17'd4088,17'd2934,17'd2934,17'd3101,17'd3252,17'd1831,17'd1967,17'd63257,17'd67451,17'd12502,17'd11886,17'd71615,17'd13433,17'd13433,17'd71310,17'd70070,17'd68645,17'd68645,17'd67574,17'd64254,17'd13184,17'd63258,17'd67308,17'd9422,17'd75491,17'd75263,17'd5652,17'd9,17'd9,17'd9,17'd9,17'd9,17'd9,17'd5651,17'd6276,17'd6731,17'd6266,17'd5962,17'd67577,17'd14069,17'd12929,17'd63260,17'd64125,17'd75261,17'd75043,17'd67308,17'd1276,17'd18,17'd18,17'd11,17'd1128,17'd18,17'd19,17'd286,17'd285,17'd286,17'd286,17'd10,17'd10,17'd11,17'd11,17'd11,17'd11,17'd11,17'd10,17'd286,17'd286,17'd7061,17'd7060,17'd7060,17'd20570,17'd7061,17'd7728,17'd9275,17'd9275,17'd6902,17'd6902,17'd6744,17'd7061,17'd7728,17'd8047,17'd8197,17'd74462,17'd75492,17'd75492,17'd51941,17'd74462,17'd8198,17'd71317,17'd75601,17'd75602,17'd75603,17'd75604,17'd75605,17'd75606,17'd61036,17'd58382,17'd75607,17'd75608,17'd75609,17'd75610,17'd75611,17'd75612,17'd75613,17'd75614,17'd75615,17'd75616,17'd75617,17'd75618,17'd75508,17'd75619,17'd75620,17'd75621,17'd75622,17'd75623,17'd75509,17'd75624,17'd75624,17'd75625,17'd75626,17'd75627,17'd75628,17'd75629,17'd75630,17'd75631,17'd75632,17'd75633,17'd75634,17'd75635,17'd75636,17'd75637,17'd75638,17'd75639,17'd75640,17'd75641,17'd75642,17'd75538,17'd75643,17'd75644,17'd75644,17'd75645,17'd75646,17'd75647,17'd75648,17'd75649,17'd75650,17'd75651,17'd75652,17'd75653,17'd75654,17'd75655,17'd75655,17'd75656,17'd75657,17'd75658,17'd75659,17'd75660,17'd75661,17'd75662,17'd75663,17'd75664,17'd74402,17'd75665,17'd74632,17'd73724,17'd72985,17'd75666,17'd73939,17'd72986,17'd73497,17'd75667,17'd75668,17'd70538,17'd128,17'd11541,17'd131,17'd131,17'd132,17'd130,17'd136,17'd136,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd133,17'd132,17'd20189,17'd75669,17'd75670,17'd75671,17'd75672,17'd75673,17'd75674,17'd75675,17'd75676,17'd75677,17'd57220,17'd52601,17'd75678,17'd17652,17'd75572,17'd75573,17'd75353,17'd75679,17'd18370,17'd75575,17'd74893,17'd75356,17'd75575,17'd73518,17'd15600,17'd15600,17'd9518,17'd10229,17'd10229,17'd10228,17'd75358,17'd12621,17'd12159,17'd12003,17'd6551,17'd6386,17'd6847,17'd7169,17'd75680,17'd7991,17'd7667,17'd6850,17'd10236,17'd10236,17'd9932,17'd9932,17'd10777,17'd10641,17'd27932,17'd27932,17'd10897,17'd10897,17'd9657,17'd9657,17'd10513,17'd10513,17'd10777,17'd10777,17'd10897,17'd10897,17'd27815,17'd10515,17'd10515,17'd10515,17'd27933,17'd27933,17'd28183,17'd28183,17'd34792,17'd31889,17'd74646,17'd73090,17'd73090,17'd73407,17'd69411,17'd69411,17'd72890,17'd72890,17'd72890,17'd69969,17'd69969,17'd69969,17'd69327,17'd75131,17'd69135,17'd69032,17'd69032,17'd69032,17'd75580,17'd75580,17'd75581,17'd75681,17'd75583,17'd74908,17'd75028,17'd75682,17'd75029,17'd74791,17'd75140,17'd75683,17'd75684,17'd75685,17'd75686,17'd75687,17'd75591,17'd75592,17'd75143,17'd75144,17'd75144,17'd75144,17'd74795,17'd74795,17'd74919,17'd74918,17'd75031,17'd74917,17'd75688,17'd75689,17'd73865,17'd74094,17'd75481,17'd73207,17'd73008,17'd75690,17'd67420,17'd66914,17'd69141,17'd63940,17'd65165,17'd65040,17'd62974,17'd63372,17'd67433,17'd65945,17'd44850,17'd16492,17'd5373,17'd4558,17'd4398,17'd796,17'd52461,17'd35059,17'd22435,17'd21944,17'd51582,17'd75253,17'd75691,17'd75692,17'd75693,17'd75376,17'd586,17'd16387,17'd463,17'd24332,17'd15626,17'd1683,17'd1683,17'd186,17'd186,17'd402,17'd1548,17'd1826,17'd638,17'd213,17'd1683,17'd24333,17'd638,17'd35208,17'd75694,17'd75695,17'd75488,17'd17186,17'd404,17'd1539,17'd426,17'd640,17'd1407,17'd1269,17'd1411,17'd70275
},
'{
17'd12,17'd3,17'd1,17'd2,17'd1127,17'd14,17'd1,17'd1412,17'd283,17'd283,17'd1275,17'd1275,17'd19,17'd18,17'd18,17'd3905,17'd466,17'd2,17'd14,17'd14,17'd1689,17'd3250,17'd4577,17'd4577,17'd27591,17'd6584,17'd4733,17'd4245,17'd2934,17'd2934,17'd2934,17'd3101,17'd2594,17'd4247,17'd3750,17'd12652,17'd11343,17'd65068,17'd63820,17'd63820,17'd67306,17'd71615,17'd71708,17'd66815,17'd12033,17'd67574,17'd66815,17'd6735,17'd6267,17'd63669,17'd3749,17'd1,17'd75696,17'd5652,17'd9,17'd9,17'd1690,17'd1691,17'd23,17'd21,17'd25,17'd5651,17'd5794,17'd6436,17'd7381,17'd5962,17'd67695,17'd63116,17'd63116,17'd63118,17'd9553,17'd67308,17'd75490,17'd1276,17'd19,17'd18,17'd18,17'd18,17'd18,17'd11,17'd285,17'd285,17'd285,17'd285,17'd285,17'd285,17'd20,17'd20,17'd11,17'd1128,17'd27,17'd27,17'd286,17'd286,17'd287,17'd27,17'd7061,17'd7060,17'd7060,17'd7061,17'd9275,17'd9275,17'd75697,17'd6902,17'd6744,17'd7061,17'd7061,17'd7555,17'd8047,17'd52025,17'd75492,17'd75492,17'd70288,17'd73111,17'd7729,17'd8048,17'd7391,17'd75047,17'd3106,17'd41008,17'd75698,17'd75699,17'd75700,17'd62583,17'd57373,17'd75701,17'd75702,17'd75703,17'd75704,17'd75705,17'd75706,17'd75707,17'd75708,17'd75709,17'd75710,17'd75711,17'd75615,17'd75712,17'd75712,17'd75712,17'd75713,17'd75713,17'd75714,17'd75715,17'd75716,17'd75717,17'd75718,17'd75719,17'd75720,17'd75721,17'd75722,17'd75723,17'd75724,17'd75725,17'd75726,17'd75727,17'd75728,17'd75729,17'd75730,17'd75731,17'd75732,17'd75733,17'd75734,17'd75735,17'd75736,17'd75737,17'd75738,17'd75739,17'd75740,17'd75741,17'd75742,17'd75743,17'd75744,17'd75745,17'd75746,17'd75747,17'd75748,17'd75749,17'd75750,17'd75751,17'd75752,17'd75753,17'd75754,17'd75661,17'd75755,17'd75756,17'd75757,17'd75758,17'd75759,17'd75760,17'd75761,17'd74521,17'd73836,17'd73939,17'd73497,17'd75762,17'd73388,17'd71260,17'd70438,17'd130,17'd132,17'd131,17'd131,17'd132,17'd132,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd134,17'd133,17'd132,17'd6531,17'd6532,17'd75763,17'd75764,17'd75765,17'd31542,17'd75766,17'd75767,17'd75768,17'd75769,17'd22570,17'd56530,17'd17372,17'd75770,17'd75771,17'd75573,17'd18130,17'd18497,17'd18618,17'd75772,17'd75240,17'd75357,17'd75240,17'd74769,17'd19477,17'd75773,17'd14044,17'd9929,17'd11031,17'd10228,17'd12156,17'd12758,17'd12159,17'd12302,17'd11851,17'd6386,17'd7826,17'd7169,17'd75680,17'd75680,17'd8931,17'd7176,17'd10236,17'd10236,17'd9931,17'd9932,17'd10777,17'd10777,17'd10641,17'd10641,17'd10897,17'd10897,17'd9657,17'd8304,17'd8304,17'd9657,17'd10513,17'd10777,17'd10897,17'd10897,17'd10515,17'd10515,17'd10515,17'd27815,17'd27815,17'd27815,17'd10516,17'd68928,17'd68929,17'd68724,17'd68825,17'd68824,17'd69325,17'd69410,17'd69410,17'd69410,17'd73197,17'd69029,17'd69029,17'd69029,17'd69129,17'd71497,17'd71497,17'd70651,17'd75021,17'd75021,17'd75774,17'd75774,17'd75775,17'd75775,17'd69032,17'd75580,17'd75582,17'd75776,17'd74786,17'd75777,17'd75778,17'd75779,17'd75030,17'd75780,17'd75781,17'd75782,17'd75783,17'd75784,17'd75590,17'd75785,17'd75369,17'd75369,17'd75479,17'd75368,17'd75786,17'd75786,17'd75787,17'd75788,17'd73756,17'd73636,17'd74444,17'd74444,17'd74443,17'd74332,17'd67915,17'd73008,17'd72167,17'd67549,17'd65037,17'd69141,17'd67285,17'd65041,17'd63942,17'd66322,17'd66927,17'd63104,17'd67048,17'd64525,17'd14060,17'd37708,17'd64647,17'd4398,17'd235,17'd36748,17'd36323,17'd2419,17'd21944,17'd21324,17'd20265,17'd75789,17'd75790,17'd75791,17'd75792,17'd31904,17'd221,17'd16496,17'd463,17'd24332,17'd15626,17'd15626,17'd15626,17'd251,17'd250,17'd250,17'd250,17'd251,17'd251,17'd213,17'd15492,17'd252,17'd75151,17'd15742,17'd30193,17'd75380,17'd75793,17'd612,17'd2588,17'd207,17'd2779,17'd1829,17'd1411,17'd14597,17'd206,17'd8188
},
'{
17'd12,17'd3,17'd1,17'd0,17'd1127,17'd1127,17'd0,17'd1412,17'd1412,17'd283,17'd283,17'd1275,17'd19,17'd19,17'd18,17'd18,17'd2,17'd2,17'd14,17'd14,17'd1689,17'd1689,17'd7711,17'd4577,17'd4577,17'd27591,17'd4733,17'd4733,17'd2934,17'd2934,17'd2934,17'd3101,17'd1831,17'd1831,17'd3250,17'd9968,17'd63519,17'd72694,17'd69723,17'd65189,17'd12928,17'd12928,17'd63978,17'd64929,17'd64254,17'd12033,17'd67574,17'd64254,17'd9419,17'd73990,17'd14069,17'd3749,17'd1276,17'd3748,17'd16389,17'd1413,17'd2937,17'd1691,17'd22,17'd22,17'd25,17'd9,17'd6277,17'd5794,17'd13941,17'd7381,17'd16865,17'd14988,17'd1127,17'd3249,17'd9553,17'd14442,17'd75491,17'd5969,17'd19,17'd18,17'd18,17'd18,17'd18,17'd19,17'd286,17'd285,17'd285,17'd285,17'd285,17'd285,17'd21,17'd21,17'd1128,17'd1128,17'd980,17'd27,17'd286,17'd286,17'd287,17'd287,17'd286,17'd7060,17'd7060,17'd7060,17'd6902,17'd9275,17'd75697,17'd73110,17'd6902,17'd6902,17'd6902,17'd7061,17'd7728,17'd8047,17'd74462,17'd74462,17'd70288,17'd73111,17'd75794,17'd70288,17'd8198,17'd7391,17'd68646,17'd5658,17'd3106,17'd14078,17'd75494,17'd75495,17'd75795,17'd56893,17'd75796,17'd75797,17'd75798,17'd75799,17'd75800,17'd861,17'd75801,17'd75802,17'd75803,17'd75804,17'd75805,17'd75806,17'd75807,17'd75807,17'd75807,17'd75808,17'd75809,17'd75810,17'd75811,17'd75812,17'd75813,17'd75814,17'd75815,17'd75816,17'd75817,17'd75818,17'd75819,17'd75820,17'd75821,17'd75822,17'd75823,17'd75824,17'd75825,17'd75826,17'd75827,17'd75828,17'd75829,17'd75830,17'd75831,17'd75832,17'd75833,17'd75834,17'd75835,17'd75836,17'd75837,17'd75838,17'd75839,17'd75747,17'd75840,17'd75750,17'd75841,17'd75842,17'd75843,17'd75844,17'd75845,17'd75846,17'd75847,17'd75848,17'd75849,17'd75850,17'd75851,17'd75852,17'd73503,17'd75853,17'd75854,17'd74877,17'd73178,17'd73072,17'd73074,17'd71954,17'd72754,17'd356,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd134,17'd133,17'd133,17'd15202,17'd2865,17'd75855,17'd75856,17'd75857,17'd75858,17'd75859,17'd75860,17'd75861,17'd75566,17'd43179,17'd23098,17'd75862,17'd75863,17'd75864,17'd75865,17'd75866,17'd18497,17'd74894,17'd75867,17'd75576,17'd75240,17'd74893,17'd74768,17'd15983,17'd15220,17'd14044,17'd14044,17'd11031,17'd10229,17'd75358,17'd12621,17'd75577,17'd12158,17'd11851,17'd11849,17'd6550,17'd7169,17'd7991,17'd75680,17'd75868,17'd8931,17'd8000,17'd10236,17'd9931,17'd9932,17'd10513,17'd10777,17'd10777,17'd10777,17'd10897,17'd10897,17'd10513,17'd9657,17'd8304,17'd8304,17'd9657,17'd10513,17'd10897,17'd27931,17'd27815,17'd27815,17'd27815,17'd27815,17'd9933,17'd27815,17'd10516,17'd10778,17'd72255,17'd72058,17'd72058,17'd68623,17'd68510,17'd68510,17'd68510,17'd68510,17'd68622,17'd68824,17'd68824,17'd68824,17'd68824,17'd69325,17'd69325,17'd69325,17'd69511,17'd69030,17'd75022,17'd75023,17'd75774,17'd75775,17'd69032,17'd75581,17'd75582,17'd75776,17'd74786,17'd75777,17'd75869,17'd75870,17'd75871,17'd75872,17'd75873,17'd75874,17'd75875,17'd75876,17'd75686,17'd75877,17'd75877,17'd75686,17'd75686,17'd75878,17'd75879,17'd75880,17'd74666,17'd74445,17'd75881,17'd75882,17'd74664,17'd75883,17'd75884,17'd74332,17'd68832,17'd67786,17'd73863,17'd65551,17'd69141,17'd63940,17'd65041,17'd15482,17'd68416,17'd16959,17'd63104,17'd65945,17'd10395,17'd48187,17'd37708,17'd4558,17'd4398,17'd628,17'd6867,17'd36323,17'd18386,17'd31099,17'd21467,17'd32405,17'd585,17'd75790,17'd75885,17'd75886,17'd75376,17'd219,17'd16387,17'd16634,17'd1542,17'd770,17'd21165,17'd770,17'd280,17'd589,17'd17423,17'd1543,17'd250,17'd250,17'd250,17'd251,17'd251,17'd280,17'd15742,17'd16635,17'd16005,17'd75887,17'd400,17'd404,17'd935,17'd270,17'd3747,17'd1124,17'd1551,17'd14597,17'd206,17'd8188
},
'{
17'd3,17'd3,17'd1,17'd0,17'd1127,17'd1127,17'd14,17'd1,17'd1,17'd283,17'd283,17'd283,17'd19,17'd19,17'd19,17'd19,17'd0,17'd2,17'd2,17'd2,17'd14,17'd1967,17'd5196,17'd6583,17'd6583,17'd4577,17'd4887,17'd4246,17'd2593,17'd2593,17'd2934,17'd3101,17'd2422,17'd2422,17'd2422,17'd2781,17'd12503,17'd9684,17'd9967,17'd63668,17'd63822,17'd13816,17'd12928,17'd65189,17'd65189,17'd13815,17'd6739,17'd71615,17'd9550,17'd75888,17'd10543,17'd63259,17'd9422,17'd1277,17'd11,17'd25,17'd467,17'd467,17'd1691,17'd1691,17'd23,17'd4,17'd1413,17'd5647,17'd5794,17'd5650,17'd7224,17'd5801,17'd17187,17'd1415,17'd9422,17'd14442,17'd5969,17'd5969,17'd1276,17'd16,17'd3905,17'd18,17'd18,17'd11,17'd20,17'd21,17'd21,17'd21,17'd21,17'd21,17'd285,17'd285,17'd27,17'd27,17'd980,17'd27,17'd19,17'd979,17'd979,17'd287,17'd286,17'd27,17'd28,17'd28,17'd28,17'd287,17'd70879,17'd70879,17'd70879,17'd70879,17'd73110,17'd6902,17'd7061,17'd7555,17'd8047,17'd74462,17'd70288,17'd70288,17'd8047,17'd8047,17'd8047,17'd7557,17'd7557,17'd10408,17'd5657,17'd5805,17'd50679,17'd75889,17'd75890,17'd14602,17'd15747,17'd75891,17'd62580,17'd75892,17'd1006,17'd679,17'd75893,17'd75894,17'd75895,17'd75896,17'd75897,17'd75898,17'd75899,17'd75900,17'd75901,17'd75902,17'd75902,17'd75903,17'd75904,17'd75905,17'd75906,17'd75907,17'd75908,17'd75909,17'd75910,17'd75910,17'd75911,17'd75912,17'd75913,17'd75914,17'd75915,17'd75916,17'd75917,17'd75918,17'd75919,17'd75920,17'd75921,17'd75922,17'd75923,17'd75924,17'd75925,17'd75926,17'd75927,17'd75928,17'd75929,17'd75930,17'd75840,17'd75750,17'd75931,17'd75932,17'd75933,17'd75934,17'd75935,17'd75936,17'd75937,17'd75938,17'd75939,17'd75940,17'd75941,17'd75942,17'd73502,17'd75943,17'd72652,17'd74877,17'd75944,17'd74878,17'd75945,17'd73388,17'd72655,17'd72754,17'd130,17'd132,17'd131,17'd131,17'd132,17'd132,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd134,17'd542,17'd133,17'd3996,17'd13534,17'd75946,17'd75947,17'd75948,17'd75949,17'd75950,17'd75951,17'd75952,17'd75953,17'd62048,17'd21909,17'd75954,17'd75955,17'd75956,17'd18017,17'd18018,17'd18497,17'd16950,17'd75957,17'd75129,17'd75575,17'd75958,17'd75867,17'd16367,17'd75773,17'd9387,17'd9387,17'd10229,17'd11031,17'd12157,17'd12621,17'd75959,17'd12159,17'd11851,17'd11849,17'd6550,17'd6550,17'd6214,17'd28532,17'd75960,17'd28532,17'd5918,17'd6851,17'd10236,17'd10236,17'd9932,17'd9932,17'd11430,17'd11430,17'd11430,17'd11430,17'd10777,17'd10513,17'd8304,17'd8933,17'd8304,17'd9657,17'd9933,17'd9933,17'd27815,17'd27815,17'd10516,17'd10516,17'd10516,17'd10516,17'd10516,17'd10778,17'd10516,17'd10778,17'd10778,17'd11038,17'd11038,17'd31402,17'd31402,17'd31402,17'd11856,17'd31402,17'd31402,17'd68622,17'd68622,17'd74202,17'd69325,17'd72771,17'd68932,17'd68932,17'd75022,17'd75023,17'd75961,17'd75962,17'd75963,17'd75964,17'd72576,17'd69333,17'd75474,17'd75243,17'd75244,17'd75361,17'd75965,17'd75871,17'd75966,17'd75872,17'd75967,17'd75873,17'd75684,17'd75684,17'd75684,17'd75968,17'd75873,17'd75969,17'd74792,17'd75970,17'd75971,17'd75971,17'd75971,17'd75972,17'd75973,17'd75974,17'd68942,17'd69519,17'd75975,17'd66912,17'd65162,17'd69417,17'd67285,17'd65041,17'd63788,17'd65932,17'd17179,17'd75976,17'd67434,17'd75977,17'd48187,17'd12485,17'd5195,17'd4398,17'd629,17'd52462,17'd24496,17'd930,17'd1087,17'd21467,17'd439,17'd586,17'd75792,17'd75978,17'd75979,17'd75980,17'd31904,17'd52107,17'd222,17'd16634,17'd16633,17'd1543,17'd770,17'd1542,17'd1542,17'd281,17'd281,17'd1116,17'd433,17'd1543,17'd250,17'd251,17'd770,17'd1116,17'd29896,17'd30046,17'd75981,17'd75982,17'd964,17'd2588,17'd273,17'd1829,17'd75983,17'd75984,17'd1410,17'd1828,17'd643,17'd426
},
'{
17'd3,17'd3,17'd1,17'd1,17'd14,17'd1127,17'd1127,17'd15,17'd1,17'd1412,17'd283,17'd283,17'd19,17'd19,17'd19,17'd19,17'd0,17'd0,17'd2,17'd2,17'd14,17'd14,17'd6419,17'd5196,17'd5196,17'd7711,17'd7545,17'd4887,17'd2782,17'd2593,17'd2593,17'd2934,17'd2593,17'd2784,17'd3250,17'd1688,17'd1689,17'd64400,17'd64668,17'd9967,17'd13185,17'd63822,17'd74232,17'd71714,17'd67693,17'd65189,17'd13433,17'd13815,17'd63821,17'd13816,17'd6433,17'd10543,17'd14069,17'd9422,17'd19,17'd11,17'd1833,17'd467,17'd467,17'd1691,17'd23,17'd4,17'd9,17'd1413,17'd5647,17'd5514,17'd6277,17'd6108,17'd75491,17'd17187,17'd1414,17'd9422,17'd1276,17'd1276,17'd1276,17'd16,17'd3905,17'd3905,17'd18,17'd18,17'd11,17'd20,17'd21,17'd21,17'd25,17'd25,17'd467,17'd467,17'd286,17'd27,17'd980,17'd980,17'd19,17'd979,17'd979,17'd979,17'd287,17'd286,17'd28,17'd28,17'd28,17'd28,17'd288,17'd70879,17'd70879,17'd70879,17'd18037,17'd18037,17'd6902,17'd7728,17'd8988,17'd8047,17'd8198,17'd8521,17'd70686,17'd8988,17'd7555,17'd50387,17'd21631,17'd7557,17'd75985,17'd12336,17'd5806,17'd13819,17'd53874,17'd75889,17'd75986,17'd75987,17'd75988,17'd75989,17'd75990,17'd75991,17'd75992,17'd75993,17'd75994,17'd75995,17'd75996,17'd75997,17'd75998,17'd75999,17'd76000,17'd76001,17'd76002,17'd76003,17'd76004,17'd76005,17'd76006,17'd76007,17'd76008,17'd76009,17'd76010,17'd76011,17'd76012,17'd76013,17'd76014,17'd76015,17'd76016,17'd76017,17'd76018,17'd76019,17'd76020,17'd76021,17'd76022,17'd76023,17'd76024,17'd76025,17'd76026,17'd76027,17'd76028,17'd76029,17'd76030,17'd76031,17'd76032,17'd75842,17'd76033,17'd76034,17'd75935,17'd75935,17'd76035,17'd76036,17'd76037,17'd76038,17'd76039,17'd76040,17'd76041,17'd73832,17'd76042,17'd73834,17'd75108,17'd73178,17'd73611,17'd76043,17'd71857,17'd71260,17'd72754,17'd1481,17'd132,17'd131,17'd131,17'd131,17'd132,17'd132,17'd130,17'd130,17'd130,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd133,17'd131,17'd132,17'd132,17'd132,17'd134,17'd542,17'd719,17'd7649,17'd6369,17'd76044,17'd76045,17'd76046,17'd30172,17'd76047,17'd76048,17'd75952,17'd76049,17'd21434,17'd62308,17'd76050,17'd76051,17'd75863,17'd76052,17'd18017,17'd17897,17'd18497,17'd16608,17'd75129,17'd75575,17'd75958,17'd75772,17'd76053,17'd19477,17'd9387,17'd9653,17'd10228,17'd11706,17'd76054,17'd12157,17'd75959,17'd12159,17'd11851,17'd11850,17'd6550,17'd6550,17'd6215,17'd6213,17'd75960,17'd75960,17'd6552,17'd6704,17'd8000,17'd8000,17'd9931,17'd9931,17'd69223,17'd69223,17'd11430,17'd11430,17'd10641,17'd10777,17'd9657,17'd8304,17'd8933,17'd8304,17'd27696,17'd27696,17'd27815,17'd27815,17'd10778,17'd10778,17'd10516,17'd10516,17'd10516,17'd10516,17'd10778,17'd10778,17'd10778,17'd11038,17'd11038,17'd31402,17'd31402,17'd31402,17'd31402,17'd76055,17'd76055,17'd76055,17'd68825,17'd72771,17'd69511,17'd69030,17'd68932,17'd75022,17'd76056,17'd74075,17'd73628,17'd74906,17'd75776,17'd69333,17'd74786,17'd75028,17'd75134,17'd76057,17'd75584,17'd76058,17'd76058,17'd76059,17'd75362,17'd75871,17'd75966,17'd75966,17'd76060,17'd76061,17'd76061,17'd75248,17'd75475,17'd76062,17'd74789,17'd74663,17'd76063,17'd76063,17'd76063,17'd76063,17'd67545,17'd76064,17'd76065,17'd66660,17'd66661,17'd65284,17'd76066,17'd76067,17'd63787,17'd65042,17'd65932,17'd17179,17'd65829,17'd67169,17'd65700,17'd76068,17'd5373,17'd64647,17'd2558,17'd3711,17'd52462,17'd35059,17'd930,17'd39034,17'd21467,17'd32405,17'd586,17'd36456,17'd76069,17'd76070,17'd76071,17'd76072,17'd76073,17'd787,17'd16634,17'd1116,17'd16633,17'd1543,17'd17298,17'd75256,17'd15742,17'd29753,17'd29753,17'd787,17'd35208,17'd433,17'd590,17'd250,17'd433,17'd15742,17'd16006,17'd76074,17'd76075,17'd770,17'd8639,17'd607,17'd803,17'd76076,17'd76077,17'd76078,17'd1410,17'd645,17'd970,17'd259
},
'{
17'd283,17'd3,17'd1,17'd1,17'd15,17'd1127,17'd1127,17'd1127,17'd0,17'd1,17'd283,17'd283,17'd19,17'd19,17'd19,17'd979,17'd1277,17'd16,17'd2,17'd2,17'd0,17'd0,17'd2,17'd1127,17'd4885,17'd5196,17'd7545,17'd7545,17'd2784,17'd2784,17'd2593,17'd2593,17'd3751,17'd2782,17'd3250,17'd4247,17'd2595,17'd14,17'd12929,17'd9684,17'd13065,17'd69723,17'd75888,17'd10264,17'd73646,17'd73541,17'd69723,17'd13184,17'd13433,17'd13433,17'd63821,17'd6433,17'd73990,17'd67452,17'd75491,17'd19,17'd286,17'd467,17'd467,17'd467,17'd25,17'd25,17'd9,17'd9,17'd4,17'd5647,17'd5651,17'd6108,17'd75490,17'd1277,17'd1414,17'd17187,17'd16,17'd1277,17'd1276,17'd16,17'd17,17'd17,17'd16,17'd18,17'd806,17'd8814,17'd2933,17'd2591,17'd25,17'd25,17'd467,17'd467,17'd285,17'd26,17'd1128,17'd1128,17'd18,17'd19,17'd1,17'd19,17'd287,17'd287,17'd287,17'd28,17'd652,17'd652,17'd29,17'd288,17'd2118,17'd2118,17'd3907,17'd4431,17'd18037,17'd6744,17'd7061,17'd7728,17'd8988,17'd8197,17'd8197,17'd8827,17'd2937,17'd7555,17'd7555,17'd7556,17'd9555,17'd70077,17'd11737,17'd13068,17'd13187,17'd76079,17'd76080,17'd76081,17'd76082,17'd75384,17'd76083,17'd76084,17'd76085,17'd76086,17'd76087,17'd76088,17'd76089,17'd76090,17'd317,17'd76091,17'd76092,17'd76093,17'd76094,17'd76095,17'd76096,17'd76097,17'd76098,17'd76099,17'd76100,17'd76101,17'd76102,17'd76103,17'd76104,17'd76105,17'd76106,17'd76107,17'd76108,17'd76017,17'd76109,17'd76110,17'd76111,17'd76112,17'd76113,17'd76114,17'd76115,17'd76116,17'd76117,17'd76117,17'd76118,17'd76119,17'd76120,17'd76121,17'd75843,17'd75934,17'd76122,17'd76123,17'd76124,17'd76125,17'd76126,17'd76127,17'd76128,17'd76129,17'd76130,17'd75102,17'd75219,17'd74402,17'd76131,17'd75108,17'd73611,17'd73078,17'd70742,17'd355,17'd127,17'd356,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd542,17'd719,17'd132,17'd2862,17'd17140,17'd76132,17'd76133,17'd76134,17'd76135,17'd76136,17'd76137,17'd35747,17'd39608,17'd61923,17'd76138,17'd10199,17'd17033,17'd16482,17'd16949,17'd76139,17'd76140,17'd74894,17'd74768,17'd75129,17'd76141,17'd75772,17'd76142,17'd17278,17'd9386,17'd10895,17'd10895,17'd9389,17'd76054,17'd76054,17'd12159,17'd12158,17'd12003,17'd11850,17'd6216,17'd6216,17'd6215,17'd6213,17'd28532,17'd28532,17'd5761,17'd5761,17'd7999,17'd8000,17'd8629,17'd9931,17'd9931,17'd9932,17'd69223,17'd11430,17'd10777,17'd10777,17'd10777,17'd10513,17'd8304,17'd8304,17'd29740,17'd27696,17'd9933,17'd27815,17'd10778,17'd11038,17'd68510,17'd68928,17'd68928,17'd69692,17'd29592,17'd29592,17'd29592,17'd27933,17'd68928,17'd10778,17'd11038,17'd68510,17'd68624,17'd68725,17'd68933,17'd76143,17'd69229,17'd76144,17'd76145,17'd69134,17'd75774,17'd75775,17'd74905,17'd76146,17'd75776,17'd74908,17'd71178,17'd76147,17'd75135,17'd75682,17'd75584,17'd76148,17'd76148,17'd76149,17'd76149,17'd76148,17'd76059,17'd75965,17'd75871,17'd75871,17'd75871,17'd75475,17'd76062,17'd74790,17'd75029,17'd76150,17'd76151,17'd71887,17'd68941,17'd68941,17'd67658,17'd76152,17'd67030,17'd66422,17'd76153,17'd70854,17'd74329,17'd71795,17'd26955,17'd15732,17'd63357,17'd14975,17'd65705,17'd65829,17'd67169,17'd76068,17'd16623,17'd4867,17'd4558,17'd18035,17'd3874,17'd18144,17'd35059,17'd53745,17'd59123,17'd21467,17'd32405,17'd75253,17'd36324,17'd75886,17'd76154,17'd33377,17'd76155,17'd76156,17'd221,17'd767,17'd75256,17'd1116,17'd16633,17'd16633,17'd15742,17'd16746,17'd29896,17'd16263,17'd76157,17'd787,17'd1116,17'd589,17'd401,17'd589,17'd281,17'd29753,17'd16140,17'd16264,17'd15742,17'd647,17'd783,17'd260,17'd1828,17'd76158,17'd76159,17'd76159,17'd76160,17'd411,17'd1823,17'd1263
},
'{
17'd283,17'd3,17'd3,17'd1,17'd1830,17'd1127,17'd4247,17'd1127,17'd15,17'd1,17'd283,17'd283,17'd19,17'd19,17'd19,17'd979,17'd1277,17'd16,17'd2,17'd2,17'd0,17'd0,17'd2,17'd466,17'd4885,17'd6419,17'd7214,17'd7545,17'd3250,17'd2592,17'd2784,17'd2593,17'd3751,17'd2593,17'd2422,17'd4247,17'd2595,17'd466,17'd1967,17'd9815,17'd10801,17'd73541,17'd67817,17'd76161,17'd10088,17'd76162,17'd13065,17'd13185,17'd13184,17'd63821,17'd63821,17'd9550,17'd6268,17'd6267,17'd67452,17'd9422,17'd5969,17'd2424,17'd1833,17'd467,17'd21,17'd25,17'd25,17'd4,17'd4,17'd23,17'd5647,17'd5651,17'd3748,17'd1276,17'd1277,17'd22965,17'd17,17'd1277,17'd1276,17'd16,17'd17,17'd17,17'd16,17'd18,17'd2423,17'd806,17'd1275,17'd2591,17'd25,17'd25,17'd467,17'd467,17'd285,17'd26,17'd1128,17'd20404,17'd18,17'd16,17'd0,17'd16,17'd287,17'd287,17'd2424,17'd287,17'd652,17'd653,17'd289,17'd29,17'd981,17'd981,17'd3907,17'd3907,17'd3907,17'd288,17'd28,17'd6902,17'd6902,17'd7728,17'd8827,17'd76163,17'd8827,17'd2937,17'd7555,17'd7728,17'd7225,17'd7556,17'd70077,17'd75047,17'd76164,17'd3106,17'd3106,17'd76165,17'd76166,17'd75890,17'd76167,17'd76168,17'd76169,17'd76170,17'd59912,17'd76171,17'd76172,17'd76173,17'd76174,17'd76175,17'd76176,17'd76177,17'd76178,17'd76179,17'd76180,17'd76180,17'd76181,17'd76182,17'd76183,17'd76184,17'd76185,17'd76186,17'd76187,17'd76188,17'd76189,17'd76190,17'd76191,17'd76192,17'd76110,17'd76193,17'd76194,17'd76195,17'd76196,17'd76197,17'd76198,17'd76199,17'd76200,17'd76201,17'd76200,17'd76202,17'd76203,17'd75933,17'd76204,17'd76204,17'd76123,17'd76205,17'd76206,17'd76207,17'd75938,17'd75939,17'd76129,17'd76130,17'd75102,17'd75219,17'd73606,17'd75853,17'd75108,17'd76208,17'd70831,17'd73283,17'd1479,17'd1481,17'd133,17'd133,17'd133,17'd133,17'd134,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd133,17'd131,17'd132,17'd132,17'd132,17'd132,17'd542,17'd1197,17'd132,17'd5311,17'd4654,17'd18931,17'd76209,17'd76210,17'd76211,17'd76212,17'd76213,17'd76214,17'd39608,17'd76215,17'd76216,17'd22244,17'd76217,17'd17150,17'd16098,17'd18253,17'd18018,17'd76140,17'd18618,17'd75957,17'd75867,17'd76141,17'd76218,17'd76053,17'd75773,17'd9388,17'd9519,17'd9519,17'd12300,17'd76219,17'd12003,17'd12158,17'd12302,17'd11851,17'd6850,17'd6216,17'd6214,17'd6213,17'd6214,17'd6213,17'd27930,17'd5613,17'd6704,17'd7999,17'd8000,17'd8629,17'd9931,17'd9931,17'd69223,17'd69223,17'd9657,17'd10777,17'd10641,17'd10777,17'd9657,17'd8304,17'd29740,17'd29740,17'd27696,17'd9933,17'd10778,17'd11038,17'd68622,17'd68624,17'd68624,17'd68510,17'd72566,17'd72566,17'd68928,17'd68928,17'd68623,17'd68623,17'd68624,17'd68724,17'd68726,17'd68935,17'd69229,17'd69134,17'd76220,17'd76221,17'd76222,17'd76223,17'd69232,17'd75132,17'd75025,17'd72674,17'd74908,17'd71178,17'd76147,17'd76224,17'd75584,17'd75360,17'd76148,17'd76148,17'd76149,17'd76149,17'd76149,17'd76149,17'd76058,17'd76059,17'd75361,17'd76059,17'd76058,17'd75360,17'd75682,17'd76225,17'd76226,17'd76227,17'd76227,17'd76227,17'd70958,17'd76228,17'd76229,17'd70369,17'd70660,17'd74555,17'd76230,17'd76231,17'd71889,17'd26955,17'd15229,17'd15100,17'd65288,17'd14857,17'd67557,17'd68410,17'd75484,17'd14736,17'd4867,17'd5938,17'd5936,17'd5628,17'd8314,17'd36748,17'd53745,17'd1524,17'd76232,17'd51582,17'd28313,17'd76233,17'd76234,17'd75979,17'd76154,17'd34511,17'd76235,17'd76236,17'd76237,17'd787,17'd15742,17'd20001,17'd20001,17'd20001,17'd16746,17'd215,17'd30046,17'd587,17'd76238,17'd619,17'd787,17'd20001,17'd17423,17'd17423,17'd18516,17'd215,17'd76239,17'd29896,17'd76240,17'd2109,17'd17787,17'd260,17'd1828,17'd76160,17'd76160,17'd76158,17'd971,17'd411,17'd1667,17'd1396
},
'{
17'd20,17'd10,17'd979,17'd1277,17'd1830,17'd3249,17'd1967,17'd2594,17'd1127,17'd0,17'd283,17'd283,17'd3,17'd283,17'd1412,17'd1,17'd283,17'd3,17'd12,17'd12,17'd12,17'd12,17'd2,17'd466,17'd2,17'd14,17'd1127,17'd1688,17'd1688,17'd3250,17'd3250,17'd3252,17'd2593,17'd2593,17'd2784,17'd2422,17'd1688,17'd1127,17'd14,17'd1967,17'd63260,17'd63258,17'd6274,17'd10543,17'd74342,17'd10264,17'd63822,17'd70278,17'd73541,17'd75888,17'd9550,17'd74232,17'd63821,17'd9550,17'd10264,17'd9552,17'd63117,17'd1276,17'd979,17'd25,17'd467,17'd1691,17'd1691,17'd1690,17'd5,17'd5,17'd5,17'd8,17'd8827,17'd4429,17'd19,17'd1416,17'd1416,17'd17,17'd16,17'd16,17'd2,17'd2,17'd2,17'd2,17'd18,17'd11,17'd11,17'd10,17'd21,17'd25,17'd9,17'd9,17'd9,17'd20,17'd20404,17'd1128,17'd19,17'd16,17'd17,17'd17,17'd28,17'd28,17'd286,17'd286,17'd28,17'd652,17'd289,17'd809,17'd288,17'd29,17'd30,17'd30,17'd654,17'd3102,17'd2118,17'd70879,17'd73110,17'd9275,17'd8988,17'd8197,17'd8197,17'd8047,17'd8047,17'd8047,17'd7386,17'd7556,17'd9555,17'd11211,17'd12336,17'd73543,17'd12506,17'd3259,17'd14748,17'd47968,17'd1971,17'd15121,17'd76241,17'd1132,17'd60891,17'd76242,17'd76243,17'd76244,17'd76245,17'd76246,17'd84,17'd76247,17'd76248,17'd76249,17'd76250,17'd76251,17'd76252,17'd76253,17'd76254,17'd76255,17'd76256,17'd76257,17'd76258,17'd76259,17'd76260,17'd76261,17'd76262,17'd76263,17'd76264,17'd76194,17'd76265,17'd76266,17'd76267,17'd76268,17'd76269,17'd76270,17'd76270,17'd76270,17'd76270,17'd76271,17'd76272,17'd76273,17'd76204,17'd75935,17'd76035,17'd76274,17'd76275,17'd75847,17'd76276,17'd76277,17'd75940,17'd74992,17'd74054,17'd73391,17'd73835,17'd75108,17'd76278,17'd70537,17'd70217,17'd4163,17'd356,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd1197,17'd134,17'd135,17'd10492,17'd6056,17'd5746,17'd76279,17'd76280,17'd76281,17'd76282,17'd76283,17'd76284,17'd21431,17'd76285,17'd76286,17'd55250,17'd16817,17'd76287,17'd76288,17'd18849,17'd18253,17'd76140,17'd76140,17'd16608,17'd18370,17'd75958,17'd76218,17'd17059,17'd15721,17'd9651,17'd75959,17'd75959,17'd12158,17'd12003,17'd12158,17'd12158,17'd12301,17'd11851,17'd68172,17'd68172,17'd7667,17'd8931,17'd6213,17'd28532,17'd50670,17'd76289,17'd76289,17'd6552,17'd6387,17'd6852,17'd10236,17'd8000,17'd9931,17'd69223,17'd76290,17'd76291,17'd11430,17'd11430,17'd10777,17'd10513,17'd9657,17'd8304,17'd9091,17'd7668,17'd10516,17'd12471,17'd12763,17'd76292,17'd76293,17'd76293,17'd76294,17'd76295,17'd68726,17'd68726,17'd68728,17'd68826,17'd68826,17'd68935,17'd75023,17'd75023,17'd69230,17'd76296,17'd76221,17'd69415,17'd76297,17'd69699,17'd69882,17'd70056,17'd69700,17'd69608,17'd71283,17'd75134,17'd75243,17'd75682,17'd75584,17'd75584,17'd75584,17'd75584,17'd75584,17'd76298,17'd76298,17'd75584,17'd76299,17'd76300,17'd76299,17'd76301,17'd71178,17'd69975,17'd74785,17'd76302,17'd72466,17'd72466,17'd76302,17'd76303,17'd76229,17'd76229,17'd76304,17'd76305,17'd66302,17'd66303,17'd66060,17'd76306,17'd14306,17'd19093,17'd18379,17'd15101,17'd17178,17'd65705,17'd15103,17'd68410,17'd14736,17'd5373,17'd50843,17'd2391,17'd69614,17'd5934,17'd6720,17'd56884,17'd1524,17'd59123,17'd1377,17'd28313,17'd76307,17'd34511,17'd36908,17'd37575,17'd76308,17'd37044,17'd76309,17'd76237,17'd76310,17'd75694,17'd75694,17'd15742,17'd15742,17'd20266,17'd435,17'd75039,17'd39035,17'd30046,17'd587,17'd619,17'd76310,17'd787,17'd15742,17'd281,17'd74929,17'd76311,17'd76312,17'd15355,17'd22267,17'd966,17'd2778,17'd260,17'd803,17'd1410,17'd1098,17'd1098,17'd1272,17'd424,17'd604,17'd604
},
'{
17'd2598,17'd11,17'd19,17'd1277,17'd1830,17'd63116,17'd1967,17'd1688,17'd1127,17'd15,17'd1412,17'd283,17'd283,17'd283,17'd1412,17'd1,17'd283,17'd3,17'd3,17'd12,17'd12,17'd12,17'd0,17'd2,17'd2,17'd0,17'd14,17'd1127,17'd1688,17'd1688,17'd1688,17'd2422,17'd2784,17'd2784,17'd2784,17'd2422,17'd1688,17'd1689,17'd14,17'd14,17'd63116,17'd14069,17'd74233,17'd63521,17'd76313,17'd76162,17'd13185,17'd13185,17'd74234,17'd67694,17'd73646,17'd74232,17'd13184,17'd63821,17'd13816,17'd75888,17'd74233,17'd68083,17'd5969,17'd10,17'd467,17'd1691,17'd21631,17'd7384,17'd5,17'd3594,17'd5,17'd5,17'd1690,17'd467,17'd10,17'd18,17'd1416,17'd17,17'd17,17'd16,17'd0,17'd2,17'd2,17'd466,17'd16,17'd18,17'd18,17'd19,17'd10,17'd25,17'd25,17'd9,17'd25,17'd21,17'd11,17'd3905,17'd16,17'd16,17'd14442,17'd16,17'd653,17'd652,17'd28,17'd287,17'd287,17'd28,17'd29,17'd30,17'd809,17'd809,17'd3102,17'd654,17'd2597,17'd2597,17'd2936,17'd17187,17'd76314,17'd73110,17'd6902,17'd7728,17'd8197,17'd8521,17'd74462,17'd52025,17'd7388,17'd7556,17'd9555,17'd75985,17'd72282,17'd76315,17'd9816,17'd11208,17'd12333,17'd12785,17'd1968,17'd1694,17'd15363,17'd475,17'd987,17'd60891,17'd76316,17'd63982,17'd76317,17'd76318,17'd76319,17'd76320,17'd76321,17'd76322,17'd76323,17'd76324,17'd76325,17'd76325,17'd76326,17'd76327,17'd76328,17'd76329,17'd76330,17'd76331,17'd76332,17'd76333,17'd76334,17'd76335,17'd76336,17'd76195,17'd76337,17'd76338,17'd76338,17'd76339,17'd76340,17'd76341,17'd76342,17'd76343,17'd76344,17'd76272,17'd76344,17'd76345,17'd76204,17'd76346,17'd76274,17'd75660,17'd76347,17'd76348,17'd76349,17'd76350,17'd76351,17'd76352,17'd76353,17'd74876,17'd73178,17'd76278,17'd70537,17'd127,17'd356,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd134,17'd132,17'd131,17'd2861,17'd76354,17'd76355,17'd76356,17'd76357,17'd76358,17'd76359,17'd76360,17'd76361,17'd76362,17'd75565,17'd76363,17'd76364,17'd76365,17'd76366,17'd76367,17'd76288,17'd76368,17'd76139,17'd76369,17'd76140,17'd76370,17'd76141,17'd76371,17'd17170,17'd76372,17'd9518,17'd76373,17'd75577,17'd12158,17'd12302,17'd12003,17'd12003,17'd71963,17'd12301,17'd11849,17'd11849,17'd7176,17'd7667,17'd6214,17'd6213,17'd50670,17'd50670,17'd27695,17'd50670,17'd5332,17'd6388,17'd7999,17'd7999,17'd8629,17'd9931,17'd69223,17'd76291,17'd11430,17'd11430,17'd10777,17'd10777,17'd10513,17'd10513,17'd10513,17'd7668,17'd10380,17'd10517,17'd10779,17'd29162,17'd76293,17'd68627,17'd68627,17'd68627,17'd76374,17'd76374,17'd76375,17'd68730,17'd75775,17'd68937,17'd74075,17'd76376,17'd69032,17'd75580,17'd76377,17'd75242,17'd75242,17'd69792,17'd70159,17'd70658,17'd71283,17'd71283,17'd71283,17'd76378,17'd76057,17'd76057,17'd76298,17'd75584,17'd75584,17'd75584,17'd75584,17'd75584,17'd75584,17'd75584,17'd76379,17'd76224,17'd76147,17'd72069,17'd76380,17'd69138,17'd76381,17'd76382,17'd76382,17'd76383,17'd76383,17'd76384,17'd76385,17'd70465,17'd76386,17'd76305,17'd66176,17'd70370,17'd65035,17'd16253,17'd14306,17'd15100,17'd63946,17'd17414,17'd76387,17'd62447,17'd63653,17'd13572,17'd12636,17'd4558,17'd4398,17'd5935,17'd61543,17'd37956,17'd53593,17'd76388,17'd52105,17'd76389,17'd19492,17'd761,17'd76390,17'd76391,17'd36457,17'd76391,17'd76308,17'd585,17'd52197,17'd20266,17'd29753,17'd29173,17'd75694,17'd76310,17'd76157,17'd39035,17'd16005,17'd16005,17'd177,17'd30046,17'd76157,17'd76157,17'd76157,17'd619,17'd76157,17'd29442,17'd76392,17'd19363,17'd15626,17'd461,17'd460,17'd801,17'd646,17'd641,17'd644,17'd803,17'd1685,17'd1272,17'd1272,17'd424,17'd1272,17'd1272
},
'{
17'd20404,17'd1128,17'd3,17'd1,17'd1830,17'd1830,17'd15,17'd1127,17'd4247,17'd14,17'd1,17'd1,17'd1412,17'd1412,17'd283,17'd3,17'd3,17'd3,17'd283,17'd3,17'd3,17'd12,17'd0,17'd1,17'd0,17'd0,17'd15,17'd1127,17'd4247,17'd4247,17'd1689,17'd1689,17'd2422,17'd2422,17'd2422,17'd1831,17'd1831,17'd1688,17'd1127,17'd14,17'd15,17'd1830,17'd14069,17'd74233,17'd63521,17'd10543,17'd76313,17'd75888,17'd73541,17'd74107,17'd71197,17'd13185,17'd13816,17'd74232,17'd74232,17'd10402,17'd10662,17'd63521,17'd76393,17'd75491,17'd1833,17'd285,17'd1832,17'd7384,17'd5,17'd5,17'd5,17'd5,17'd4,17'd25,17'd808,17'd10,17'd3905,17'd4089,17'd17,17'd17,17'd0,17'd0,17'd14,17'd466,17'd17,17'd17,17'd18,17'd18,17'd11,17'd10,17'd25,17'd25,17'd9,17'd1413,17'd808,17'd20404,17'd4089,17'd17,17'd16,17'd16,17'd4089,17'd3905,17'd16,17'd1276,17'd287,17'd287,17'd652,17'd809,17'd1693,17'd11207,17'd76394,17'd655,17'd2597,17'd2258,17'd2258,17'd2597,17'd76395,17'd981,17'd28,17'd286,17'd8047,17'd74462,17'd74462,17'd52025,17'd8047,17'd8047,17'd9276,17'd9555,17'd75985,17'd72282,17'd10269,17'd11210,17'd11208,17'd2430,17'd1968,17'd1694,17'd76241,17'd76396,17'd59497,17'd65585,17'd63823,17'd76171,17'd76397,17'd76398,17'd76399,17'd76319,17'd76319,17'd76400,17'd76401,17'd76402,17'd76403,17'd76404,17'd76405,17'd76330,17'd76406,17'd76407,17'd76408,17'd76409,17'd76410,17'd76411,17'd76412,17'd76413,17'd76414,17'd76415,17'd76416,17'd76417,17'd76417,17'd76418,17'd76419,17'd76420,17'd76421,17'd76422,17'd76423,17'd76424,17'd76425,17'd76426,17'd76427,17'd76428,17'd75846,17'd76429,17'd75939,17'd76349,17'd75940,17'd76351,17'd75219,17'd73606,17'd76131,17'd73929,17'd73292,17'd71954,17'd72754,17'd20762,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd134,17'd132,17'd132,17'd3168,17'd18578,17'd4654,17'd19047,17'd76430,17'd76431,17'd76432,17'd76433,17'd76434,17'd76435,17'd76436,17'd34493,17'd76437,17'd76438,17'd13021,17'd76439,17'd76440,17'd17774,17'd18253,17'd76140,17'd18497,17'd16608,17'd76370,17'd76441,17'd76441,17'd76053,17'd75773,17'd20112,17'd76442,17'd76443,17'd76444,17'd11849,17'd11849,17'd71963,17'd71963,17'd11850,17'd11850,17'd6850,17'd7176,17'd6215,17'd6214,17'd5915,17'd5915,17'd27695,17'd76289,17'd5613,17'd5761,17'd6552,17'd6704,17'd8000,17'd9931,17'd76290,17'd76290,17'd69223,17'd11430,17'd11430,17'd11430,17'd69223,17'd10513,17'd10777,17'd8780,17'd9934,17'd11039,17'd8001,17'd7012,17'd76445,17'd68512,17'd68628,17'd76446,17'd76447,17'd76448,17'd73960,17'd76449,17'd76450,17'd76451,17'd76452,17'd76452,17'd75025,17'd75583,17'd72674,17'd75026,17'd76453,17'd76454,17'd71178,17'd71178,17'd71178,17'd76301,17'd76301,17'd76455,17'd76456,17'd76456,17'd76457,17'd76456,17'd76456,17'd76456,17'd76301,17'd76147,17'd76147,17'd76458,17'd76459,17'd76460,17'd69975,17'd74785,17'd74784,17'd76461,17'd68732,17'd68732,17'd68732,17'd68051,17'd67657,17'd76462,17'd76463,17'd76463,17'd66783,17'd76464,17'd76465,17'd76466,17'd72578,17'd76467,17'd14056,17'd18748,17'd18030,17'd65690,17'd62702,17'd65947,17'd13689,17'd12483,17'd11049,17'd2558,17'd629,17'd9247,17'd33999,17'd58129,17'd76468,17'd52105,17'd76389,17'd52197,17'd76233,17'd76469,17'd37575,17'd36604,17'd36325,17'd76071,17'd76470,17'd52023,17'd439,17'd29753,17'd32724,17'd790,17'd767,17'd76471,17'd39330,17'd398,17'd30945,17'd32883,17'd618,17'd75253,17'd16263,17'd16263,17'd76157,17'd76157,17'd75599,17'd76472,17'd76473,17'd179,17'd22267,17'd76474,17'd460,17'd263,17'd1268,17'd273,17'd643,17'd803,17'd971,17'd1685,17'd424,17'd424,17'd1272,17'd1272
},
'{
17'd3905,17'd18,17'd12,17'd12,17'd1,17'd1830,17'd15,17'd14,17'd4247,17'd1127,17'd14,17'd0,17'd1412,17'd1412,17'd283,17'd3,17'd3,17'd3,17'd283,17'd3,17'd12,17'd12,17'd1,17'd1412,17'd0,17'd0,17'd1830,17'd14,17'd4247,17'd4247,17'd1689,17'd1967,17'd1689,17'd1688,17'd1831,17'd1831,17'd1831,17'd1688,17'd1127,17'd14,17'd1830,17'd15,17'd1830,17'd63117,17'd67452,17'd14187,17'd73768,17'd74342,17'd75888,17'd76162,17'd71197,17'd71709,17'd73541,17'd10264,17'd10402,17'd75888,17'd6103,17'd6267,17'd5967,17'd9274,17'd5515,17'd286,17'd1832,17'd7383,17'd24,17'd24,17'd5,17'd5,17'd4,17'd4,17'd9,17'd16389,17'd1128,17'd3905,17'd4089,17'd1416,17'd2,17'd15,17'd14,17'd1127,17'd1415,17'd17,17'd17,17'd18,17'd19,17'd11,17'd10,17'd25,17'd25,17'd1413,17'd16389,17'd11,17'd4089,17'd1416,17'd17,17'd17,17'd3905,17'd17,17'd17187,17'd16,17'd287,17'd287,17'd28,17'd288,17'd76394,17'd11207,17'd470,17'd470,17'd3752,17'd3429,17'd52621,17'd12195,17'd982,17'd31,17'd2118,17'd287,17'd286,17'd7385,17'd52025,17'd8197,17'd8197,17'd8988,17'd9276,17'd9555,17'd9555,17'd6903,17'd6903,17'd6598,17'd3907,17'd3431,17'd2260,17'd1553,17'd296,17'd816,17'd60519,17'd63823,17'd76475,17'd76476,17'd76477,17'd76400,17'd76478,17'd76479,17'd76480,17'd76480,17'd76481,17'd76482,17'd76483,17'd76484,17'd76485,17'd76486,17'd76408,17'd76487,17'd76488,17'd76489,17'd76490,17'd76338,17'd76338,17'd76491,17'd76339,17'd76339,17'd76492,17'd76492,17'd76492,17'd76493,17'd76494,17'd76424,17'd75752,17'd76495,17'd76496,17'd75844,17'd76497,17'd76498,17'd76499,17'd76500,17'd76429,17'd76501,17'd76039,17'd76502,17'd75941,17'd75664,17'd73607,17'd73835,17'd74050,17'd73292,17'd72655,17'd72754,17'd20762,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd1197,17'd134,17'd132,17'd131,17'd3168,17'd4336,17'd76503,17'd18818,17'd76504,17'd30022,17'd31235,17'd76505,17'd32866,17'd17621,17'd76506,17'd37545,17'd76507,17'd76508,17'd12883,17'd76509,17'd76510,17'd16605,17'd17404,17'd16607,17'd16607,17'd74894,17'd18618,17'd17899,17'd76441,17'd76511,17'd19477,17'd76512,17'd76513,17'd76514,17'd76443,17'd11851,17'd11849,17'd68926,17'd68926,17'd11850,17'd11850,17'd6850,17'd7176,17'd6215,17'd6214,17'd5916,17'd5916,17'd50670,17'd76289,17'd52268,17'd5613,17'd5761,17'd5918,17'd7999,17'd8000,17'd8629,17'd76515,17'd76290,17'd76290,17'd69223,17'd69223,17'd69223,17'd69223,17'd10513,17'd10513,17'd27696,17'd9934,17'd10380,17'd10517,17'd68625,17'd68626,17'd68514,17'd76516,17'd74775,17'd76517,17'd76518,17'd74076,17'd73743,17'd73743,17'd76146,17'd76519,17'd76520,17'd75776,17'd74908,17'd72069,17'd75027,17'd71178,17'd71178,17'd76147,17'd76147,17'd76301,17'd76455,17'd76455,17'd76301,17'd76147,17'd76301,17'd76147,17'd76458,17'd74909,17'd74909,17'd71060,17'd71060,17'd76521,17'd70160,17'd76302,17'd68940,17'd76522,17'd68732,17'd68404,17'd68404,17'd68404,17'd68404,17'd67911,17'd76523,17'd76524,17'd76525,17'd65925,17'd67029,17'd76526,17'd65160,17'd76527,17'd76528,17'd13684,17'd17290,17'd19229,17'd76529,17'd76530,17'd14175,17'd14176,17'd60399,17'd4557,17'd4398,17'd9403,17'd9247,17'd76531,17'd39030,17'd52534,17'd52196,17'd76389,17'd766,17'd52023,17'd76469,17'd75980,17'd37045,17'd36604,17'd34003,17'd34667,17'd76469,17'd220,17'd76310,17'd615,17'd32724,17'd790,17'd787,17'd219,17'd32408,17'd76532,17'd176,17'd32085,17'd618,17'd19240,17'd39035,17'd615,17'd76157,17'd16263,17'd75379,17'd76533,17'd74801,17'd252,17'd805,17'd456,17'd265,17'd257,17'd272,17'd272,17'd644,17'd803,17'd971,17'd971,17'd424,17'd424,17'd424,17'd424
},
'{
17'd2,17'd0,17'd12,17'd12,17'd3,17'd1,17'd1,17'd14,17'd1127,17'd1688,17'd1689,17'd15,17'd1,17'd1412,17'd283,17'd1275,17'd12,17'd3,17'd3,17'd3,17'd12,17'd12,17'd3,17'd283,17'd0,17'd0,17'd1,17'd0,17'd1127,17'd4247,17'd1127,17'd14,17'd14,17'd1127,17'd4247,17'd2594,17'd2594,17'd4247,17'd1127,17'd14,17'd16,17'd16,17'd16,17'd14442,17'd14988,17'd67695,17'd5963,17'd67577,17'd6433,17'd64667,17'd14441,17'd70076,17'd63387,17'd10543,17'd6267,17'd6267,17'd63520,17'd10662,17'd76534,17'd76535,17'd75262,17'd75696,17'd2937,17'd1690,17'd284,17'd24,17'd5,17'd6,17'd5,17'd4,17'd4,17'd9,17'd21,17'd1128,17'd4089,17'd22965,17'd466,17'd14,17'd15,17'd14,17'd14,17'd2,17'd2,17'd12,17'd18,17'd11,17'd10,17'd10,17'd10,17'd10,17'd808,17'd808,17'd19,17'd4089,17'd1416,17'd17,17'd14442,17'd9969,17'd1415,17'd17,17'd18,17'd19,17'd287,17'd76536,17'd2118,17'd654,17'd469,17'd292,17'd293,17'd293,17'd11071,17'd10925,17'd10925,17'd3593,17'd10092,17'd2118,17'd28,17'd27,17'd285,17'd2937,17'd8047,17'd8988,17'd8988,17'd7728,17'd7556,17'd7225,17'd7225,17'd7225,17'd9555,17'd10093,17'd11208,17'd2939,17'd39,17'd76537,17'd76538,17'd76172,17'd76539,17'd76540,17'd76541,17'd76542,17'd76543,17'd76544,17'd76545,17'd76546,17'd76547,17'd76548,17'd76549,17'd76332,17'd76333,17'd76334,17'd76550,17'd76551,17'd76552,17'd76553,17'd76554,17'd76555,17'd76555,17'd76556,17'd76557,17'd76558,17'd76559,17'd76494,17'd76560,17'd76271,17'd76561,17'd76562,17'd75937,17'd76563,17'd76563,17'd76564,17'd76565,17'd76566,17'd76500,17'd75660,17'd76567,17'd76568,17'd76040,17'd76569,17'd74054,17'd76570,17'd73600,17'd72986,17'd76043,17'd71477,17'd20762,17'd1481,17'd130,17'd132,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd1197,17'd134,17'd132,17'd132,17'd3168,17'd76571,17'd13534,17'd76572,17'd76573,17'd76574,17'd76575,17'd76576,17'd76577,17'd76578,17'd76579,17'd76580,17'd34326,17'd76581,17'd76582,17'd45901,17'd76583,17'd75863,17'd17774,17'd16244,17'd16117,17'd16367,17'd16486,17'd76053,17'd17776,17'd76511,17'd16367,17'd19982,17'd21613,17'd76442,17'd76442,17'd75959,17'd12302,17'd76584,17'd76584,17'd68621,17'd10379,17'd7176,17'd7176,17'd7667,17'd7667,17'd6552,17'd6552,17'd5915,17'd50670,17'd52268,17'd52268,17'd27930,17'd5761,17'd6552,17'd9523,17'd8629,17'd8629,17'd9931,17'd9931,17'd9932,17'd9932,17'd9932,17'd9931,17'd69223,17'd10513,17'd10513,17'd8780,17'd9933,17'd10380,17'd10380,17'd10517,17'd68626,17'd29300,17'd76585,17'd76585,17'd76516,17'd76517,17'd76586,17'd76518,17'd76587,17'd76587,17'd76588,17'd76381,17'd68940,17'd74785,17'd74785,17'd69975,17'd76589,17'd76460,17'd76589,17'd76589,17'd76590,17'd76591,17'd76459,17'd76460,17'd76460,17'd69975,17'd70160,17'd74785,17'd76302,17'd68940,17'd76383,17'd76383,17'd68051,17'd68732,17'd67911,17'd76592,17'd76593,17'd76593,17'd76593,17'd76593,17'd76593,17'd76594,17'd67543,17'd76595,17'd65925,17'd76596,17'd65680,17'd13927,17'd76597,17'd76598,17'd73528,17'd76599,17'd76600,17'd13568,17'd73422,17'd67173,17'd67292,17'd76601,17'd4711,17'd5936,17'd8314,17'd9102,17'd24496,17'd52195,17'd20711,17'd18759,17'd76602,17'd19602,17'd38073,17'd31904,17'd35062,17'd37575,17'd396,17'd36325,17'd35209,17'd35909,17'd76603,17'd220,17'd16263,17'd29753,17'd18633,17'd36907,17'd76604,17'd36324,17'd33540,17'd76605,17'd76606,17'd76607,17'd76233,17'd35617,17'd177,17'd30046,17'd39628,17'd76608,17'd76609,17'd76610,17'd76611,17'd279,17'd278,17'd278,17'd1274,17'd263,17'd1407,17'd270,17'd1828,17'd1828,17'd971,17'd1685,17'd971,17'd971,17'd971,17'd971
},
'{
17'd1689,17'd14,17'd0,17'd12,17'd3,17'd283,17'd1,17'd0,17'd14,17'd1688,17'd1688,17'd1967,17'd15,17'd1,17'd283,17'd1275,17'd3,17'd3,17'd3,17'd3,17'd12,17'd12,17'd3,17'd3,17'd0,17'd0,17'd1,17'd1,17'd15,17'd1127,17'd1127,17'd14,17'd15,17'd14,17'd1127,17'd4247,17'd4247,17'd4247,17'd1127,17'd14,17'd17,17'd1277,17'd1276,17'd16,17'd0,17'd4732,17'd13814,17'd75159,17'd10543,17'd64930,17'd63520,17'd10662,17'd63521,17'd63258,17'd63387,17'd6267,17'd64930,17'd64930,17'd10090,17'd76612,17'd5968,17'd6276,17'd8827,17'd1691,17'd23,17'd24,17'd5,17'd6,17'd6,17'd6,17'd4,17'd4,17'd9,17'd21,17'd20404,17'd4089,17'd466,17'd1127,17'd1967,17'd1967,17'd14,17'd14,17'd2,17'd0,17'd16,17'd19,17'd979,17'd10,17'd808,17'd10,17'd10,17'd16389,17'd3748,17'd3905,17'd27442,17'd2425,17'd10092,17'd10092,17'd2936,17'd1414,17'd1416,17'd17,17'd288,17'd76536,17'd29,17'd981,17'd654,17'd1834,17'd293,17'd294,17'd12505,17'd12196,17'd16501,17'd11888,17'd10924,17'd3429,17'd654,17'd288,17'd28,17'd27,17'd1833,17'd7728,17'd7728,17'd7728,17'd7556,17'd7388,17'd7386,17'd7225,17'd6903,17'd10093,17'd11073,17'd2942,17'd1694,17'd815,17'd76613,17'd76614,17'd76615,17'd76616,17'd76617,17'd76618,17'd76619,17'd76620,17'd76621,17'd76622,17'd76623,17'd76624,17'd76625,17'd76626,17'd76627,17'd76628,17'd76629,17'd76630,17'd76631,17'd76489,17'd76632,17'd76633,17'd76558,17'd76634,17'd76635,17'd76636,17'd76420,17'd76424,17'd76561,17'd76637,17'd76638,17'd76639,17'd76640,17'd76641,17'd75753,17'd76206,17'd76500,17'd76642,17'd75938,17'd76348,17'd76643,17'd76644,17'd75850,17'd76645,17'd76570,17'd74877,17'd74188,17'd71669,17'd126,17'd1481,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd132,17'd3168,17'd6055,17'd13534,17'd75561,17'd75562,17'd76646,17'd76647,17'd76648,17'd76649,17'd76650,17'd76651,17'd76652,17'd33359,17'd76363,17'd76653,17'd76654,17'd76655,17'd17149,17'd16949,17'd16732,17'd72888,17'd16367,17'd16486,17'd16486,17'd17527,17'd76511,17'd76053,17'd76656,17'd20112,17'd76442,17'd76443,17'd75959,17'd12159,17'd12301,17'd76219,17'd68621,17'd68621,17'd6850,17'd7176,17'd7667,17'd7667,17'd5918,17'd5918,17'd5916,17'd50670,17'd5613,17'd52268,17'd52268,17'd5613,17'd27930,17'd27930,17'd7999,17'd29591,17'd8629,17'd9931,17'd9932,17'd9932,17'd9932,17'd9931,17'd69223,17'd69223,17'd10513,17'd10513,17'd9933,17'd9933,17'd9933,17'd27815,17'd69692,17'd68625,17'd68625,17'd68511,17'd29300,17'd76585,17'd76657,17'd76658,17'd76659,17'd76660,17'd76518,17'd68939,17'd76588,17'd73418,17'd76381,17'd68940,17'd76380,17'd76380,17'd76380,17'd76380,17'd76380,17'd76380,17'd74785,17'd76302,17'd68940,17'd76383,17'd76382,17'd76661,17'd68939,17'd68939,17'd76662,17'd67781,17'd68284,17'd68284,17'd74775,17'd74775,17'd76663,17'd76663,17'd76663,17'd76663,17'd67656,17'd76664,17'd74429,17'd76595,17'd76665,17'd65680,17'd64763,17'd76666,17'd76667,17'd73528,17'd17540,17'd20854,17'd13288,17'd65044,17'd66540,17'd62203,17'd67431,17'd50498,17'd10524,17'd5935,17'd76668,17'd76669,17'd929,17'd20711,17'd765,17'd52464,17'd19492,17'd38073,17'd31904,17'd76670,17'd33377,17'd37304,17'd396,17'd34003,17'd34345,17'd76607,17'd32560,17'd587,17'd76671,17'd20266,17'd766,17'd19492,17'd76672,17'd75693,17'd76673,17'd76605,17'd76674,17'd76675,17'd31255,17'd76233,17'd586,17'd177,17'd76472,17'd76472,17'd76676,17'd76677,17'd76678,17'd253,17'd278,17'd460,17'd263,17'd257,17'd270,17'd273,17'd1828,17'd1410,17'd971,17'd971,17'd971,17'd971,17'd972,17'd972
},
'{
17'd1689,17'd1689,17'd2,17'd13,17'd3,17'd1275,17'd283,17'd1,17'd15,17'd1688,17'd2422,17'd1689,17'd15,17'd1,17'd3,17'd1275,17'd283,17'd3,17'd3,17'd12,17'd3,17'd3,17'd3,17'd3,17'd3,17'd3,17'd1,17'd1412,17'd1,17'd0,17'd466,17'd2,17'd1,17'd0,17'd14,17'd1127,17'd1127,17'd1127,17'd1127,17'd1127,17'd1415,17'd16,17'd1277,17'd979,17'd19,17'd11,17'd16389,17'd5653,17'd76679,17'd76680,17'd9552,17'd6589,17'd6101,17'd67452,17'd63258,17'd6274,17'd69255,17'd63387,17'd14867,17'd67452,17'd6275,17'd7224,17'd6277,17'd9,17'd8,17'd4,17'd24,17'd24,17'd5,17'd6,17'd5,17'd5,17'd4,17'd25,17'd11,17'd3905,17'd466,17'd1127,17'd1689,17'd1689,17'd14,17'd14,17'd14,17'd2,17'd0,17'd12,17'd3,17'd3,17'd75696,17'd3748,17'd10,17'd808,17'd3748,17'd19,17'd26344,17'd63522,17'd3101,17'd2784,17'd2781,17'd1689,17'd2257,17'd2257,17'd1415,17'd16,17'd19,17'd19,17'd16,17'd2936,17'd293,17'd34,17'd294,17'd36,17'd14320,17'd58016,17'd57896,17'd11888,17'd11072,17'd10407,17'd9969,17'd981,17'd287,17'd286,17'd7728,17'd7555,17'd7557,17'd7388,17'd7388,17'd7225,17'd10269,17'd76315,17'd11073,17'd9816,17'd12036,17'd15119,17'd59497,17'd76613,17'd76681,17'd76682,17'd76683,17'd76684,17'd76685,17'd76686,17'd76687,17'd76548,17'd76688,17'd76549,17'd76689,17'd76690,17'd76691,17'd76692,17'd76263,17'd76693,17'd76409,17'd76552,17'd76553,17'd76265,17'd76633,17'd76338,17'd76694,17'd76695,17'd76696,17'd76697,17'd76698,17'd76497,17'd76699,17'd76699,17'd76700,17'd76700,17'd76701,17'd76702,17'd76703,17'd76704,17'd76705,17'd76706,17'd76707,17'd75219,17'd76708,17'd76709,17'd76710,17'd73178,17'd70831,17'd126,17'd1481,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd134,17'd132,17'd132,17'd10492,17'd3812,17'd4816,17'd76711,17'd76712,17'd76713,17'd76714,17'd76715,17'd76716,17'd76717,17'd76578,17'd76718,17'd34326,17'd76719,17'd21905,17'd76720,17'd76721,17'd76722,17'd76723,17'd76724,17'd15983,17'd16245,17'd16245,17'd16486,17'd76725,17'd76725,17'd76726,17'd20111,17'd21768,17'd76727,17'd76443,17'd76443,17'd12158,17'd75577,17'd11312,17'd11312,17'd10512,17'd6850,17'd7176,17'd7176,17'd5918,17'd5918,17'd6552,17'd5761,17'd50670,17'd76289,17'd27695,17'd27695,17'd76289,17'd5613,17'd26218,17'd6389,17'd7999,17'd8000,17'd10236,17'd10236,17'd9931,17'd9931,17'd9932,17'd9932,17'd10513,17'd10513,17'd10513,17'd10513,17'd27931,17'd27931,17'd10897,17'd10897,17'd29592,17'd31718,17'd31718,17'd68625,17'd68625,17'd68511,17'd76445,17'd68512,17'd68512,17'd68513,17'd76446,17'd68828,17'd76518,17'd74076,17'd76461,17'd76461,17'd68732,17'd76461,17'd76461,17'd76461,17'd76728,17'd76728,17'd76518,17'd76586,17'd76660,17'd76660,17'd76659,17'd76516,17'd76516,17'd76729,17'd76657,17'd76657,17'd68403,17'd68403,17'd76730,17'd76730,17'd76730,17'd76731,17'd76732,17'd67279,17'd76733,17'd76734,17'd14855,17'd64763,17'd12765,17'd18377,17'd25883,17'd76735,17'd76736,17'd22256,17'd12910,17'd76737,17'd76738,17'd67166,17'd45403,17'd4865,17'd69614,17'd76739,17'd33999,17'd24164,17'd20863,17'd765,17'd19602,17'd28313,17'd26721,17'd28427,17'd76740,17'd76071,17'd37045,17'd396,17'd36604,17'd76741,17'd76742,17'd76743,17'd32560,17'd16006,17'd76671,17'd16263,17'd28313,17'd52277,17'd36749,17'd76069,17'd38074,17'd34511,17'd76742,17'd38461,17'd76607,17'd76744,17'd76745,17'd16264,17'd76239,17'd76746,17'd76747,17'd76678,17'd73325,17'd27824,17'd278,17'd460,17'd266,17'd266,17'd968,17'd272,17'd1828,17'd1828,17'd1828,17'd1410,17'd1410,17'd1410,17'd803,17'd803
},
'{
17'd2592,17'd2781,17'd14,17'd2,17'd3,17'd1275,17'd650,17'd1412,17'd1830,17'd1689,17'd2422,17'd3250,17'd1967,17'd15,17'd3,17'd1275,17'd283,17'd3,17'd12,17'd12,17'd3,17'd283,17'd3,17'd3,17'd283,17'd3,17'd1412,17'd4884,17'd4884,17'd1,17'd2,17'd2,17'd1,17'd0,17'd14,17'd14,17'd1127,17'd1127,17'd1127,17'd1127,17'd17187,17'd1414,17'd17,17'd979,17'd808,17'd11,17'd21,17'd5652,17'd6275,17'd76679,17'd6107,17'd67577,17'd6100,17'd5964,17'd74233,17'd64125,17'd63258,17'd14867,17'd67452,17'd67307,17'd5801,17'd5653,17'd5653,17'd5651,17'd5647,17'd4,17'd23,17'd284,17'd5,17'd6,17'd6,17'd5,17'd4,17'd23,17'd21,17'd18,17'd2,17'd1127,17'd1688,17'd1689,17'd14,17'd14,17'd14,17'd14,17'd2,17'd0,17'd0,17'd3,17'd18,17'd19,17'd11,17'd11,17'd75696,17'd6108,17'd979,17'd22965,17'd76748,17'd3251,17'd3250,17'd2781,17'd3752,17'd3429,17'd2597,17'd1416,17'd979,17'd1128,17'd3905,17'd1415,17'd1693,17'd293,17'd471,17'd15878,17'd58504,17'd14989,17'd14989,17'd58504,17'd13944,17'd76749,17'd76750,17'd10544,17'd2118,17'd287,17'd1833,17'd8047,17'd8047,17'd7557,17'd7388,17'd7556,17'd10093,17'd72282,17'd9554,17'd9554,17'd11073,17'd12333,17'd1279,17'd76751,17'd76752,17'd76753,17'd76754,17'd76755,17'd76756,17'd76757,17'd76758,17'd76759,17'd76760,17'd76761,17'd76762,17'd76763,17'd76764,17'd76765,17'd76766,17'd76767,17'd76768,17'd76769,17'd76770,17'd76771,17'd76772,17'd76773,17'd76774,17'd76775,17'd76776,17'd76777,17'd75845,17'd75936,17'd76778,17'd76700,17'd76497,17'd76779,17'd76780,17'd76781,17'd76782,17'd76783,17'd76784,17'd76785,17'd76786,17'd76787,17'd76788,17'd74877,17'd72986,17'd72654,17'd71260,17'd1481,17'd132,17'd11541,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd134,17'd132,17'd132,17'd2861,17'd3512,17'd6532,17'd76789,17'd76790,17'd76791,17'd76792,17'd76793,17'd31705,17'd76794,17'd76795,17'd76796,17'd17493,17'd76797,17'd76798,17'd76799,17'd76800,17'd18968,17'd76801,17'd15219,17'd19220,17'd15849,17'd15983,17'd16245,17'd76802,17'd76802,17'd76803,17'd20111,17'd76804,17'd21768,17'd76443,17'd76444,17'd12158,17'd12003,17'd76805,17'd11570,17'd11312,17'd10512,17'd6850,17'd7176,17'd6704,17'd6704,17'd5918,17'd5918,17'd5916,17'd5915,17'd76289,17'd76289,17'd76289,17'd76289,17'd5003,17'd5159,17'd28304,17'd7999,17'd8000,17'd8000,17'd8629,17'd29591,17'd8629,17'd9931,17'd10513,17'd10513,17'd10777,17'd10513,17'd50487,17'd50487,17'd76291,17'd76291,17'd28533,17'd76806,17'd31888,17'd29593,17'd31718,17'd31718,17'd68625,17'd68625,17'd68625,17'd68511,17'd29300,17'd29300,17'd76585,17'd76729,17'd76660,17'd68629,17'd68629,17'd76658,17'd76659,17'd76659,17'd76659,17'd76807,17'd76807,17'd76808,17'd76809,17'd76810,17'd76445,17'd76445,17'd68626,17'd68626,17'd76811,17'd76811,17'd29300,17'd76585,17'd29027,17'd76812,17'd76813,17'd76731,17'd76732,17'd74652,17'd74545,17'd14169,17'd13413,17'd76814,17'd12766,17'd27939,17'd24806,17'd13052,17'd62310,17'd62561,17'd12769,17'd66185,17'd11865,17'd67043,17'd65942,17'd76815,17'd76531,17'd37956,17'd24164,17'd18758,17'd26009,17'd76816,17'd51858,17'd28427,17'd52277,17'd76670,17'd76817,17'd36750,17'd76818,17'd396,17'd36325,17'd34345,17'd76819,17'd76820,17'd31412,17'd16140,17'd30046,17'd16264,17'd76821,17'd75980,17'd76154,17'd75979,17'd38074,17'd33848,17'd34667,17'd38461,17'd76606,17'd76607,17'd30945,17'd39329,17'd16746,17'd68847,17'd279,17'd182,17'd73644,17'd15240,17'd804,17'd254,17'd265,17'd262,17'd7539,17'd640,17'd1687,17'd1687,17'd1828,17'd1828,17'd1410,17'd1828,17'd803,17'd644
},
'{
17'd2784,17'd2592,17'd1689,17'd14,17'd12,17'd806,17'd283,17'd1412,17'd1830,17'd3249,17'd3250,17'd2422,17'd1688,17'd1830,17'd283,17'd3,17'd283,17'd3,17'd3,17'd3,17'd3,17'd3,17'd3,17'd3,17'd3,17'd283,17'd650,17'd650,17'd650,17'd283,17'd12,17'd13,17'd2,17'd0,17'd1,17'd1,17'd14,17'd1127,17'd1127,17'd1127,17'd17187,17'd16,17'd18,17'd19,17'd10,17'd25,17'd1690,17'd2937,17'd5652,17'd5801,17'd5799,17'd75044,17'd5967,17'd76535,17'd14187,17'd14187,17'd63117,17'd14988,17'd76822,17'd76823,17'd75696,17'd75696,17'd6108,17'd75696,17'd1413,17'd8,17'd4,17'd23,17'd24,17'd24,17'd3594,17'd3753,17'd5,17'd4,17'd25,17'd808,17'd18,17'd22965,17'd2594,17'd4247,17'd15,17'd14,17'd1127,17'd14,17'd15,17'd1,17'd0,17'd2,17'd979,17'd19,17'd18,17'd19,17'd979,17'd3748,17'd808,17'd3748,17'd4247,17'd76824,17'd76825,17'd2934,17'd68191,17'd6265,17'd3250,17'd4247,17'd17,17'd1277,17'd19,17'd16,17'd1414,17'd10268,17'd76826,17'd12653,17'd58504,17'd66091,17'd76827,17'd76828,17'd76828,17'd14598,17'd13945,17'd76829,17'd10544,17'd2118,17'd287,17'd7555,17'd7555,17'd7555,17'd7728,17'd8988,17'd7061,17'd7061,17'd7060,17'd6744,17'd76830,17'd11209,17'd35,17'd59497,17'd76831,17'd76832,17'd76833,17'd76834,17'd76835,17'd76836,17'd76837,17'd76837,17'd76838,17'd76762,17'd76839,17'd76840,17'd76841,17'd76766,17'd76768,17'd76769,17'd76770,17'd76842,17'd76843,17'd76844,17'd76845,17'd76846,17'd76271,17'd76700,17'd76847,17'd75446,17'd76848,17'd76849,17'd76850,17'd76851,17'd76702,17'd76703,17'd75938,17'd76501,17'd76568,17'd76785,17'd76852,17'd73832,17'd73502,17'd73713,17'd75451,17'd75452,17'd72654,17'd73073,17'd127,17'd134,17'd131,17'd131,17'd132,17'd130,17'd130,17'd130,17'd132,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd1197,17'd133,17'd132,17'd135,17'd132,17'd3168,17'd4814,17'd2865,17'd3029,17'd76853,17'd76854,17'd76855,17'd76856,17'd76857,17'd76858,17'd76859,17'd76860,17'd76212,17'd76861,17'd76862,17'd31086,17'd76863,17'd76864,17'd76865,17'd20111,17'd76866,17'd76867,17'd76868,17'd76869,17'd76870,17'd76802,17'd76871,17'd19981,17'd20533,17'd15078,17'd76872,17'd76873,17'd76874,17'd76444,17'd76875,17'd11178,17'd11312,17'd11570,17'd11570,17'd10512,17'd6705,17'd6705,17'd6704,17'd5918,17'd5916,17'd5915,17'd50670,17'd50670,17'd5914,17'd50670,17'd5003,17'd5612,17'd5158,17'd5332,17'd6388,17'd6387,17'd6707,17'd6707,17'd8303,17'd8154,17'd8154,17'd9090,17'd9394,17'd9394,17'd10513,17'd10513,17'd27931,17'd27931,17'd27931,17'd9933,17'd10380,17'd10380,17'd10380,17'd10380,17'd10380,17'd10380,17'd10380,17'd10779,17'd10779,17'd7012,17'd29163,17'd29163,17'd29163,17'd29163,17'd29163,17'd68173,17'd29163,17'd29299,17'd29299,17'd29299,17'd29299,17'd12625,17'd12625,17'd12625,17'd10779,17'd12625,17'd12625,17'd12625,17'd68626,17'd68282,17'd68173,17'd76876,17'd7180,17'd76877,17'd76878,17'd29028,17'd76879,17'd76880,17'd15097,17'd76881,17'd17176,17'd30334,17'd26115,17'd76882,17'd13052,17'd12171,17'd12631,17'd12769,17'd76883,17'd18754,17'd10905,17'd43462,17'd3872,17'd39178,17'd2738,17'd59766,17'd18759,17'd76884,17'd51674,17'd52277,17'd761,17'd761,17'd76885,17'd27821,17'd36750,17'd396,17'd396,17'd36457,17'd33377,17'd35909,17'd76603,17'd76233,17'd618,17'd16140,17'd76074,17'd31412,17'd38461,17'd36457,17'd76886,17'd36750,17'd76887,17'd76887,17'd34667,17'd36182,17'd76607,17'd176,17'd39329,17'd588,17'd68749,17'd68960,17'd182,17'd639,17'd1683,17'd639,17'd804,17'd804,17'd969,17'd459,17'd968,17'd272,17'd643,17'd644,17'd1687,17'd1828,17'd1963,17'd24165,17'd645,17'd643
},
'{
17'd63254,17'd2782,17'd3250,17'd1689,17'd2,17'd12,17'd3,17'd1412,17'd1830,17'd15,17'd1689,17'd2422,17'd1688,17'd15,17'd1,17'd3,17'd283,17'd283,17'd3,17'd3,17'd3,17'd3,17'd3,17'd3,17'd283,17'd283,17'd283,17'd650,17'd650,17'd283,17'd3,17'd12,17'd0,17'd1,17'd1,17'd1,17'd14,17'd1127,17'd1127,17'd1127,17'd1415,17'd16,17'd18,17'd19,17'd10,17'd25,17'd1691,17'd1690,17'd1413,17'd5651,17'd5653,17'd75158,17'd6275,17'd75046,17'd14187,17'd75159,17'd76888,17'd76822,17'd4732,17'd4732,17'd3748,17'd75696,17'd75490,17'd3748,17'd16389,17'd9,17'd4,17'd4,17'd24,17'd24,17'd3594,17'd3753,17'd6,17'd5,17'd4,17'd25,17'd19,17'd1416,17'd2595,17'd4247,17'd1127,17'd1127,17'd14,17'd14,17'd14,17'd14,17'd2,17'd2,17'd1277,17'd19,17'd19,17'd19,17'd19,17'd979,17'd10,17'd808,17'd650,17'd2594,17'd76825,17'd60150,17'd3901,17'd67808,17'd7371,17'd2781,17'd52621,17'd2597,17'd16,17'd1276,17'd1277,17'd1414,17'd3593,17'd12196,17'd4893,17'd66091,17'd76889,17'd76890,17'd76891,17'd76892,17'd15361,17'd58504,17'd76893,17'd10092,17'd1415,17'd2938,17'd653,17'd74808,17'd71091,17'd74808,17'd8988,17'd7728,17'd7061,17'd4430,17'd4431,17'd3754,17'd2427,17'd76894,17'd76895,17'd76896,17'd76897,17'd76898,17'd76899,17'd76900,17'd76901,17'd76902,17'd76903,17'd76904,17'd76905,17'd76906,17'd76907,17'd76908,17'd76909,17'd76845,17'd76910,17'd76911,17'd76560,17'd76344,17'd76912,17'd75935,17'd76500,17'd76913,17'd76914,17'd76915,17'd76916,17'd76917,17'd76918,17'd76207,17'd75938,17'd76919,17'd75555,17'd76351,17'd76920,17'd76921,17'd73607,17'd76922,17'd76923,17'd74520,17'd76924,17'd76925,17'd73073,17'd72754,17'd130,17'd132,17'd132,17'd134,17'd130,17'd130,17'd136,17'd130,17'd132,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd1197,17'd133,17'd133,17'd134,17'd132,17'd357,17'd4336,17'd13534,17'd76926,17'd76927,17'd6371,17'd76928,17'd76929,17'd76930,17'd76575,17'd76931,17'd76932,17'd76933,17'd76934,17'd76935,17'd76936,17'd76799,17'd76937,17'd76938,17'd76865,17'd76939,17'd76804,17'd76940,17'd76869,17'd76869,17'd76870,17'd76941,17'd76940,17'd20533,17'd21768,17'd76942,17'd76943,17'd76944,17'd6385,17'd11034,17'd11311,17'd11178,17'd11035,17'd10512,17'd10512,17'd6705,17'd6704,17'd6552,17'd5918,17'd5917,17'd5916,17'd50670,17'd76289,17'd5914,17'd6384,17'd5611,17'd5612,17'd5612,17'd5158,17'd5331,17'd5332,17'd6553,17'd6553,17'd8303,17'd8303,17'd8154,17'd8154,17'd9090,17'd9394,17'd9394,17'd10513,17'd10513,17'd27931,17'd9933,17'd9933,17'd10380,17'd10380,17'd10380,17'd10380,17'd10380,17'd10380,17'd10380,17'd10380,17'd10516,17'd10779,17'd10779,17'd10779,17'd10779,17'd10779,17'd10779,17'd10779,17'd10779,17'd10779,17'd10779,17'd10779,17'd10516,17'd10516,17'd10516,17'd10516,17'd10516,17'd10779,17'd10779,17'd10779,17'd68511,17'd76945,17'd7013,17'd76876,17'd76877,17'd76878,17'd29028,17'd76946,17'd66529,17'd76947,17'd13284,17'd17069,17'd30490,17'd30033,17'd23983,17'd12313,17'd12171,17'd30034,17'd12479,17'd76948,17'd66792,17'd68743,17'd46596,17'd40099,17'd54422,17'd37956,17'd24164,17'd24953,17'd26009,17'd76949,17'd76950,17'd76951,17'd51859,17'd76952,17'd76953,17'd76071,17'd36604,17'd76818,17'd396,17'd76954,17'd33848,17'd76885,17'd31564,17'd31564,17'd586,17'd586,17'd32883,17'd31255,17'd34668,17'd37305,17'd37046,17'd34003,17'd36604,17'd36750,17'd36182,17'd35062,17'd33376,17'd218,17'd619,17'd223,17'd76955,17'd462,17'd1826,17'd1548,17'd1826,17'd639,17'd965,17'd965,17'd49713,17'd265,17'd257,17'd272,17'd643,17'd643,17'd1687,17'd1828,17'd645,17'd1963,17'd803,17'd206
},
'{
17'd3904,17'd3904,17'd4246,17'd7214,17'd466,17'd12,17'd3,17'd3,17'd1412,17'd1830,17'd1967,17'd1688,17'd1831,17'd1689,17'd15,17'd1,17'd283,17'd283,17'd283,17'd3,17'd3,17'd3,17'd3,17'd3,17'd283,17'd3,17'd1275,17'd465,17'd651,17'd651,17'd1275,17'd806,17'd12,17'd3,17'd1,17'd1,17'd15,17'd14,17'd14,17'd14,17'd2,17'd2,17'd18,17'd11,17'd21,17'd25,17'd1691,17'd1691,17'd5,17'd4,17'd1413,17'd5651,17'd75262,17'd75158,17'd5799,17'd5799,17'd76956,17'd6277,17'd5652,17'd808,17'd10,17'd3748,17'd5969,17'd979,17'd808,17'd9,17'd4,17'd4,17'd5,17'd5,17'd3594,17'd3594,17'd6,17'd5,17'd4,17'd9,17'd808,17'd18,17'd3430,17'd15745,17'd2594,17'd4247,17'd14,17'd14,17'd14,17'd1127,17'd14,17'd2,17'd2,17'd0,17'd1,17'd1,17'd18,17'd18,17'd19,17'd808,17'd977,17'd806,17'd17917,17'd37047,17'd15877,17'd13943,17'd76957,17'd76957,17'd2593,17'd3101,17'd1831,17'd15,17'd1276,17'd1415,17'd2597,17'd10546,17'd4738,17'd14443,17'd76958,17'd76959,17'd76960,17'd76961,17'd76962,17'd76963,17'd14744,17'd12505,17'd10092,17'd30,17'd30,17'd981,17'd76964,17'd76964,17'd76965,17'd76965,17'd76965,17'd288,17'd4091,17'd3755,17'd655,17'd76966,17'd76967,17'd76968,17'd76969,17'd76970,17'd76971,17'd76972,17'd76973,17'd76974,17'd76975,17'd76975,17'd76341,17'd76976,17'd76561,17'd76977,17'd76978,17'd76979,17'd76980,17'd76037,17'd76981,17'd76982,17'd76983,17'd76919,17'd75755,17'd76130,17'd76984,17'd76985,17'd76986,17'd76981,17'd76207,17'd76347,17'd76349,17'd76987,17'd76988,17'd76989,17'd76990,17'd74872,17'd76991,17'd73504,17'd73724,17'd72986,17'd71578,17'd76992,17'd71477,17'd136,17'd130,17'd132,17'd132,17'd128,17'd130,17'd136,17'd136,17'd136,17'd130,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd133,17'd133,17'd134,17'd132,17'd135,17'd76993,17'd5466,17'd76994,17'd76995,17'd76996,17'd76997,17'd76998,17'd76999,17'd77000,17'd17864,17'd77001,17'd77002,17'd77003,17'd76212,17'd77004,17'd77005,17'd17030,17'd77006,17'd77007,17'd77008,17'd76865,17'd77009,17'd76726,17'd77010,17'd76656,17'd77011,17'd77011,17'd19981,17'd76942,17'd14152,17'd77012,17'd77013,17'd6845,17'd23630,17'd23112,17'd23283,17'd24481,17'd24481,17'd23976,17'd11035,17'd7176,17'd5761,17'd6552,17'd5916,17'd5916,17'd5915,17'd50670,17'd5914,17'd6384,17'd5481,17'd5611,17'd5611,17'd5611,17'd5612,17'd5331,17'd5332,17'd6388,17'd6218,17'd6218,17'd6553,17'd6553,17'd5919,17'd6221,17'd6392,17'd28058,17'd8780,17'd8780,17'd8780,17'd7668,17'd7500,17'd7500,17'd7669,17'd7669,17'd8780,17'd8780,17'd8780,17'd8780,17'd8780,17'd7669,17'd7669,17'd7669,17'd7669,17'd7669,17'd7669,17'd7669,17'd7669,17'd7669,17'd7669,17'd7669,17'd8471,17'd8471,17'd8471,17'd8471,17'd8471,17'd8155,17'd13281,17'd13281,17'd7013,17'd7013,17'd7502,17'd7014,17'd7015,17'd16374,17'd14427,17'd14576,17'd13680,17'd13283,17'd12627,17'd77014,17'd25882,17'd24156,17'd77015,17'd61930,17'd12013,17'd77016,17'd77017,17'd66187,17'd11046,17'd77018,17'd3870,17'd7025,17'd22956,17'd35768,17'd1236,17'd61026,17'd76950,17'd583,17'd583,17'd77019,17'd52367,17'd760,17'd76817,17'd77020,17'd77021,17'd77022,17'd396,17'd36750,17'd77023,17'd52465,17'd31904,17'd38335,17'd77024,17'd76233,17'd31255,17'd34345,17'd37305,17'd77025,17'd77026,17'd77027,17'd77028,17'd77029,17'd77030,17'd32884,17'd438,17'd615,17'd1238,17'd39627,17'd612,17'd213,17'd251,17'd250,17'd180,17'd252,17'd181,17'd1123,17'd73987,17'd969,17'd257,17'd646,17'd270,17'd272,17'd644,17'd803,17'd645,17'd645,17'd803,17'd206
},
'{
17'd65576,17'd4088,17'd4245,17'd4246,17'd1688,17'd2,17'd1,17'd1,17'd1412,17'd3749,17'd1830,17'd1689,17'd1831,17'd1688,17'd1967,17'd1830,17'd1412,17'd283,17'd283,17'd3,17'd3,17'd12,17'd3,17'd3,17'd283,17'd3,17'd806,17'd1275,17'd651,17'd77031,17'd465,17'd1275,17'd3,17'd3,17'd283,17'd1,17'd1,17'd15,17'd15,17'd0,17'd2,17'd12,17'd19,17'd10,17'd21,17'd25,17'd1691,17'd7384,17'd3594,17'd5,17'd4,17'd9,17'd6108,17'd75263,17'd5653,17'd5653,17'd6277,17'd6277,17'd5512,17'd5647,17'd10,17'd11,17'd19,17'd19,17'd10,17'd25,17'd9,17'd4,17'd4,17'd5,17'd5,17'd3594,17'd6,17'd5,17'd4,17'd8,17'd9,17'd10,17'd16636,17'd8971,17'd77032,17'd2594,17'd1127,17'd1127,17'd1127,17'd1127,17'd14,17'd14,17'd2,17'd0,17'd0,17'd0,17'd16,17'd18,17'd19,17'd11,17'd2933,17'd465,17'd1412,17'd3250,17'd15496,17'd15359,17'd64116,17'd4737,17'd76957,17'd3901,17'd34512,17'd3252,17'd2936,17'd9969,17'd17187,17'd10092,17'd2783,17'd64117,17'd77033,17'd77034,17'd77035,17'd76960,17'd76961,17'd76962,17'd77036,17'd14744,17'd4738,17'd77037,17'd10407,17'd469,17'd1693,17'd3102,17'd77038,17'd77039,17'd77040,17'd77039,17'd76830,17'd9554,17'd981,17'd1693,17'd77041,17'd76967,17'd77042,17'd77043,17'd77044,17'd77045,17'd77046,17'd77047,17'd77048,17'd77049,17'd77050,17'd77051,17'd77052,17'd77053,17'd77054,17'd77055,17'd77056,17'd77057,17'd77058,17'd77058,17'd76783,17'd77059,17'd77060,17'd77061,17'd77062,17'd77063,17'd76918,17'd76126,17'd76982,17'd76348,17'd74869,17'd74750,17'd74994,17'd75759,17'd75759,17'd77064,17'd73829,17'd74521,17'd75108,17'd72871,17'd77065,17'd139,17'd130,17'd130,17'd132,17'd132,17'd130,17'd130,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd133,17'd133,17'd132,17'd132,17'd132,17'd10492,17'd77066,17'd3659,17'd19169,17'd77067,17'd77068,17'd77069,17'd77070,17'd17982,17'd77071,17'd30321,17'd77072,17'd77073,17'd77074,17'd77075,17'd31711,17'd77076,17'd77077,17'd77078,17'd77079,17'd77080,17'd77081,17'd76939,17'd76726,17'd76867,17'd76940,17'd76871,17'd77082,17'd20533,17'd14152,17'd14284,17'd77083,17'd7328,17'd6211,17'd6384,17'd23461,17'd24150,17'd6068,17'd24481,17'd6850,17'd7176,17'd5918,17'd5761,17'd76289,17'd50670,17'd5915,17'd5916,17'd6384,17'd5913,17'd5481,17'd5481,17'd5611,17'd5611,17'd5612,17'd5158,17'd5331,17'd5331,17'd6389,17'd6389,17'd6389,17'd6218,17'd5614,17'd5615,17'd6221,17'd6221,17'd28058,17'd8780,17'd7668,17'd7668,17'd7668,17'd7500,17'd7500,17'd8780,17'd8780,17'd10513,17'd10513,17'd10513,17'd9657,17'd7668,17'd7668,17'd7668,17'd7669,17'd7669,17'd7500,17'd7500,17'd7500,17'd7500,17'd7500,17'd7500,17'd6557,17'd6557,17'd6557,17'd8155,17'd8155,17'd7179,17'd7179,17'd7179,17'd7013,17'd68049,17'd7014,17'd66419,17'd77084,17'd7504,17'd13680,17'd13411,17'd77085,17'd77086,17'd77087,17'd74653,17'd24946,17'd11861,17'd11715,17'd19354,17'd77088,17'd77089,17'd65692,17'd10522,17'd18980,17'd48558,17'd6866,17'd77090,17'd77091,17'd77092,17'd77093,17'd77019,17'd77094,17'd77095,17'd77096,17'd52278,17'd77097,17'd27821,17'd580,17'd77098,17'd77022,17'd77022,17'd36457,17'd76071,17'd77099,17'd761,17'd76672,17'd76672,17'd31564,17'd76740,17'd34345,17'd37447,17'd77100,17'd77101,17'd77102,17'd77103,17'd77104,17'd77105,17'd77106,17'd39184,17'd20266,17'd1541,17'd27948,17'd635,17'd19102,17'd250,17'd280,17'd24000,17'd23489,17'd20271,17'd182,17'd1683,17'd1123,17'd595,17'd256,17'd257,17'd270,17'd272,17'd644,17'd803,17'd645,17'd645,17'd644,17'd643
},
'{
17'd65576,17'd9960,17'd4428,17'd4245,17'd2422,17'd1689,17'd15,17'd1,17'd1412,17'd1412,17'd1412,17'd14,17'd1688,17'd1831,17'd1689,17'd3249,17'd1,17'd283,17'd283,17'd3,17'd3,17'd12,17'd3,17'd3,17'd283,17'd3,17'd806,17'd1275,17'd977,17'd807,17'd977,17'd2591,17'd1275,17'd1275,17'd1275,17'd283,17'd283,17'd3,17'd3,17'd12,17'd12,17'd12,17'd806,17'd2933,17'd25,17'd4,17'd5,17'd5,17'd3594,17'd3594,17'd5,17'd4,17'd9,17'd16389,17'd16389,17'd16389,17'd5652,17'd5652,17'd6277,17'd5651,17'd808,17'd11,17'd19,17'd18,17'd11,17'd21,17'd25,17'd4,17'd4,17'd5,17'd5,17'd5,17'd5,17'd5,17'd5,17'd8,17'd8,17'd1413,17'd21,17'd20404,17'd15745,17'd15745,17'd2594,17'd4247,17'd1127,17'd14,17'd14,17'd14,17'd14,17'd14,17'd14,17'd2,17'd0,17'd1,17'd12,17'd12,17'd10,17'd16389,17'd4732,17'd1,17'd3252,17'd61679,17'd15359,17'd6730,17'd14071,17'd3751,17'd3592,17'd15496,17'd2934,17'd7371,17'd3249,17'd3249,17'd76826,17'd76893,17'd77107,17'd14189,17'd76889,17'd77108,17'd77109,17'd77110,17'd77111,17'd76892,17'd76827,17'd64660,17'd76957,17'd77041,17'd77037,17'd10407,17'd2936,17'd65450,17'd77112,17'd77112,17'd77113,17'd77039,17'd9554,17'd3595,17'd31,17'd1834,17'd12784,17'd77114,17'd77115,17'd77116,17'd77117,17'd77118,17'd77119,17'd77120,17'd76272,17'd76561,17'd76700,17'd76703,17'd77121,17'd77122,17'd77058,17'd76783,17'd77123,17'd77123,17'd77124,17'd77125,17'd77061,17'd77126,17'd76981,17'd77127,17'd77128,17'd76428,17'd77129,17'd75848,17'd77130,17'd76786,17'd77131,17'd77132,17'd75851,17'd77133,17'd76042,17'd75854,17'd74050,17'd72654,17'd67858,17'd130,17'd132,17'd132,17'd128,17'd128,17'd130,17'd130,17'd130,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd2698,17'd77134,17'd3512,17'd77135,17'd77136,17'd77137,17'd77138,17'd77139,17'd77140,17'd77141,17'd77142,17'd76999,17'd77143,17'd77144,17'd77145,17'd33196,17'd35465,17'd77146,17'd77147,17'd77148,17'd77149,17'd77150,17'd14152,17'd19981,17'd76803,17'd77151,17'd76726,17'd77152,17'd77153,17'd77154,17'd77154,17'd14548,17'd77155,17'd24480,17'd6547,17'd6212,17'd23629,17'd23630,17'd5916,17'd8931,17'd7667,17'd7176,17'd8931,17'd5613,17'd5613,17'd50670,17'd5915,17'd5914,17'd5913,17'd50670,17'd50670,17'd50670,17'd76289,17'd5158,17'd5158,17'd5158,17'd5158,17'd5331,17'd5331,17'd26218,17'd26218,17'd5332,17'd5332,17'd6387,17'd6707,17'd9090,17'd9090,17'd9090,17'd6220,17'd6220,17'd6220,17'd6391,17'd6391,17'd6391,17'd9090,17'd9657,17'd9657,17'd9657,17'd9657,17'd9657,17'd7668,17'd7500,17'd7500,17'd7500,17'd7500,17'd7500,17'd7500,17'd6555,17'd6555,17'd77156,17'd77156,17'd77157,17'd77157,17'd6560,17'd30032,17'd30032,17'd7671,17'd7014,17'd7014,17'd7181,17'd7503,17'd31090,17'd12472,17'd12310,17'd12007,17'd12007,17'd77158,17'd25632,17'd24658,17'd20549,17'd77159,17'd11438,17'd11324,17'd77160,17'd77161,17'd5350,17'd67561,17'd7849,17'd3868,17'd77162,17'd21159,17'd77163,17'd77164,17'd77165,17'd77166,17'd77167,17'd77166,17'd77168,17'd77169,17'd77168,17'd581,17'd77170,17'd77171,17'd77025,17'd77172,17'd76741,17'd35909,17'd31255,17'd31904,17'd38335,17'd31730,17'd76885,17'd759,17'd37447,17'd77100,17'd77173,17'd77174,17'd395,17'd77175,17'd77029,17'd77176,17'd76532,17'd15874,17'd223,17'd612,17'd963,17'd591,17'd77177,17'd250,17'd75485,17'd77178,17'd23489,17'd24000,17'd15626,17'd402,17'd1123,17'd595,17'd256,17'd256,17'd270,17'd272,17'd644,17'd803,17'd645,17'd803,17'd644,17'd643
},
'{
17'd65576,17'd9960,17'd3903,17'd4428,17'd2935,17'd3250,17'd1967,17'd1830,17'd1,17'd283,17'd1412,17'd1,17'd1127,17'd1831,17'd3250,17'd1967,17'd0,17'd3,17'd283,17'd283,17'd3,17'd12,17'd12,17'd3,17'd3,17'd3,17'd806,17'd1275,17'd2591,17'd977,17'd977,17'd977,17'd465,17'd465,17'd1275,17'd1275,17'd650,17'd283,17'd283,17'd3,17'd3,17'd806,17'd2933,17'd2591,17'd23,17'd4,17'd5,17'd6,17'd5,17'd5,17'd5,17'd5,17'd4,17'd23,17'd25,17'd25,17'd5651,17'd16389,17'd16389,17'd16389,17'd808,17'd808,17'd10,17'd20404,17'd11,17'd11,17'd25,17'd9,17'd4,17'd4,17'd5,17'd5,17'd5,17'd5,17'd5,17'd5,17'd8,17'd8,17'd9,17'd10,17'd13,17'd2595,17'd2594,17'd2594,17'd1127,17'd14,17'd14,17'd14,17'd15,17'd14,17'd1127,17'd1127,17'd0,17'd1,17'd12,17'd13,17'd1277,17'd1277,17'd283,17'd5051,17'd63116,17'd2784,17'd15496,17'd53228,17'd5511,17'd4737,17'd70968,17'd6730,17'd5203,17'd3901,17'd2592,17'd2781,17'd10406,17'd76826,17'd76893,17'd12784,17'd64660,17'd76889,17'd77179,17'd77180,17'd77181,17'd77182,17'd77183,17'd77184,17'd76828,17'd4737,17'd76893,17'd10545,17'd2597,17'd2596,17'd9969,17'd76395,17'd77185,17'd77112,17'd77186,17'd18037,17'd652,17'd289,17'd2597,17'd12196,17'd77187,17'd77188,17'd77189,17'd77190,17'd76334,17'd77191,17'd77192,17'd77193,17'd76696,17'd77194,17'd77195,17'd77196,17'd77197,17'd77198,17'd77199,17'd77200,17'd77125,17'd77201,17'd76349,17'd77202,17'd77203,17'd77128,17'd77204,17'd76918,17'd76919,17'd77205,17'd76785,17'd77206,17'd73606,17'd76787,17'd74053,17'd73391,17'd74405,17'd75451,17'd75667,17'd72655,17'd138,17'd132,17'd132,17'd132,17'd130,17'd130,17'd130,17'd132,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd134,17'd77207,17'd3812,17'd4816,17'd77208,17'd77209,17'd77210,17'd77211,17'd77212,17'd77213,17'd77214,17'd77215,17'd77216,17'd77217,17'd77218,17'd77219,17'd77220,17'd77076,17'd77221,17'd77222,17'd77223,17'd77224,17'd77225,17'd14284,17'd76866,17'd76512,17'd77151,17'd76940,17'd77226,17'd77227,17'd14408,17'd14548,17'd77227,17'd46126,17'd23975,17'd26827,17'd6382,17'd23630,17'd6384,17'd6213,17'd7176,17'd7667,17'd7667,17'd6552,17'd27930,17'd76289,17'd27695,17'd6549,17'd5913,17'd76289,17'd76289,17'd50670,17'd50670,17'd27930,17'd5158,17'd5158,17'd5612,17'd5158,17'd5158,17'd26218,17'd26218,17'd5158,17'd5331,17'd5332,17'd6388,17'd7999,17'd29591,17'd8154,17'd8154,17'd6219,17'd6219,17'd6220,17'd6220,17'd6220,17'd8154,17'd8304,17'd8304,17'd8304,17'd8304,17'd9657,17'd7668,17'd7500,17'd7500,17'd7500,17'd7500,17'd7500,17'd7177,17'd6222,17'd6222,17'd6393,17'd6393,17'd77228,17'd77228,17'd11040,17'd6561,17'd6561,17'd6856,17'd6856,17'd7330,17'd7841,17'd12626,17'd12006,17'd33693,17'd11857,17'd11041,17'd11581,17'd11435,17'd10902,17'd21935,17'd10242,17'd10243,17'd10068,17'd77229,17'd77230,17'd77231,17'd5023,17'd5772,17'd4053,17'd55881,17'd57102,17'd77232,17'd1522,17'd26963,17'd77233,17'd77171,17'd77234,17'd77020,17'd77235,17'd77236,17'd581,17'd77020,17'd77172,17'd77022,17'd77237,17'd579,17'd77238,17'd76740,17'd31255,17'd36324,17'd38335,17'd77239,17'd77097,17'd77240,17'd77241,17'd77242,17'd77243,17'd77244,17'd395,17'd77245,17'd77246,17'd77247,17'd15874,17'd75486,17'd68960,17'd638,17'd19102,17'd68846,17'd590,17'd1397,17'd463,17'd75597,17'd17298,17'd1543,17'd17185,17'd15492,17'd15240,17'd456,17'd266,17'd256,17'd270,17'd272,17'd644,17'd645,17'd645,17'd644,17'd644,17'd644
},
'{
17'd7042,17'd9960,17'd3903,17'd4892,17'd3427,17'd2935,17'd1689,17'd1,17'd12,17'd3,17'd283,17'd1412,17'd15,17'd1688,17'd2422,17'd3250,17'd2,17'd3,17'd283,17'd283,17'd3,17'd12,17'd12,17'd12,17'd806,17'd806,17'd1275,17'd1275,17'd2591,17'd2591,17'd2421,17'd978,17'd977,17'd2591,17'd2933,17'd2933,17'd465,17'd465,17'd1275,17'd806,17'd806,17'd8814,17'd2933,17'd2933,17'd23,17'd4,17'd6,17'd6,17'd6,17'd6,17'd6,17'd3594,17'd5,17'd24,17'd23,17'd25,17'd5652,17'd3748,17'd3748,17'd3748,17'd979,17'd10,17'd10,17'd1128,17'd2423,17'd806,17'd21,17'd25,17'd23,17'd4,17'd5,17'd5,17'd5,17'd5,17'd5,17'd5,17'd5,17'd6,17'd8,17'd25,17'd3,17'd0,17'd466,17'd15745,17'd2594,17'd4247,17'd1967,17'd1967,17'd3249,17'd1967,17'd1127,17'd1127,17'd2,17'd2,17'd0,17'd0,17'd1415,17'd1415,17'd0,17'd4884,17'd5051,17'd1412,17'd1831,17'd61411,17'd77248,17'd5201,17'd77249,17'd77249,17'd15117,17'd6730,17'd4086,17'd2934,17'd10407,17'd10092,17'd10545,17'd76826,17'd2783,17'd64660,17'd7544,17'd77250,17'd77251,17'd77252,17'd77253,17'd77254,17'd76891,17'd66213,17'd4086,17'd3101,17'd1831,17'd2257,17'd2596,17'd2596,17'd3102,17'd76964,17'd75697,17'd6902,17'd6744,17'd73110,17'd77038,17'd77255,17'd77256,17'd77257,17'd77258,17'd77259,17'd77260,17'd77261,17'd77262,17'd76415,17'd76424,17'd75659,17'd76348,17'd75448,17'd77263,17'd75556,17'd75941,17'd77264,17'd77265,17'd76128,17'd77266,17'd77267,17'd77268,17'd77204,17'd77269,17'd77270,17'd74748,17'd77271,17'd76989,17'd74994,17'd76787,17'd73933,17'd77272,17'd75943,17'd75560,17'd75453,17'd70537,17'd20762,17'd1481,17'd133,17'd133,17'd133,17'd1481,17'd1481,17'd132,17'd11541,17'd131,17'd131,17'd131,17'd131,17'd132,17'd130,17'd136,17'd136,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd77273,17'd4973,17'd6532,17'd3514,17'd77274,17'd77275,17'd77276,17'd77277,17'd77278,17'd13146,17'd77279,17'd77280,17'd77281,17'd77282,17'd77283,17'd33196,17'd77284,17'd77285,17'd77077,17'd15967,17'd76938,17'd77225,17'd14152,17'd76804,17'd76512,17'd76804,17'd77009,17'd77153,17'd77286,17'd14408,17'd77287,17'd15831,17'd77288,17'd77289,17'd6545,17'd6547,17'd5914,17'd5914,17'd6213,17'd6216,17'd8931,17'd7667,17'd5918,17'd5761,17'd76289,17'd52352,17'd6548,17'd6549,17'd6843,17'd6843,17'd75960,17'd76289,17'd50670,17'd50670,17'd27930,17'd27930,17'd5158,17'd5331,17'd5331,17'd5331,17'd5158,17'd5158,17'd5331,17'd5331,17'd28056,17'd28304,17'd6218,17'd6218,17'd5614,17'd37434,17'd6853,17'd6708,17'd6708,17'd6219,17'd6219,17'd6219,17'd9091,17'd7177,17'd7177,17'd7177,17'd6222,17'd6222,17'd6222,17'd6222,17'd6220,17'd6220,17'd6222,17'd6708,17'd6708,17'd6223,17'd6224,17'd6224,17'd6394,17'd8305,17'd8305,17'd8157,17'd8306,17'd9396,17'd10518,17'd9240,17'd11320,17'd8940,17'd19990,17'd11435,17'd11435,17'd8941,17'd34159,17'd9242,17'd77290,17'd5175,17'd4214,17'd4217,17'd3696,17'd6080,17'd8480,17'd51856,17'd51580,17'd57102,17'd77291,17'd1522,17'd77096,17'd77233,17'd77292,17'd578,17'd77293,17'd77294,17'd580,17'd580,17'd77170,17'd77233,17'd77295,17'd578,17'd77174,17'd77296,17'd77297,17'd77298,17'd76469,17'd398,17'd36324,17'd76670,17'd77299,17'd77025,17'd77300,17'd77301,17'd77302,17'd77303,17'd77304,17'd77305,17'd35347,17'd16497,17'd77306,17'd77307,17'd24000,17'd17422,17'd19241,17'd17423,17'd433,17'd620,17'd16634,17'd16634,17'd16633,17'd649,17'd1543,17'd180,17'd27824,17'd254,17'd459,17'd257,17'd270,17'd270,17'd644,17'd645,17'd803,17'd643,17'd643,17'd643
},
'{
17'd3903,17'd3903,17'd3903,17'd4244,17'd15496,17'd3427,17'd3250,17'd3249,17'd2,17'd12,17'd283,17'd650,17'd1830,17'd1688,17'd2422,17'd3250,17'd14,17'd0,17'd283,17'd283,17'd3,17'd12,17'd12,17'd12,17'd12,17'd3,17'd283,17'd1275,17'd1275,17'd2591,17'd2421,17'd7725,17'd977,17'd2591,17'd2933,17'd2591,17'd977,17'd651,17'd465,17'd1275,17'd8814,17'd8814,17'd2933,17'd2933,17'd25,17'd4,17'd8,17'd6,17'd7,17'd7,17'd6,17'd3594,17'd22268,17'd24,17'd5,17'd4,17'd10,17'd10,17'd75696,17'd75696,17'd10,17'd11,17'd20,17'd20,17'd2423,17'd806,17'd21,17'd25,17'd23,17'd4,17'd5,17'd5,17'd5,17'd6,17'd5,17'd24,17'd5,17'd6,17'd8,17'd9,17'd465,17'd283,17'd12,17'd2595,17'd77032,17'd2594,17'd1127,17'd3249,17'd1967,17'd1967,17'd14,17'd14,17'd1127,17'd466,17'd0,17'd1830,17'd1415,17'd17187,17'd14,17'd466,17'd12,17'd650,17'd1830,17'd2422,17'd27441,17'd4888,17'd14745,17'd76828,17'd77249,17'd14598,17'd14598,17'd5203,17'd2934,17'd10545,17'd10407,17'd10546,17'd2593,17'd4738,17'd14598,17'd77308,17'd77309,17'd77310,17'd77311,17'd77310,17'd77312,17'd77313,17'd5959,17'd5203,17'd2784,17'd3250,17'd10268,17'd10268,17'd1693,17'd3102,17'd18037,17'd6744,17'd6902,17'd75697,17'd76964,17'd76394,17'd12197,17'd77314,17'd12784,17'd77315,17'd77316,17'd77317,17'd77318,17'd76489,17'd76975,17'd77319,17'd77320,17'd74869,17'd77321,17'd77322,17'd77322,17'd77323,17'd75660,17'd77324,17'd77325,17'd76696,17'd77128,17'd77326,17'd77327,17'd77328,17'd77329,17'd77330,17'd77331,17'd74513,17'd74296,17'd73502,17'd73826,17'd75451,17'd73828,17'd70537,17'd356,17'd133,17'd133,17'd133,17'd1197,17'd1197,17'd1481,17'd133,17'd132,17'd131,17'd131,17'd131,17'd131,17'd131,17'd132,17'd130,17'd136,17'd136,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd132,17'd132,17'd1759,17'd77332,17'd6369,17'd77333,17'd77334,17'd14695,17'd77209,17'd77335,17'd77336,17'd77337,17'd77212,17'd77338,17'd77339,17'd77340,17'd77341,17'd77342,17'd77343,17'd77344,17'd15966,17'd76937,17'd15708,17'd77345,17'd15455,17'd14284,17'd19981,17'd19981,17'd14549,17'd14549,17'd77346,17'd14701,17'd77347,17'd77348,17'd77349,17'd77289,17'd7324,17'd24650,17'd7008,17'd6212,17'd7166,17'd6846,17'd6214,17'd8931,17'd6552,17'd5761,17'd5915,17'd76289,17'd6548,17'd5149,17'd9368,17'd9368,17'd77350,17'd75960,17'd76289,17'd50670,17'd27930,17'd27930,17'd5158,17'd5331,17'd5332,17'd5332,17'd5158,17'd5158,17'd5158,17'd5331,17'd5613,17'd28056,17'd6389,17'd6389,17'd27935,17'd36887,17'd37434,17'd53214,17'd6853,17'd6853,17'd6390,17'd6390,17'd6708,17'd6708,17'd6708,17'd6708,17'd6222,17'd6222,17'd6222,17'd6222,17'd6708,17'd6708,17'd6708,17'd6223,17'd6223,17'd35760,17'd8630,17'd8473,17'd8473,17'd9395,17'd9395,17'd9239,17'd64502,17'd9784,17'd34795,17'd9658,17'd62682,17'd62682,17'd9935,17'd77351,17'd9936,17'd8005,17'd8942,17'd60617,17'd9787,17'd9243,17'd7510,17'd4705,17'd4862,17'd77352,17'd41158,17'd51183,17'd56665,17'd77353,17'd77354,17'd77355,17'd77356,17'd77357,17'd77358,17'd31725,17'd77359,17'd77360,17'd77361,17'd77170,17'd77233,17'd77172,17'd77362,17'd578,17'd77101,17'd77363,17'd77364,17'd38461,17'd37446,17'd36456,17'd33376,17'd35909,17'd77361,17'd77365,17'd77366,17'd77367,17'd77300,17'd77368,17'd77369,17'd75979,17'd32560,17'd77306,17'd223,17'd280,17'd17423,17'd400,17'd17423,17'd613,17'd463,17'd18515,17'd787,17'd20266,17'd35208,17'd1543,17'd280,17'd20271,17'd278,17'd804,17'd265,17'd268,17'd269,17'd270,17'd644,17'd803,17'd803,17'd643,17'd206,17'd643
},
'{
17'd6264,17'd4428,17'd65576,17'd4427,17'd4087,17'd9960,17'd4088,17'd6096,17'd14,17'd3,17'd806,17'd1275,17'd283,17'd1830,17'd2596,17'd3429,17'd1689,17'd14,17'd0,17'd3,17'd3,17'd806,17'd2423,17'd12,17'd13,17'd3,17'd979,17'd19,17'd11,17'd25,17'd4,17'd5,17'd5206,17'd8,17'd8,17'd4,17'd4,17'd9,17'd9,17'd9,17'd808,17'd10,17'd1275,17'd2933,17'd2933,17'd4242,17'd2421,17'd7373,17'd7,17'd7,17'd6,17'd6,17'd5,17'd5,17'd24,17'd23,17'd23,17'd25,17'd9,17'd25,17'd25,17'd25,17'd22,17'd21,17'd11,17'd11,17'd20,17'd20,17'd22,17'd23,17'd24,17'd5,17'd5,17'd5,17'd5,17'd5,17'd6,17'd6,17'd7,17'd5206,17'd9,17'd25,17'd11,17'd1128,17'd4089,17'd22965,17'd2594,17'd2594,17'd1689,17'd1967,17'd1967,17'd1967,17'd1689,17'd1127,17'd1127,17'd466,17'd1,17'd0,17'd2,17'd466,17'd2,17'd0,17'd1830,17'd64400,17'd6265,17'd77370,17'd77371,17'd77372,17'd5960,17'd72788,17'd77373,17'd77034,17'd15117,17'd13943,17'd2782,17'd7371,17'd10268,17'd10546,17'd12504,17'd66091,17'd77374,17'd77375,17'd77310,17'd77311,17'd77376,17'd77377,17'd77254,17'd77313,17'd14744,17'd4738,17'd63384,17'd77041,17'd293,17'd470,17'd9816,17'd73110,17'd6744,17'd7061,17'd6902,17'd73110,17'd11073,17'd1834,17'd34,17'd77378,17'd77379,17'd77380,17'd77317,17'd77381,17'd77382,17'd77383,17'd77384,17'd77385,17'd77386,17'd77387,17'd77388,17'd77389,17'd77390,17'd77391,17'd76774,17'd77392,17'd76123,17'd77393,17'd77394,17'd76351,17'd76920,17'd75334,17'd74750,17'd75103,17'd77395,17'd73606,17'd73835,17'd73497,17'd71954,17'd138,17'd132,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd3025,17'd77396,17'd5466,17'd18816,17'd77397,17'd77398,17'd77399,17'd77400,17'd77401,17'd77402,17'd77403,17'd77404,17'd77405,17'd77406,17'd77407,17'd77408,17'd77409,17'd77410,17'd77411,17'd77412,17'd77413,17'd77414,17'd77415,17'd15076,17'd77416,17'd77417,17'd77009,17'd20533,17'd77418,17'd14701,17'd77419,17'd77420,17'd77421,17'd77422,17'd38841,17'd8142,17'd8911,17'd7493,17'd62184,17'd25224,17'd7328,17'd6214,17'd6552,17'd27930,17'd76289,17'd50670,17'd5610,17'd4994,17'd6211,17'd6547,17'd5149,17'd6548,17'd4844,17'd5611,17'd5612,17'd5158,17'd5331,17'd5331,17'd5331,17'd5331,17'd6552,17'd6552,17'd5915,17'd50670,17'd5482,17'd5482,17'd5482,17'd5482,17'd5482,17'd5336,17'd5336,17'd5762,17'd5336,17'd5336,17'd5168,17'd37434,17'd37434,17'd37434,17'd37434,17'd37434,17'd5614,17'd5614,17'd5337,17'd5337,17'd5338,17'd35197,17'd35197,17'd35197,17'd52833,17'd52762,17'd52687,17'd5618,17'd5618,17'd6225,17'd5483,17'd34794,17'd9784,17'd5341,17'd5341,17'd4539,17'd5017,17'd5485,17'd4540,17'd4540,17'd4541,17'd5487,17'd77423,17'd9787,17'd6077,17'd4387,17'd3694,17'd4221,17'd54603,17'd77424,17'd51019,17'd77425,17'd77426,17'd55170,17'd53155,17'd25893,17'd77427,17'd31896,17'd576,17'd30941,17'd77428,17'd77293,17'd77429,17'd77101,17'd77430,17'd578,17'd77101,17'd77026,17'd77027,17'd77431,17'd38461,17'd34511,17'd76670,17'd76470,17'd77432,17'd77433,17'd77244,17'd77434,17'd77435,17'd77436,17'd77437,17'd77438,17'd77176,17'd77439,17'd77440,17'd75377,17'd1542,17'd16633,17'd17186,17'd1543,17'd589,17'd214,17'd1116,17'd787,17'd16263,17'd16263,17'd281,17'd1543,17'd20868,17'd20271,17'd27824,17'd804,17'd459,17'd268,17'd269,17'd272,17'd273,17'd273,17'd273,17'd273,17'd272,17'd269
},
'{
17'd4245,17'd3904,17'd9960,17'd4736,17'd9959,17'd4087,17'd9960,17'd6584,17'd1967,17'd0,17'd806,17'd1275,17'd283,17'd1,17'd2936,17'd2258,17'd1689,17'd1967,17'd15,17'd1,17'd3,17'd806,17'd806,17'd12,17'd0,17'd1,17'd1276,17'd1276,17'd979,17'd25,17'd1690,17'd7383,17'd5206,17'd8,17'd8,17'd4,17'd4,17'd4,17'd9,17'd9,17'd808,17'd10,17'd1275,17'd1275,17'd2933,17'd2591,17'd2421,17'd978,17'd7,17'd5205,17'd6,17'd6,17'd6,17'd5,17'd5,17'd24,17'd23,17'd23,17'd23,17'd23,17'd23,17'd23,17'd22,17'd21,17'd11,17'd11,17'd20,17'd20,17'd5518,17'd22,17'd23,17'd24,17'd5,17'd5,17'd5,17'd5,17'd6,17'd6,17'd7,17'd7,17'd8,17'd4,17'd21,17'd20,17'd20404,17'd4089,17'd2595,17'd4247,17'd1688,17'd1689,17'd1967,17'd1967,17'd1689,17'd1688,17'd4247,17'd4247,17'd466,17'd466,17'd466,17'd466,17'd466,17'd14,17'd1830,17'd63118,17'd3750,17'd7371,17'd15496,17'd77441,17'd77442,17'd77443,17'd77444,17'd77111,17'd77036,17'd14744,17'd4086,17'd2783,17'd10546,17'd10545,17'd11072,17'd12504,17'd76958,17'd77445,17'd77446,17'd77447,17'd77448,17'd77448,17'd77449,17'd77450,17'd77451,17'd76958,17'd77033,17'd64793,17'd77107,17'd77452,17'd655,17'd30,17'd29,17'd4430,17'd6744,17'd73110,17'd11073,17'd11209,17'd2427,17'd2120,17'd15629,17'd77453,17'd77454,17'd77455,17'd77456,17'd77457,17'd77458,17'd77459,17'd77460,17'd77461,17'd77462,17'd77463,17'd77464,17'd77465,17'd76491,17'd76494,17'd77466,17'd77467,17'd77124,17'd77060,17'd75449,17'd77468,17'd77469,17'd77470,17'd77471,17'd76042,17'd73929,17'd72872,17'd67858,17'd132,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd1197,17'd77472,17'd77473,17'd19424,17'd19425,17'd77474,17'd77475,17'd76927,17'd77400,17'd77476,17'd77477,17'd77139,17'd77478,17'd77479,17'd14277,17'd77480,17'd77481,17'd77482,17'd77483,17'd15582,17'd77484,17'd77485,17'd77486,17'd77487,17'd77488,17'd77489,17'd14152,17'd20533,17'd77418,17'd22760,17'd77490,17'd13267,17'd24648,17'd38697,17'd45281,17'd77491,17'd8607,17'd23457,17'd8911,17'd7659,17'd7494,17'd6844,17'd50670,17'd5917,17'd5917,17'd5914,17'd5478,17'd5326,17'd26827,17'd26827,17'd5149,17'd6549,17'd5609,17'd4843,17'd4843,17'd5003,17'd5612,17'd5612,17'd5612,17'd5158,17'd5761,17'd6552,17'd5916,17'd5915,17'd5482,17'd5482,17'd5481,17'd5481,17'd5481,17'd5158,17'd5335,17'd5335,17'd5335,17'd5335,17'd5167,17'd5167,17'd5167,17'd36887,17'd36887,17'd36887,17'd28185,17'd28185,17'd36887,17'd51930,17'd35197,17'd35197,17'd52762,17'd52762,17'd34923,17'd34923,17'd77492,17'd77492,17'd35479,17'd63490,17'd63490,17'd5016,17'd62424,17'd6226,17'd77493,17'd4539,17'd35761,17'd6564,17'd6227,17'd6072,17'd77494,17'd4543,17'd5623,17'd6233,17'd77495,17'd77496,17'd4221,17'd77497,17'd55655,17'd77498,17'd77499,17'd77500,17'd55271,17'd54783,17'd33845,17'd77501,17'd77502,17'd77503,17'd31098,17'd31098,17'd575,17'd77504,17'd77362,17'd77237,17'd77504,17'd578,17'd77237,17'd77172,17'd36325,17'd77299,17'd35909,17'd34511,17'd34511,17'd76742,17'd77505,17'd77026,17'd77506,17'd77434,17'd77507,17'd77508,17'd77509,17'd34931,17'd77510,17'd77511,17'd77512,17'd1116,17'd17076,17'd17186,17'd16633,17'd74673,17'd281,17'd1116,17'd20266,17'd29753,17'd76157,17'd30046,17'd1116,17'd24000,17'd252,17'd1826,17'd26728,17'd2255,17'd257,17'd256,17'd269,17'd272,17'd273,17'd272,17'd272,17'd272,17'd270,17'd640
},
'{
17'd4892,17'd3904,17'd4244,17'd7042,17'd4736,17'd5646,17'd9960,17'd4245,17'd2781,17'd15,17'd3,17'd283,17'd283,17'd1412,17'd15,17'd1689,17'd1688,17'd1127,17'd2,17'd3,17'd806,17'd806,17'd3,17'd12,17'd0,17'd0,17'd1277,17'd979,17'd808,17'd25,17'd23,17'd5,17'd5206,17'd8,17'd8,17'd4,17'd4,17'd4,17'd9,17'd9,17'd808,17'd808,17'd1275,17'd1275,17'd2933,17'd2591,17'd2421,17'd7373,17'd3753,17'd5205,17'd5205,17'd5205,17'd6,17'd6,17'd5,17'd5,17'd24,17'd24,17'd23,17'd23,17'd23,17'd23,17'd22,17'd22,17'd21,17'd11,17'd20,17'd20,17'd20,17'd22,17'd23,17'd23,17'd4,17'd4,17'd5,17'd5,17'd6,17'd6,17'd7,17'd7,17'd7,17'd6,17'd4,17'd21,17'd11,17'd18,17'd17,17'd1416,17'd4247,17'd1127,17'd14,17'd14,17'd14,17'd1127,17'd4247,17'd2594,17'd1688,17'd1689,17'd1967,17'd14,17'd1127,17'd4247,17'd14,17'd15,17'd3749,17'd64400,17'd6424,17'd52704,17'd77513,17'd77514,17'd77308,17'd77515,17'd7370,17'd7544,17'd66091,17'd64116,17'd4738,17'd63254,17'd6424,17'd67808,17'd4737,17'd66091,17'd7370,17'd77516,17'd77517,17'd77518,17'd77519,17'd77448,17'd77520,17'd77181,17'd77521,17'd77114,17'd77522,17'd13945,17'd11071,17'd469,17'd31,17'd31,17'd654,17'd3102,17'd76395,17'd77523,17'd77524,17'd77255,17'd76966,17'd58016,17'd77036,17'd77525,17'd77526,17'd77527,17'd77528,17'd77529,17'd77530,17'd77531,17'd77532,17'd77533,17'd77534,17'd76555,17'd77535,17'd76696,17'd76037,17'd77536,17'd77124,17'd77537,17'd77538,17'd75449,17'd74054,17'd75450,17'd76991,17'd75337,17'd73292,17'd71477,17'd136,17'd132,17'd132,17'd134,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd2698,17'd77473,17'd2862,17'd77539,17'd3029,17'd77540,17'd77541,17'd77542,17'd77137,17'd77543,17'd77544,17'd77545,17'd77546,17'd3518,17'd77547,17'd77548,17'd77549,17'd77550,17'd77551,17'd77552,17'd77553,17'd15967,17'd77554,17'd13151,17'd77555,17'd14701,17'd77227,17'd77556,17'd77348,17'd13267,17'd77557,17'd77558,17'd77558,17'd77559,17'd77559,17'd7656,17'd54497,17'd6840,17'd24309,17'd7007,17'd6211,17'd23629,17'd6384,17'd6384,17'd6384,17'd5914,17'd6549,17'd6546,17'd7007,17'd5325,17'd4994,17'd5326,17'd5478,17'd5150,17'd25770,17'd5002,17'd5002,17'd5005,17'd5002,17'd5611,17'd5481,17'd5482,17'd5482,17'd5335,17'd5335,17'd5160,17'd5160,17'd5160,17'd30638,17'd28185,17'd28185,17'd36887,17'd36887,17'd36887,17'd36887,17'd37434,17'd37434,17'd37434,17'd37434,17'd36887,17'd5167,17'd5012,17'd5012,17'd5013,17'd5013,17'd5339,17'd5339,17'd5171,17'd5171,17'd53579,17'd36032,17'd52763,17'd77560,17'd77560,17'd52834,17'd77561,17'd36033,17'd36312,17'd37033,17'd77562,17'd36034,17'd77563,17'd60264,17'd77564,17'd4700,17'd5927,17'd77565,17'd64907,17'd3558,17'd41904,17'd52193,17'd77566,17'd35615,17'd77567,17'd55474,17'd53009,17'd52466,17'd77568,17'd77569,17'd77570,17'd77571,17'd77572,17'd77573,17'd77574,17'd31725,17'd77292,17'd31725,17'd77243,17'd77575,17'd77025,17'd77098,17'd76391,17'd77432,17'd34511,17'd34667,17'd77364,17'd77576,17'd77577,17'd77368,17'd77578,17'd77579,17'd77580,17'd77581,17'd34511,17'd77582,17'd77583,17'd77584,17'd16387,17'd615,17'd74929,17'd18516,17'd20001,17'd435,17'd76157,17'd77585,17'd16006,17'd16140,17'd16263,17'd29173,17'd68847,17'd648,17'd180,17'd17422,17'd18387,17'd460,17'd263,17'd262,17'd270,17'd272,17'd272,17'd272,17'd270,17'd270,17'd268,17'd256
},
'{
17'd27713,17'd3903,17'd3903,17'd77586,17'd4736,17'd4891,17'd4892,17'd6420,17'd3250,17'd1967,17'd0,17'd1,17'd1412,17'd1412,17'd1,17'd14,17'd1688,17'd1689,17'd14,17'd0,17'd3,17'd1275,17'd3,17'd3,17'd0,17'd2,17'd16,17'd1276,17'd3748,17'd21,17'd23,17'd5,17'd8,17'd8,17'd8,17'd8,17'd4,17'd4,17'd9,17'd9,17'd808,17'd808,17'd1275,17'd1275,17'd2591,17'd2591,17'd2421,17'd7215,17'd3753,17'd3753,17'd5205,17'd5205,17'd7,17'd6,17'd6,17'd5,17'd24,17'd24,17'd23,17'd23,17'd23,17'd23,17'd23,17'd23,17'd21,17'd10,17'd20,17'd2598,17'd2598,17'd20,17'd21,17'd22,17'd4,17'd4,17'd4,17'd5,17'd6,17'd6,17'd6,17'd6,17'd7,17'd7,17'd8,17'd4,17'd21,17'd11,17'd18,17'd16,17'd466,17'd14,17'd14,17'd14,17'd14,17'd1127,17'd4247,17'd4247,17'd3252,17'd2422,17'd2781,17'd1967,17'd1689,17'd4247,17'd4247,17'd15745,17'd15,17'd1967,17'd6265,17'd63255,17'd64116,17'd77587,17'd77588,17'd77589,17'd77308,17'd77313,17'd8337,17'd76827,17'd66091,17'd4893,17'd14071,17'd67808,17'd63384,17'd4737,17'd5645,17'd7047,17'd77110,17'd77590,17'd77591,17'd77592,17'd77593,17'd77594,17'd77447,17'd77312,17'd8337,17'd76828,17'd4737,17'd3751,17'd2782,17'd76826,17'd10545,17'd10407,17'd10267,17'd77523,17'd77523,17'd77523,17'd1834,17'd77255,17'd77041,17'd13944,17'd77595,17'd77596,17'd77597,17'd77598,17'd77599,17'd77600,17'd76332,17'd76334,17'd77533,17'd77601,17'd76342,17'd77602,17'd77603,17'd77604,17'd77605,17'd77606,17'd75941,17'd76041,17'd75450,17'd73608,17'd74404,17'd73078,17'd72552,17'd20762,17'd130,17'd132,17'd130,17'd128,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd135,17'd76571,17'd2862,17'd6532,17'd19425,17'd77607,17'd77608,17'd77609,17'd19297,17'd19048,17'd77335,17'd77610,17'd77546,17'd77611,17'd14947,17'd77612,17'd77613,17'd77614,17'd36880,17'd77615,17'd77616,17'd76937,17'd16704,17'd77617,17'd13151,17'd15076,17'd16227,17'd77618,17'd77619,17'd77557,17'd12739,17'd13019,17'd13388,17'd8758,17'd9066,17'd77491,17'd8142,17'd54497,17'd7005,17'd77620,17'd7007,17'd23799,17'd6212,17'd5913,17'd6384,17'd5915,17'd5913,17'd6547,17'd7007,17'd77621,17'd5324,17'd4994,17'd5326,17'd5478,17'd5150,17'd4845,17'd5002,17'd5005,17'd5005,17'd4843,17'd4843,17'd4843,17'd4843,17'd25627,17'd5004,17'd25627,17'd25627,17'd25627,17'd30638,17'd30638,17'd28185,17'd36887,17'd36887,17'd36887,17'd37434,17'd37434,17'd53214,17'd53214,17'd37434,17'd5167,17'd5167,17'd5012,17'd5011,17'd37697,17'd37697,17'd52603,17'd52603,17'd37945,17'd77622,17'd52095,17'd52095,17'd38192,17'd52522,17'd52522,17'd57868,17'd57868,17'd52907,17'd37561,17'd37700,17'd77623,17'd77624,17'd6073,17'd6229,17'd5925,17'd77625,17'd77565,17'd64777,17'd3558,17'd46238,17'd64644,17'd50592,17'd57360,17'd77626,17'd53747,17'd53518,17'd77627,17'd77628,17'd77569,17'd77629,17'd77571,17'd77630,17'd77631,17'd77632,17'd77633,17'd576,17'd77634,17'd77244,17'd77243,17'd77575,17'd395,17'd77098,17'd77096,17'd77432,17'd77094,17'd34345,17'd77635,17'd77636,17'd77637,17'd77638,17'd77639,17'd77640,17'd77641,17'd28655,17'd77642,17'd28191,17'd222,17'd77585,17'd30046,17'd30046,17'd18633,17'd33539,17'd32559,17'd619,17'd15874,17'd32407,17'd77643,17'd75379,17'd588,17'd39950,17'd77644,17'd24332,17'd401,17'd402,17'd804,17'd255,17'd262,17'd262,17'd269,17'd270,17'd272,17'd270,17'd269,17'd269,17'd257,17'd262
},
'{
17'd4244,17'd3902,17'd65576,17'd9960,17'd3903,17'd3903,17'd27713,17'd25384,17'd2935,17'd3250,17'd3249,17'd1830,17'd1,17'd1412,17'd1,17'd0,17'd4247,17'd1127,17'd466,17'd0,17'd3,17'd3,17'd3,17'd3,17'd1,17'd2,17'd16,17'd979,17'd10,17'd21,17'd23,17'd4,17'd8,17'd8,17'd6,17'd6,17'd6,17'd5,17'd4,17'd4,17'd9,17'd25,17'd25,17'd25,17'd23,17'd23,17'd7215,17'd7215,17'd3753,17'd3753,17'd5205,17'd5205,17'd7,17'd7,17'd6,17'd6,17'd5,17'd24,17'd24,17'd24,17'd23,17'd23,17'd23,17'd23,17'd25,17'd21,17'd20,17'd20,17'd1128,17'd11,17'd11,17'd21,17'd25,17'd23,17'd4,17'd4,17'd6,17'd6,17'd3753,17'd3753,17'd5205,17'd5205,17'd6,17'd4,17'd23,17'd21,17'd11,17'd19,17'd18,17'd16,17'd16,17'd17,17'd17,17'd17,17'd17,17'd1415,17'd14070,17'd14070,17'd3252,17'd1831,17'd1689,17'd1127,17'd1127,17'd4247,17'd17917,17'd1689,17'd9815,17'd68191,17'd63384,17'd14443,17'd67065,17'd77645,17'd77646,17'd77250,17'd77521,17'd77313,17'd8337,17'd5959,17'd64392,17'd4737,17'd76957,17'd14071,17'd3903,17'd5201,17'd7544,17'd77516,17'd77590,17'd77647,17'd77648,17'd77649,17'd77650,17'd77519,17'd77651,17'd77652,17'd72788,17'd5645,17'd71304,17'd64251,17'd76957,17'd76826,17'd10545,17'd10545,17'd10092,17'd655,17'd77523,17'd11208,17'd469,17'd32,17'd12505,17'd14072,17'd77653,17'd77654,17'd77655,17'd77656,17'd77657,17'd77658,17'd77659,17'd77660,17'd77661,17'd77662,17'd77663,17'd77664,17'd76502,17'd75663,17'd77665,17'd77666,17'd73829,17'd73929,17'd75668,17'd71477,17'd1481,17'd134,17'd134,17'd132,17'd130,17'd128,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd10492,17'd3812,17'd6369,17'd20059,17'd18817,17'd19169,17'd77667,17'd77609,17'd77668,17'd77669,17'd77335,17'd77670,17'd77671,17'd77672,17'd77673,17'd31238,17'd9365,17'd33033,17'd77674,17'd77675,17'd77676,17'd77677,17'd77678,17'd77679,17'd77617,17'd13390,17'd77680,17'd77681,17'd77682,17'd77683,17'd77684,17'd16463,17'd32716,17'd32238,17'd8758,17'd6542,17'd77685,17'd4520,17'd4186,17'd53056,17'd5322,17'd24944,17'd23629,17'd6384,17'd50670,17'd5914,17'd31088,17'd5608,17'd24649,17'd24649,17'd24649,17'd5323,17'd4840,17'd4688,17'd4688,17'd4845,17'd4845,17'd4845,17'd4687,17'd4686,17'd4842,17'd28418,17'd28418,17'd28418,17'd28418,17'd28418,17'd4842,17'd4842,17'd5005,17'd30637,17'd5004,17'd25627,17'd5163,17'd5163,17'd5163,17'd37030,17'd37030,17'd37030,17'd77686,17'd56308,17'd77687,17'd77687,17'd50835,17'd50835,17'd50918,17'd50918,17'd50488,17'd50488,17'd50488,17'd51248,17'd51248,17'd51177,17'd51177,17'd51177,17'd38445,17'd56203,17'd77688,17'd77689,17'd60388,17'd7335,17'd35054,17'd77690,17'd63500,17'd19859,17'd49107,17'd3208,17'd45514,17'd52533,17'd50592,17'd77691,17'd77692,17'd77693,17'd53071,17'd77501,17'd77628,17'd26720,17'd77694,17'd77695,17'd77695,17'd77696,17'd77697,17'd392,17'd77698,17'd77699,17'd576,17'd77700,17'd77701,17'd77243,17'd77292,17'd77233,17'd77702,17'd77094,17'd36750,17'd77703,17'd77704,17'd77705,17'd77706,17'd77707,17'd77708,17'd37045,17'd1235,17'd926,17'd51582,17'd767,17'd76310,17'd16263,17'd618,17'd52197,17'd52107,17'd788,17'd75253,17'd77709,17'd31412,17'd76745,17'd77643,17'd16635,17'd77710,17'd77711,17'd23489,17'd17423,17'd19241,17'd180,17'd20009,17'd456,17'd265,17'd256,17'd968,17'd1407,17'd1407,17'd1407,17'd268,17'd268,17'd263,17'd459
},
'{
17'd7042,17'd3902,17'd65576,17'd9960,17'd3903,17'd9960,17'd27590,17'd4243,17'd3427,17'd2784,17'd2781,17'd3249,17'd1830,17'd1412,17'd283,17'd3,17'd14,17'd1127,17'd466,17'd2,17'd12,17'd3,17'd3,17'd3,17'd1,17'd0,17'd16,17'd16,17'd19,17'd10,17'd25,17'd4,17'd8,17'd8,17'd6,17'd6,17'd6,17'd6,17'd4,17'd4,17'd9,17'd9,17'd25,17'd25,17'd23,17'd23,17'd7215,17'd7215,17'd3753,17'd3753,17'd5205,17'd5205,17'd7,17'd7,17'd7,17'd6,17'd5,17'd5,17'd5,17'd24,17'd23,17'd23,17'd23,17'd23,17'd25,17'd25,17'd21,17'd20,17'd11,17'd1128,17'd11,17'd11,17'd10,17'd25,17'd25,17'd4,17'd6,17'd6,17'd3753,17'd3753,17'd3753,17'd3753,17'd6,17'd6,17'd4,17'd23,17'd21,17'd11,17'd10,17'd19,17'd19,17'd16,17'd16,17'd16,17'd16,17'd17187,17'd1689,17'd2422,17'd3252,17'd10535,17'd1831,17'd1688,17'd1689,17'd1688,17'd1831,17'd1688,17'd3250,17'd2784,17'd75260,17'd63385,17'd64251,17'd6263,17'd77712,17'd30947,17'd77713,17'd77714,17'd77521,17'd77313,17'd76892,17'd76958,17'd64116,17'd14071,17'd6892,17'd4736,17'd5376,17'd77373,17'd77521,17'd77252,17'd77715,17'd77716,17'd77648,17'd77717,17'd77718,17'd77719,17'd77720,17'd8509,17'd7541,17'd70486,17'd69718,17'd4738,17'd2783,17'd2593,17'd10669,17'd3593,17'd33,17'd293,17'd293,17'd11071,17'd16501,17'd77721,17'd63670,17'd77722,17'd76681,17'd77723,17'd77724,17'd76549,17'd77725,17'd77726,17'd77727,17'd77728,17'd77729,17'd77730,17'd77606,17'd75941,17'd77731,17'd76042,17'd77732,17'd73602,17'd71477,17'd20762,17'd132,17'd131,17'd132,17'd132,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd357,17'd4814,17'd77733,17'd77734,17'd77735,17'd5595,17'd77736,17'd77737,17'd19297,17'd77137,17'd18933,17'd77476,17'd77738,17'd77739,17'd77740,17'd77741,17'd77742,17'd77743,17'd77744,17'd77745,17'd77746,17'd32072,17'd42768,17'd61391,17'd61391,17'd77747,17'd15583,17'd77748,17'd77749,17'd77750,17'd32716,17'd77751,17'd11420,17'd77752,17'd77753,17'd11983,17'd77754,17'd8141,17'd5911,17'd33041,17'd53278,17'd24795,17'd26827,17'd5914,17'd6384,17'd5914,17'd25225,17'd25628,17'd24944,17'd4992,17'd24798,17'd53352,17'd42910,17'd32552,17'd4840,17'd32552,17'd4688,17'd4687,17'd4687,17'd4686,17'd4686,17'd4686,17'd4841,17'd4841,17'd4841,17'd4841,17'd4841,17'd4841,17'd4841,17'd28418,17'd28418,17'd28418,17'd37153,17'd37153,17'd37153,17'd29024,17'd37288,17'd37288,17'd38567,17'd4528,17'd50488,17'd50488,17'd50488,17'd50488,17'd50488,17'd50488,17'd4528,17'd4527,17'd50587,17'd55457,17'd52011,17'd51010,17'd51010,17'd52688,17'd56203,17'd38322,17'd37809,17'd77755,17'd77756,17'd35200,17'd77757,17'd77758,17'd3548,17'd77759,17'd42646,17'd41770,17'd2893,17'd63103,17'd62844,17'd77760,17'd77761,17'd77762,17'd77568,17'd77763,17'd77764,17'd77765,17'd77766,17'd77767,17'd387,17'd77768,17'd77769,17'd77696,17'd77770,17'd77633,17'd77574,17'd77771,17'd77701,17'd77701,17'd77292,17'd77772,17'd77773,17'd77170,17'd77233,17'd77774,17'd77775,17'd77776,17'd77777,17'd77778,17'd36182,17'd77779,17'd77780,17'd18759,17'd51496,17'd16263,17'd16005,17'd16005,17'd16497,17'd219,17'd38335,17'd76073,17'd52023,17'd76233,17'd32883,17'd586,17'd16263,17'd769,17'd77711,17'd280,17'd400,17'd17423,17'd251,17'd964,17'd2420,17'd804,17'd265,17'd257,17'd74675,17'd968,17'd1407,17'd268,17'd268,17'd257,17'd459,17'd969
},
'{
17'd77781,17'd10533,17'd47270,17'd77781,17'd9960,17'd9960,17'd3902,17'd4891,17'd4892,17'd4088,17'd6424,17'd3750,17'd3249,17'd1,17'd1275,17'd806,17'd0,17'd14,17'd466,17'd466,17'd12,17'd3,17'd1,17'd1,17'd1,17'd1,17'd0,17'd13,17'd1128,17'd10,17'd25,17'd23,17'd4,17'd5,17'd6,17'd6,17'd6,17'd6,17'd8,17'd8,17'd9,17'd9,17'd9,17'd25,17'd23,17'd4,17'd5,17'd5,17'd3753,17'd3753,17'd3753,17'd5205,17'd5205,17'd5205,17'd5205,17'd5205,17'd6,17'd5,17'd5,17'd24,17'd24,17'd24,17'd23,17'd4,17'd25,17'd25,17'd21,17'd21,17'd11,17'd1128,17'd18,17'd1128,17'd10,17'd21,17'd25,17'd4,17'd5,17'd6,17'd3594,17'd3594,17'd3753,17'd3753,17'd5205,17'd3753,17'd6,17'd4,17'd23,17'd21,17'd25,17'd10,17'd11,17'd19,17'd19,17'd19,17'd19,17'd16,17'd9422,17'd17187,17'd1127,17'd1831,17'd1831,17'd2422,17'd2422,17'd1831,17'd1689,17'd3250,17'd3252,17'd3252,17'd2784,17'd7371,17'd6424,17'd14071,17'd5052,17'd77782,17'd31256,17'd77720,17'd77783,17'd77309,17'd77714,17'd77313,17'd7544,17'd5376,17'd69718,17'd69718,17'd7212,17'd70486,17'd77373,17'd77784,17'd77785,17'd77717,17'd77786,17'd77787,17'd77788,17'd77789,17'd77790,17'd77791,17'd77792,17'd7370,17'd5960,17'd5201,17'd6730,17'd4086,17'd16392,17'd14320,17'd14989,17'd14190,17'd14321,17'd14322,17'd63670,17'd77793,17'd77794,17'd77795,17'd77796,17'd77797,17'd77798,17'd77799,17'd77800,17'd77801,17'd77802,17'd77803,17'd76981,17'd77729,17'd77804,17'd77805,17'd74403,17'd73610,17'd77806,17'd72655,17'd137,17'd128,17'd134,17'd132,17'd132,17'd132,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd76993,17'd3169,17'd77807,17'd77808,17'd77809,17'd3172,17'd77810,17'd77811,17'd19297,17'd77137,17'd77812,17'd77813,17'd77814,17'd77815,17'd77816,17'd9497,17'd77817,17'd77818,17'd77819,17'd31395,17'd77820,17'd24145,17'd12134,17'd58481,17'd77821,17'd77822,17'd15829,17'd77823,17'd77824,17'd77825,17'd41885,17'd77826,17'd77827,17'd37146,17'd6377,17'd77828,17'd4986,17'd5142,17'd4363,17'd4521,17'd38441,17'd77829,17'd4993,17'd6382,17'd6382,17'd25225,17'd31088,17'd5479,17'd5326,17'd5325,17'd77621,17'd53352,17'd53352,17'd5145,17'd6067,17'd4682,17'd4683,17'd4683,17'd4683,17'd4840,17'd32552,17'd44614,17'd44614,17'd39166,17'd5757,17'd4840,17'd4840,17'd4840,17'd4840,17'd4683,17'd5328,17'd5328,17'd5328,17'd5328,17'd5328,17'd5328,17'd4684,17'd49995,17'd49995,17'd49995,17'd4527,17'd4527,17'd4527,17'd4527,17'd4527,17'd4690,17'd4690,17'd49896,17'd4371,17'd51327,17'd50836,17'd38322,17'd77830,17'd38448,17'd58974,17'd77831,17'd77832,17'd77833,17'd77834,17'd77835,17'd77836,17'd2884,17'd2536,17'd77837,17'd2729,17'd37166,17'd77838,17'd77839,17'd53155,17'd77840,17'd77841,17'd77842,17'd77843,17'd77844,17'd77845,17'd77846,17'd28542,17'd77847,17'd77847,17'd77848,17'd77696,17'd77631,17'd77631,17'd77633,17'd77771,17'd77849,17'd77850,17'd577,17'd77851,17'd77851,17'd77237,17'd77237,17'd77026,17'd77103,17'd37447,17'd77305,17'd76235,17'd77852,17'd77853,17'd77854,17'd76604,17'd32726,17'd36046,17'd75691,17'd35617,17'd16497,17'd586,17'd31730,17'd77024,17'd76233,17'd31730,17'd586,17'd29753,17'd35208,17'd51335,17'd280,17'd19363,17'd76312,17'd614,17'd638,17'd612,17'd639,17'd804,17'd265,17'd266,17'd262,17'd257,17'd268,17'd268,17'd263,17'd801,17'd254,17'd965
},
'{
17'd33216,17'd30047,17'd4889,17'd47270,17'd65576,17'd3903,17'd9960,17'd3902,17'd3902,17'd9960,17'd67808,17'd7371,17'd3249,17'd1,17'd1275,17'd806,17'd1,17'd15,17'd466,17'd466,17'd13,17'd3,17'd1,17'd1,17'd1,17'd1,17'd0,17'd466,17'd3905,17'd10,17'd808,17'd25,17'd4,17'd5,17'd6,17'd6,17'd6,17'd6,17'd8,17'd8,17'd1413,17'd9,17'd9,17'd9,17'd4,17'd4,17'd5,17'd5,17'd3753,17'd3753,17'd3753,17'd3753,17'd5205,17'd5205,17'd5205,17'd5205,17'd6,17'd6,17'd5,17'd5,17'd24,17'd24,17'd23,17'd4,17'd25,17'd25,17'd25,17'd21,17'd11,17'd11,17'd18,17'd3905,17'd10,17'd10,17'd808,17'd9,17'd4,17'd5,17'd5,17'd3594,17'd3753,17'd3753,17'd5205,17'd5205,17'd6,17'd5,17'd23,17'd23,17'd21,17'd21,17'd10,17'd10,17'd10,17'd979,17'd18,17'd3905,17'd18,17'd16,17'd0,17'd14,17'd1689,17'd3250,17'd2422,17'd2422,17'd3250,17'd2781,17'd2781,17'd14070,17'd14188,17'd14070,17'd2422,17'd4887,17'd77855,17'd5644,17'd77856,17'd30947,17'd77181,17'd77783,17'd77309,17'd77714,17'd77451,17'd77857,17'd5374,17'd70486,17'd77858,17'd77859,17'd5792,17'd77443,17'd77860,17'd77861,17'd77718,17'd77862,17'd77863,17'd77788,17'd77864,17'd77865,17'd77866,17'd8189,17'd77313,17'd6261,17'd5960,17'd14598,17'd14598,17'd76828,17'd77184,17'd77374,17'd76891,17'd77308,17'd77182,17'd77520,17'd77867,17'd77868,17'd77869,17'd77870,17'd77871,17'd77872,17'd77873,17'd77874,17'd77875,17'd77876,17'd77877,17'd77121,17'd75849,17'd75851,17'd74755,17'd73602,17'd71954,17'd67858,17'd136,17'd128,17'd128,17'd132,17'd132,17'd1759,17'd1197,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd132,17'd5898,17'd6055,17'd3812,17'd77734,17'd77878,17'd5595,17'd77879,17'd76132,17'd77209,17'd77880,17'd77813,17'd77881,17'd77813,17'd77882,17'd77883,17'd14696,17'd77884,17'd77885,17'd31240,17'd77819,17'd77886,17'd77887,17'd77888,17'd77889,17'd77889,17'd77890,17'd77616,17'd10881,17'd13389,17'd6208,17'd77891,17'd77892,17'd36577,17'd39005,17'd10357,17'd77893,17'd39462,17'd4986,17'd33531,17'd33205,17'd4522,17'd53280,17'd53056,17'd7324,17'd23975,17'd31088,17'd5478,17'd5326,17'd5479,17'd31088,17'd4993,17'd77894,17'd77895,17'd4997,17'd38442,17'd5144,17'd5144,17'd5145,17'd42910,17'd4995,17'd4839,17'd34156,17'd34156,17'd5606,17'd5606,17'd4839,17'd5757,17'd5757,17'd5757,17'd4840,17'd4840,17'd4840,17'd4840,17'd4840,17'd4840,17'd4840,17'd4683,17'd4684,17'd4527,17'd4527,17'd49995,17'd49995,17'd49995,17'd49995,17'd58971,17'd57867,17'd57867,17'd49805,17'd51403,17'd77896,17'd38448,17'd58352,17'd59746,17'd4033,17'd59747,17'd59748,17'd60141,17'd77897,17'd64096,17'd48470,17'd77898,17'd51015,17'd77899,17'd37571,17'd77900,17'd57607,17'd77901,17'd53155,17'd77902,17'd77903,17'd77904,17'd77843,17'd77905,17'd1081,17'd77906,17'd77907,17'd77847,17'd77847,17'd77908,17'd77909,17'd77910,17'd77911,17'd77912,17'd77913,17'd77633,17'd77914,17'd77915,17'd577,17'd77916,17'd77917,17'd77244,17'd77918,17'd77237,17'd37170,17'd76391,17'd77919,17'd77920,17'd77921,17'd77853,17'd586,17'd16388,17'd76675,17'd76675,17'd32883,17'd586,17'd35617,17'd16388,17'd77922,17'd37446,17'd33214,17'd76233,17'd76604,17'd76232,17'd1238,17'd613,17'd77923,17'd75982,17'd20001,17'd35208,17'd280,17'd638,17'd182,17'd1095,17'd595,17'd265,17'd262,17'd256,17'd268,17'd967,17'd801,17'd460,17'd804,17'd26728
},
'{
17'd6421,17'd5199,17'd30047,17'd47270,17'd4244,17'd3903,17'd3903,17'd9960,17'd4087,17'd4244,17'd3751,17'd6424,17'd9815,17'd1830,17'd283,17'd3,17'd1,17'd1830,17'd0,17'd2,17'd2,17'd2,17'd0,17'd1,17'd1,17'd1,17'd1,17'd0,17'd18,17'd11,17'd10,17'd9,17'd4,17'd5,17'd6,17'd6,17'd6,17'd6,17'd6,17'd6,17'd4,17'd4,17'd9,17'd9,17'd4,17'd4,17'd5,17'd5,17'd6,17'd6,17'd6,17'd6,17'd3753,17'd3753,17'd5205,17'd8190,17'd5205,17'd3753,17'd24,17'd24,17'd24,17'd24,17'd23,17'd23,17'd4,17'd4,17'd25,17'd25,17'd10,17'd11,17'd18,17'd18,17'd18,17'd1128,17'd11,17'd21,17'd2591,17'd2421,17'd2421,17'd16009,17'd6,17'd6,17'd6,17'd7,17'd7,17'd6,17'd5,17'd284,17'd22,17'd22,17'd25,17'd25,17'd25,17'd10,17'd10,17'd11,17'd1128,17'd1128,17'd18,17'd16,17'd1415,17'd2936,17'd1689,17'd1689,17'd1831,17'd1689,17'd1967,17'd1689,17'd1831,17'd77924,17'd77924,17'd3252,17'd25384,17'd77925,17'd77926,17'd7368,17'd77180,17'd77927,17'd77446,17'd77446,17'd77446,17'd77312,17'd77451,17'd8337,17'd72788,17'd73013,17'd73013,17'd70486,17'd8337,17'd77928,17'd77929,17'd77310,17'd77930,17'd77931,17'd77788,17'd77932,17'd77933,17'd77934,17'd77935,17'd77652,17'd77936,17'd76892,17'd76892,17'd77453,17'd77183,17'd77521,17'd77182,17'd77783,17'd77937,17'd77938,17'd77939,17'd77649,17'd76482,17'd76686,17'd76687,17'd77940,17'd77941,17'd77942,17'd77943,17'd77944,17'd77945,17'd75938,17'd77946,17'd74518,17'd77947,17'd71260,17'd71260,17'd71372,17'd71477,17'd141,17'd129,17'd132,17'd132,17'd131,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd77948,17'd4336,17'd77949,17'd3513,17'd77950,17'd3030,17'd77951,17'd3515,17'd77952,17'd77953,17'd77881,17'd77954,17'd77955,17'd12598,17'd77956,17'd77957,17'd3823,17'd77958,17'd11419,17'd77959,17'd37548,17'd77960,17'd9763,17'd77961,17'd11690,17'd12279,17'd8288,17'd8910,17'd8758,17'd77962,17'd77963,17'd77964,17'd77965,17'd77966,17'd77967,17'd6205,17'd6539,17'd39462,17'd77968,17'd34920,17'd33205,17'd4520,17'd54497,17'd5322,17'd4994,17'd5478,17'd5478,17'd5609,17'd31088,17'd31088,17'd5608,17'd24649,17'd77969,17'd77970,17'd77971,17'd77972,17'd4188,17'd4838,17'd4991,17'd4188,17'd4838,17'd4676,17'd4837,17'd4837,17'd4681,17'd4681,17'd24649,17'd5323,17'd5323,17'd4992,17'd4839,17'd5757,17'd5757,17'd5757,17'd5757,17'd5757,17'd5156,17'd5156,17'd4689,17'd5156,17'd4690,17'd58971,17'd57867,17'd49598,17'd49805,17'd54499,17'd53860,17'd38572,17'd58352,17'd59746,17'd36738,17'd49402,17'd77973,17'd77974,17'd77975,17'd63502,17'd3049,17'd77976,17'd51407,17'd2374,17'd52696,17'd2547,17'd2548,17'd36321,17'd77977,17'd54518,17'd77978,17'd77979,17'd77980,17'd77981,17'd77982,17'd77983,17'd77984,17'd26336,17'd163,17'd77985,17'd77986,17'd77987,17'd77988,17'd77989,17'd77911,17'd77990,17'd77770,17'd77991,17'd77915,17'd77992,17'd77701,17'd77993,17'd77300,17'd77302,17'd77102,17'd77022,17'd37045,17'd52367,17'd77994,17'd77995,17'd28313,17'd32883,17'd77996,17'd77997,17'd76606,17'd76156,17'd76469,17'd75376,17'd36046,17'd32883,17'd176,17'd77998,17'd36046,17'd220,17'd77999,17'd78000,17'd78001,17'd78002,17'd464,17'd281,17'd1116,17'd620,17'd280,17'd213,17'd639,17'd17551,17'd595,17'd2255,17'd459,17'd265,17'd967,17'd2588,17'd460,17'd253,17'd639,17'd401
},
'{
17'd5510,17'd5790,17'd33216,17'd30047,17'd4427,17'd4244,17'd3903,17'd9960,17'd4427,17'd4427,17'd13943,17'd2782,17'd2781,17'd15,17'd3,17'd3,17'd1,17'd1830,17'd0,17'd0,17'd2,17'd2,17'd0,17'd1,17'd1,17'd1,17'd1,17'd1,17'd18,17'd19,17'd10,17'd25,17'd23,17'd5,17'd5,17'd6,17'd6,17'd6,17'd6,17'd6,17'd4,17'd4,17'd9,17'd9,17'd4,17'd4,17'd5,17'd5,17'd6,17'd6,17'd6,17'd6,17'd3753,17'd3753,17'd5205,17'd5205,17'd5205,17'd3753,17'd5,17'd24,17'd24,17'd24,17'd23,17'd23,17'd23,17'd23,17'd25,17'd25,17'd10,17'd11,17'd19,17'd18,17'd4089,17'd3905,17'd11,17'd10,17'd465,17'd2591,17'd977,17'd2421,17'd4,17'd5,17'd6,17'd6,17'd7,17'd7,17'd6,17'd5,17'd23,17'd23,17'd25,17'd25,17'd25,17'd21,17'd10,17'd10,17'd20,17'd20,17'd11,17'd19,17'd1277,17'd16,17'd15,17'd15,17'd1127,17'd1127,17'd1127,17'd1127,17'd4247,17'd2594,17'd17917,17'd27714,17'd14743,17'd78003,17'd77925,17'd5199,17'd7047,17'd77589,17'd77927,17'd78004,17'd77446,17'd77446,17'd77713,17'd77110,17'd77308,17'd6261,17'd70486,17'd77858,17'd7212,17'd5960,17'd77928,17'd78005,17'd77866,17'd77592,17'd78006,17'd78007,17'd78008,17'd78009,17'd77448,17'd77866,17'd77309,17'd77254,17'd78010,17'd78011,17'd78012,17'd77714,17'd77783,17'd77791,17'd78013,17'd78014,17'd78015,17'd78016,17'd78017,17'd78018,17'd78019,17'd78020,17'd78021,17'd78022,17'd78023,17'd78024,17'd76699,17'd78025,17'd78026,17'd78027,17'd73395,17'd70742,17'd72757,17'd71477,17'd78028,17'd141,17'd130,17'd132,17'd131,17'd131,17'd133,17'd133,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd52246,17'd76993,17'd78029,17'd77734,17'd12876,17'd13383,17'd78030,17'd78031,17'd18213,17'd77952,17'd78032,17'd78033,17'd77137,17'd78034,17'd78035,17'd78036,17'd9210,17'd78037,17'd78038,17'd78039,17'd78040,17'd8138,17'd31395,17'd78041,17'd77826,17'd78042,17'd6837,17'd7160,17'd12279,17'd32398,17'd35467,17'd37280,17'd78043,17'd8284,17'd77966,17'd46981,17'd78044,17'd77893,17'd78045,17'd78046,17'd10195,17'd36730,17'd4989,17'd53280,17'd77969,17'd5146,17'd4993,17'd4994,17'd4994,17'd24944,17'd24944,17'd25083,17'd5608,17'd4992,17'd5322,17'd52761,17'd38846,17'd38846,17'd4187,17'd33367,17'd38846,17'd38846,17'd4187,17'd4187,17'd33367,17'd4997,17'd77969,17'd77969,17'd24649,17'd24649,17'd6067,17'd6067,17'd6067,17'd6067,17'd6067,17'd4525,17'd4525,17'd41459,17'd49804,17'd49496,17'd55351,17'd55351,17'd52183,17'd51489,17'd51664,17'd52605,17'd38061,17'd4204,17'd3847,17'd78047,17'd36038,17'd60503,17'd77975,17'd78048,17'd3049,17'd64908,17'd44741,17'd2539,17'd40407,17'd52458,17'd59495,17'd78049,17'd36321,17'd78050,17'd78051,17'd78052,17'd78053,17'd78054,17'd78055,17'd26226,17'd78056,17'd78057,17'd78058,17'd78059,17'd163,17'd78060,17'd77987,17'd78061,17'd386,17'd78062,17'd77911,17'd77631,17'd77912,17'd77573,17'd78063,17'd78064,17'd77242,17'd77993,17'd77302,17'd77701,17'd77025,17'd77021,17'd27821,17'd1235,17'd26721,17'd51858,17'd76672,17'd398,17'd78065,17'd76744,17'd78066,17'd76817,17'd75980,17'd31255,17'd33214,17'd76532,17'd176,17'd78067,17'd32883,17'd31412,17'd78068,17'd76238,17'd437,17'd78069,17'd75253,17'd20266,17'd75256,17'd35208,17'd770,17'd251,17'd639,17'd181,17'd254,17'd2255,17'd265,17'd801,17'd801,17'd1095,17'd253,17'd20271,17'd15492,17'd78070
},
'{
17'd5375,17'd6422,17'd5644,17'd33216,17'd30047,17'd47270,17'd4736,17'd4736,17'd4736,17'd4427,17'd4244,17'd4088,17'd2592,17'd1967,17'd0,17'd0,17'd1412,17'd1,17'd1,17'd0,17'd2,17'd2,17'd0,17'd1,17'd1,17'd1412,17'd283,17'd283,17'd3,17'd3,17'd11,17'd21,17'd23,17'd4,17'd5,17'd6,17'd6,17'd6,17'd6,17'd6,17'd4,17'd4,17'd9,17'd9,17'd4,17'd4,17'd4,17'd4,17'd6,17'd6,17'd6,17'd6,17'd6,17'd6,17'd5205,17'd5205,17'd5205,17'd5205,17'd6,17'd5,17'd5,17'd24,17'd4,17'd4,17'd23,17'd23,17'd25,17'd25,17'd21,17'd21,17'd11,17'd11,17'd4089,17'd4089,17'd13,17'd2423,17'd1275,17'd465,17'd651,17'd2591,17'd4,17'd4,17'd4,17'd8,17'd6,17'd6,17'd6,17'd6,17'd5,17'd5,17'd23,17'd23,17'd23,17'd23,17'd25,17'd25,17'd21,17'd21,17'd10,17'd10,17'd979,17'd979,17'd10,17'd10,17'd2423,17'd12,17'd13,17'd2,17'd1127,17'd1127,17'd1831,17'd3252,17'd14743,17'd6420,17'd4428,17'd9960,17'd69718,17'd5960,17'd78071,17'd78072,17'd77927,17'd77181,17'd77713,17'd77312,17'd77110,17'd77451,17'd8337,17'd5960,17'd5377,17'd5377,17'd5792,17'd77373,17'd77784,17'd77377,17'd78073,17'd78074,17'd77717,17'd78075,17'd77650,17'd78076,17'd78077,17'd78078,17'd77937,17'd78079,17'd78080,17'd78081,17'd77446,17'd78082,17'd77933,17'd78083,17'd78084,17'd78085,17'd78086,17'd78087,17'd76687,17'd78088,17'd78089,17'd78090,17'd76552,17'd76416,17'd76426,17'd76913,17'd77946,17'd78091,17'd78092,17'd73612,17'd71765,17'd72988,17'd78093,17'd78028,17'd130,17'd131,17'd131,17'd131,17'd1481,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd133,17'd133,17'd133,17'd1759,17'd77472,17'd5744,17'd5745,17'd76994,17'd2868,17'd78094,17'd18460,17'd78095,17'd6200,17'd78096,17'd78097,17'd8133,17'd78098,17'd78099,17'd76997,17'd78100,17'd78101,17'd32711,17'd10193,17'd10356,17'd9498,17'd78102,17'd78103,17'd36729,17'd78104,17'd38310,17'd78105,17'd8756,17'd8756,17'd8286,17'd36578,17'd46980,17'd78043,17'd7321,17'd78106,17'd33687,17'd78107,17'd78108,17'd7653,17'd5603,17'd78109,17'd5142,17'd4520,17'd52761,17'd77894,17'd24798,17'd24649,17'd5607,17'd24944,17'd25083,17'd25083,17'd78110,17'd78110,17'd78111,17'd24647,17'd4680,17'd6210,17'd4990,17'd33367,17'd33838,17'd41891,17'd5144,17'd5145,17'd6067,17'd4995,17'd4995,17'd4683,17'd4995,17'd4995,17'd4526,17'd4526,17'd4526,17'd49895,17'd49804,17'd49496,17'd49704,17'd4368,17'd55555,17'd55745,17'd49599,17'd55867,17'd38571,17'd53141,17'd56204,17'd56771,17'd78112,17'd61533,17'd60267,17'd61273,17'd78113,17'd63094,17'd3049,17'd2718,17'd65699,17'd78114,17'd55075,17'd21942,17'd58747,17'd2549,17'd78115,17'd78116,17'd78117,17'd78118,17'd34508,17'd78119,17'd77981,17'd77982,17'd78120,17'd78121,17'd78122,17'd78123,17'd78124,17'd78125,17'd78126,17'd78061,17'd77910,17'd77910,17'd78127,17'd77911,17'd78128,17'd77573,17'd78129,17'd78130,17'd77992,17'd77241,17'd77368,17'd78131,17'd78132,17'd78133,17'd77171,17'd77020,17'd76953,17'd78134,17'd77239,17'd584,17'd75376,17'd77998,17'd78065,17'd76674,17'd77097,17'd27821,17'd76390,17'd78135,17'd35347,17'd76532,17'd32408,17'd16388,17'd32726,17'd78136,17'd76820,17'd33376,17'd78137,17'd30945,17'd32560,17'd76471,17'd15742,17'd20001,17'd1543,17'd280,17'd24333,17'd182,17'd804,17'd254,17'd456,17'd78138,17'd456,17'd182,17'd20271,17'd24000,17'd400,17'd178
},
'{
17'd7046,17'd6423,17'd5510,17'd5644,17'd33216,17'd30047,17'd9959,17'd4736,17'd7042,17'd4736,17'd4244,17'd4428,17'd2935,17'd2781,17'd14,17'd15,17'd1412,17'd1412,17'd1,17'd1,17'd0,17'd0,17'd0,17'd0,17'd1,17'd1,17'd283,17'd283,17'd283,17'd3,17'd11,17'd10,17'd25,17'd23,17'd5,17'd6,17'd6,17'd6,17'd6,17'd6,17'd4,17'd4,17'd9,17'd9,17'd4,17'd4,17'd4,17'd4,17'd6,17'd6,17'd6,17'd6,17'd6,17'd6,17'd3753,17'd5205,17'd5205,17'd5205,17'd7,17'd6,17'd5,17'd24,17'd4,17'd4,17'd23,17'd23,17'd25,17'd25,17'd25,17'd21,17'd10,17'd11,17'd18,17'd4089,17'd8971,17'd8971,17'd12,17'd283,17'd650,17'd1275,17'd25,17'd25,17'd25,17'd4,17'd4,17'd6,17'd6,17'd6,17'd6,17'd5,17'd4,17'd23,17'd23,17'd23,17'd25,17'd25,17'd21,17'd21,17'd10,17'd808,17'd808,17'd25,17'd25,17'd25,17'd2933,17'd8814,17'd2423,17'd12,17'd0,17'd14,17'd1689,17'd3250,17'd7545,17'd14743,17'd15746,17'd4245,17'd4088,17'd4427,17'd5376,17'd6261,17'd78139,17'd77180,17'd77713,17'd77713,17'd77312,17'd77110,17'd77451,17'd78140,17'd5197,17'd5645,17'd5792,17'd7540,17'd77111,17'd78141,17'd78142,17'd77718,17'd77592,17'd78143,17'd77787,17'd78144,17'd78145,17'd78145,17'd78008,17'd78146,17'd78147,17'd78148,17'd78149,17'd77867,17'd78150,17'd78151,17'd78152,17'd78153,17'd78154,17'd78155,17'd78156,17'd76836,17'd78157,17'd78090,17'd76335,17'd78158,17'd76699,17'd78159,17'd74992,17'd73607,17'd72866,17'd72869,17'd71476,17'd78160,17'd78161,17'd359,17'd2698,17'd131,17'd131,17'd131,17'd1481,17'd1481,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd133,17'd1197,17'd133,17'd133,17'd134,17'd2698,17'd12875,17'd5466,17'd19294,17'd12734,17'd8903,17'd3030,17'd78162,17'd78163,17'd77952,17'd6533,17'd4500,17'd78164,17'd15703,17'd78165,17'd78166,17'd78167,17'd78168,17'd78169,17'd78170,17'd78171,17'd78172,17'd33033,17'd78173,17'd10357,17'd39005,17'd6835,17'd78174,17'd78175,17'd78176,17'd78177,17'd78178,17'd34327,17'd5752,17'd77966,17'd78179,17'd78180,17'd78181,17'd10041,17'd7820,17'd78182,17'd78183,17'd42630,17'd78184,17'd54497,17'd53506,17'd24148,17'd4680,17'd24648,17'd24797,17'd24648,17'd24797,17'd24797,17'd78111,17'd78111,17'd44845,17'd24478,17'd4676,17'd5754,17'd4189,17'd4999,17'd5145,17'd6067,17'd4682,17'd4683,17'd4840,17'd4840,17'd4995,17'd4526,17'd4526,17'd49597,17'd49597,17'd4369,17'd55351,17'd55351,17'd55555,17'd78185,17'd78186,17'd4031,17'd39020,17'd56204,17'd57348,17'd57094,17'd59608,17'd58731,17'd59233,17'd36594,17'd78187,17'd63235,17'd78188,17'd2881,17'd42475,17'd41768,17'd54874,17'd61162,17'd60148,17'd56780,17'd78189,17'd78190,17'd78191,17'd1939,17'd54331,17'd1938,17'd78192,17'd78193,17'd78194,17'd78195,17'd78196,17'd78195,17'd78197,17'd78059,17'd78198,17'd1519,17'd78199,17'd78200,17'd386,17'd77696,17'd78201,17'd77770,17'd77991,17'd78202,17'd78203,17'd77992,17'd77174,17'd77237,17'd77237,17'd77101,17'd77101,17'd77101,17'd579,17'd77433,17'd76390,17'd27821,17'd78204,17'd78204,17'd75980,17'd35618,17'd76605,17'd76605,17'd78205,17'd52108,17'd76390,17'd77432,17'd35909,17'd35618,17'd33214,17'd76603,17'd78206,17'd78207,17'd77176,17'd78208,17'd34931,17'd78207,17'd32560,17'd15874,17'd75694,17'd281,17'd589,17'd251,17'd639,17'd639,17'd965,17'd254,17'd966,17'd460,17'd253,17'd20271,17'd23489,17'd1116,17'd74929,17'd399
},
'{
17'd7883,17'd7046,17'd6423,17'd5510,17'd5644,17'd5199,17'd30047,17'd78209,17'd7042,17'd4736,17'd4244,17'd4428,17'd14743,17'd7711,17'd3750,17'd14,17'd1277,17'd19,17'd1,17'd1,17'd0,17'd0,17'd0,17'd0,17'd12,17'd3,17'd1275,17'd1275,17'd1275,17'd1275,17'd283,17'd1275,17'd25,17'd23,17'd5,17'd5,17'd6,17'd6,17'd6,17'd6,17'd4,17'd4,17'd9,17'd9,17'd4,17'd4,17'd4,17'd4,17'd4,17'd4,17'd6,17'd6,17'd6,17'd6,17'd6,17'd6,17'd6,17'd7,17'd7,17'd7,17'd4,17'd4,17'd4,17'd4,17'd23,17'd23,17'd23,17'd23,17'd25,17'd21,17'd10,17'd10,17'd283,17'd12,17'd2595,17'd15745,17'd2595,17'd466,17'd1,17'd1412,17'd650,17'd465,17'd465,17'd977,17'd9,17'd8,17'd6,17'd6,17'd6,17'd5,17'd5,17'd24,17'd23,17'd23,17'd4,17'd4,17'd21,17'd21,17'd21,17'd21,17'd21,17'd23,17'd23,17'd24,17'd284,17'd22,17'd2591,17'd1275,17'd3,17'd0,17'd1967,17'd1967,17'd1967,17'd2781,17'd2422,17'd14188,17'd34512,17'd3592,17'd4427,17'd7212,17'd7710,17'd77589,17'd78072,17'd77180,17'd78072,17'd77110,17'd7882,17'd7883,17'd6261,17'd7047,17'd7047,17'd72788,17'd78210,17'd77928,17'd78005,17'd77929,17'd77934,17'd78211,17'd77862,17'd77648,17'd78212,17'd78213,17'd78213,17'd78213,17'd78214,17'd78215,17'd78216,17'd76753,17'd78217,17'd78218,17'd78219,17'd76623,17'd78220,17'd78221,17'd78222,17'd76901,17'd78223,17'd78224,17'd78225,17'd78226,17'd77128,17'd78227,17'd75941,17'd74994,17'd75221,17'd74188,17'd76925,17'd73184,17'd77065,17'd71372,17'd720,17'd132,17'd131,17'd131,17'd130,17'd130,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd132,17'd132,17'd134,17'd135,17'd10492,17'd5744,17'd78228,17'd78229,17'd12734,17'd9900,17'd76789,17'd78230,17'd78163,17'd6533,17'd78231,17'd5133,17'd78232,17'd9061,17'd78233,17'd78234,17'd78235,17'd78236,17'd78237,17'd78238,17'd77282,17'd77481,17'd33034,17'd9903,17'd78239,17'd78240,17'd78241,17'd36881,17'd7820,17'd37687,17'd8139,17'd8603,17'd10626,17'd9366,17'd78242,17'd8449,17'd47760,17'd4665,17'd43456,17'd34497,17'd78243,17'd78244,17'd36166,17'd36022,17'd39610,17'd78184,17'd78184,17'd4522,17'd5605,17'd5606,17'd78245,17'd78246,17'd5606,17'd5606,17'd78247,17'd5755,17'd4676,17'd4523,17'd4358,17'd4834,17'd33991,17'd33838,17'd4189,17'd4999,17'd4999,17'd4525,17'd5000,17'd42181,17'd42181,17'd55454,17'd49497,17'd51844,17'd55745,17'd78186,17'd78248,17'd78249,17'd39618,17'd55748,17'd37811,17'd37564,17'd37159,17'd3542,17'd59614,17'd51576,17'd78250,17'd22430,17'd78251,17'd78252,17'd78253,17'd65698,17'd37706,17'd62334,17'd78254,17'd78255,17'd78256,17'd78257,17'd78258,17'd78259,17'd78260,17'd53597,17'd53597,17'd78261,17'd78262,17'd78263,17'd78264,17'd78265,17'd78266,17'd78267,17'd78268,17'd78269,17'd78270,17'd384,17'd78061,17'd78061,17'd77696,17'd77696,17'd78271,17'd78272,17'd77992,17'd78273,17'd77362,17'd77429,17'd78274,17'd78275,17'd78276,17'd78277,17'd77027,17'd37046,17'd77703,17'd77238,17'd76741,17'd76887,17'd76887,17'd34345,17'd36182,17'd36182,17'd35910,17'd34345,17'd77019,17'd78278,17'd27821,17'd76817,17'd77298,17'd76742,17'd34667,17'd78066,17'd76742,17'd78279,17'd78280,17'd78281,17'd76606,17'd78282,17'd32407,17'd16006,17'd75694,17'd29173,17'd16633,17'd24332,17'd24333,17'd639,17'd965,17'd254,17'd460,17'd804,17'd181,17'd252,17'd1542,17'd29442,17'd29442,17'd76157
},
'{
17'd7709,17'd7883,17'd7046,17'd6423,17'd6422,17'd5790,17'd5199,17'd30047,17'd4736,17'd3903,17'd4428,17'd6420,17'd6420,17'd4246,17'd2592,17'd1967,17'd16,17'd19,17'd1,17'd1,17'd1,17'd0,17'd0,17'd0,17'd12,17'd12,17'd806,17'd1275,17'd1275,17'd1275,17'd283,17'd1275,17'd25,17'd23,17'd5,17'd5,17'd6,17'd6,17'd6,17'd6,17'd4,17'd4,17'd9,17'd9,17'd4,17'd4,17'd4,17'd23,17'd23,17'd4,17'd6,17'd6,17'd6,17'd6,17'd6,17'd6,17'd6,17'd6,17'd7,17'd7,17'd8,17'd4,17'd4,17'd4,17'd23,17'd23,17'd23,17'd23,17'd25,17'd25,17'd10,17'd10,17'd3,17'd283,17'd1,17'd466,17'd78283,17'd77924,17'd1127,17'd1830,17'd1,17'd283,17'd650,17'd651,17'd9,17'd1413,17'd8,17'd7,17'd6,17'd5,17'd5,17'd24,17'd23,17'd23,17'd4,17'd4,17'd23,17'd21,17'd21,17'd21,17'd22,17'd22,17'd22,17'd23,17'd23,17'd23,17'd2421,17'd2591,17'd1275,17'd3,17'd1,17'd1830,17'd15,17'd3249,17'd1689,17'd27714,17'd38864,17'd3427,17'd4428,17'd4736,17'd5377,17'd6261,17'd78071,17'd77179,17'd77179,17'd77110,17'd8336,17'd8508,17'd77589,17'd77451,17'd77857,17'd8337,17'd77928,17'd77928,17'd77928,17'd77515,17'd78284,17'd78285,17'd78286,17'd78287,17'd78288,17'd76686,17'd78289,17'd78290,17'd78291,17'd78292,17'd76683,17'd78008,17'd78293,17'd78294,17'd78295,17'd78296,17'd78297,17'd78298,17'd78299,17'd78300,17'd78301,17'd78302,17'd78303,17'd78304,17'd78305,17'd78306,17'd77538,17'd76787,17'd73938,17'd73389,17'd72869,17'd71954,17'd78307,17'd67858,17'd136,17'd132,17'd132,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd134,17'd134,17'd5898,17'd76571,17'd5466,17'd3813,17'd78308,17'd9361,17'd78094,17'd77810,17'd78309,17'd17247,17'd17980,17'd78310,17'd78232,17'd78163,17'd14402,17'd78311,17'd78312,17'd78313,17'd78314,17'd9497,17'd78315,17'd32546,17'd78316,17'd77481,17'd8907,17'd12737,17'd78317,17'd78318,17'd78319,17'd37935,17'd9499,17'd8139,17'd8139,17'd78174,17'd78319,17'd8284,17'd5319,17'd4179,17'd78320,17'd78321,17'd41148,17'd78322,17'd78323,17'd78324,17'd78109,17'd78325,17'd41890,17'd4989,17'd4520,17'd4523,17'd5756,17'd5756,17'd5606,17'd5756,17'd4681,17'd4676,17'd4676,17'd4190,17'd4366,17'd4019,17'd4359,17'd4359,17'd4190,17'd4360,17'd4524,17'd49295,17'd4517,17'd4675,17'd78326,17'd78327,17'd78328,17'd78329,17'd78330,17'd78331,17'd78332,17'd55062,17'd56205,17'd52273,17'd53001,17'd52187,17'd36742,17'd78333,17'd51757,17'd78334,17'd52838,17'd78335,17'd26716,17'd64113,17'd78336,17'd54873,17'd53939,17'd78337,17'd56426,17'd78338,17'd78339,17'd78340,17'd78341,17'd78342,17'd78343,17'd54425,17'd78344,17'd78262,17'd78345,17'd78346,17'd78347,17'd78348,17'd78349,17'd78350,17'd78350,17'd78349,17'd78060,17'd78270,17'd78126,17'd78061,17'd78351,17'd78271,17'd77991,17'd77914,17'd78352,17'd78353,17'd77240,17'd78354,17'd78354,17'd77773,17'd77433,17'd78355,17'd36909,17'd37046,17'd78356,17'd77774,17'd78356,17'd78357,17'd77238,17'd77238,17'd76741,17'd36325,17'd34003,17'd77299,17'd27821,17'd27821,17'd76817,17'd78358,17'd78357,17'd78359,17'd78356,17'd37046,17'd78360,17'd78360,17'd77369,17'd35771,17'd76819,17'd77922,17'd16140,17'd29896,17'd29173,17'd15742,17'd1542,17'd24332,17'd180,17'd639,17'd965,17'd254,17'd804,17'd15240,17'd252,17'd770,17'd74929,17'd30046,17'd619,17'd16263
},
'{
17'd8508,17'd7709,17'd7883,17'd6423,17'd5375,17'd5643,17'd6421,17'd5200,17'd4427,17'd3903,17'd4428,17'd6420,17'd6420,17'd4245,17'd6584,17'd2781,17'd16,17'd18,17'd1,17'd1,17'd1,17'd1,17'd0,17'd0,17'd12,17'd12,17'd806,17'd806,17'd1275,17'd1275,17'd283,17'd1275,17'd25,17'd23,17'd24,17'd5,17'd5,17'd6,17'd6,17'd6,17'd4,17'd4,17'd9,17'd9,17'd9,17'd9,17'd23,17'd23,17'd23,17'd23,17'd4,17'd8,17'd5,17'd5,17'd6,17'd6,17'd5,17'd5,17'd6,17'd6,17'd8,17'd8,17'd4,17'd23,17'd23,17'd23,17'd23,17'd23,17'd23,17'd23,17'd21,17'd21,17'd806,17'd283,17'd1412,17'd0,17'd4247,17'd10535,17'd10535,17'd1831,17'd466,17'd13,17'd3,17'd1275,17'd2591,17'd2591,17'd2421,17'd978,17'd5,17'd5,17'd5,17'd5,17'd24,17'd24,17'd23,17'd23,17'd4,17'd23,17'd23,17'd22,17'd21,17'd21,17'd25,17'd23,17'd4,17'd23,17'd23,17'd25,17'd2591,17'd465,17'd1275,17'd283,17'd16,17'd1415,17'd1127,17'd1688,17'd2422,17'd3101,17'd6420,17'd9960,17'd71304,17'd7212,17'd5792,17'd6261,17'd7046,17'd29754,17'd78361,17'd31256,17'd30195,17'd8189,17'd8038,17'd8189,17'd77516,17'd77515,17'd77111,17'd77936,17'd8509,17'd77792,17'd78362,17'd78363,17'd78364,17'd78365,17'd78366,17'd78367,17'd76686,17'd78368,17'd78145,17'd78369,17'd77788,17'd78370,17'd78290,17'd78155,17'd78371,17'd76764,17'd78372,17'd78373,17'd78374,17'd78375,17'd78376,17'd78377,17'd78378,17'd78379,17'd75556,17'd73934,17'd73179,17'd73389,17'd71033,17'd71765,17'd72753,17'd72753,17'd141,17'd136,17'd132,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd2698,17'd76993,17'd3169,17'd6056,17'd78380,17'd78381,17'd16091,17'd78382,17'd78383,17'd78097,17'd78384,17'd17980,17'd17247,17'd78031,17'd78385,17'd78386,17'd78387,17'd78388,17'd78389,17'd78390,17'd78391,17'd8135,17'd78392,17'd78169,17'd78393,17'd12439,17'd78394,17'd78395,17'd37022,17'd78396,17'd33985,17'd40074,17'd10626,17'd8139,17'd37548,17'd5907,17'd78397,17'd33037,17'd41301,17'd78398,17'd78399,17'd78400,17'd78401,17'd3829,17'd78323,17'd4354,17'd4015,17'd41890,17'd45393,17'd33533,17'd42180,17'd33991,17'd4999,17'd34155,17'd34155,17'd4524,17'd4359,17'd43183,17'd78402,17'd48724,17'd78402,17'd78402,17'd48803,17'd48803,17'd78403,17'd4021,17'd4196,17'd4029,17'd78404,17'd78405,17'd78406,17'd39943,17'd51665,17'd39171,17'd55257,17'd53000,17'd3541,17'd78407,17'd78408,17'd52911,17'd47378,17'd3047,17'd78409,17'd41901,17'd78410,17'd2528,17'd65837,17'd56323,17'd62335,17'd2080,17'd78411,17'd53435,17'd67563,17'd78412,17'd78413,17'd78414,17'd78415,17'd78416,17'd55888,17'd2085,17'd54087,17'd78417,17'd78418,17'd78346,17'd78419,17'd78420,17'd78421,17'd78422,17'd78423,17'd1080,17'd78424,17'd78425,17'd78126,17'd78200,17'd78351,17'd77770,17'd77699,17'd77428,17'd78426,17'd77773,17'd78357,17'd77299,17'd78427,17'd77095,17'd76887,17'd76741,17'd37046,17'd77028,17'd77027,17'd77028,17'd77296,17'd78356,17'd77703,17'd77703,17'd36325,17'd36457,17'd78356,17'd77238,17'd34667,17'd36182,17'd77364,17'd76741,17'd37046,17'd77237,17'd78428,17'd78429,17'd78430,17'd77174,17'd77431,17'd75980,17'd76233,17'd16140,17'd215,17'd78431,17'd76746,17'd78432,17'd17298,17'd280,17'd15626,17'd17789,17'd965,17'd804,17'd17789,17'd15240,17'd15626,17'd17076,17'd15873,17'd30046,17'd15874,17'd32726
},
'{
17'd8508,17'd7709,17'd7883,17'd8509,17'd6423,17'd6422,17'd5643,17'd4890,17'd4426,17'd4244,17'd4428,17'd6420,17'd25384,17'd6420,17'd4733,17'd6260,17'd14,17'd18,17'd1,17'd1,17'd1,17'd1,17'd0,17'd0,17'd12,17'd12,17'd806,17'd806,17'd1275,17'd1275,17'd283,17'd1275,17'd25,17'd23,17'd24,17'd5,17'd5,17'd6,17'd6,17'd6,17'd8,17'd4,17'd9,17'd9,17'd9,17'd25,17'd23,17'd23,17'd22,17'd23,17'd4,17'd4,17'd5,17'd5,17'd5,17'd6,17'd5,17'd24,17'd5,17'd6,17'd8,17'd8,17'd4,17'd23,17'd23,17'd23,17'd23,17'd23,17'd23,17'd23,17'd21,17'd21,17'd806,17'd3,17'd0,17'd1830,17'd3249,17'd1689,17'd14070,17'd78433,17'd77924,17'd15745,17'd3430,17'd12,17'd806,17'd2933,17'd10260,17'd4242,17'd5,17'd5,17'd5,17'd5,17'd5,17'd24,17'd23,17'd23,17'd6,17'd5,17'd23,17'd23,17'd21,17'd25,17'd25,17'd25,17'd9,17'd25,17'd22,17'd22,17'd977,17'd977,17'd2591,17'd806,17'd979,17'd17,17'd4247,17'd1967,17'd2781,17'd3101,17'd25384,17'd3903,17'd4427,17'd7212,17'd77859,17'd78434,17'd6585,17'd7046,17'd7369,17'd7883,17'd77792,17'd77935,17'd78435,17'd77935,17'd77312,17'd77110,17'd77308,17'd7370,17'd7046,17'd6729,17'd78436,17'd78437,17'd78438,17'd78439,17'd78440,17'd78441,17'd78442,17'd78443,17'd78444,17'd78445,17'd78446,17'd78447,17'd78448,17'd78088,17'd78449,17'd78450,17'd78451,17'd78452,17'd78453,17'd78454,17'd78455,17'd78456,17'd78457,17'd78458,17'd77385,17'd78459,17'd78460,17'd73717,17'd73388,17'd71954,17'd72988,17'd78307,17'd67858,17'd138,17'd130,17'd131,17'd131,17'd131,17'd131,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd132,17'd135,17'd2860,17'd6055,17'd3812,17'd19294,17'd78461,17'd78462,17'd78463,17'd14826,17'd4656,17'd17247,17'd78164,17'd4342,17'd78464,17'd78465,17'd78466,17'd78467,17'd77671,17'd78468,17'd78469,17'd78470,17'd78471,17'd78472,17'd5136,17'd9635,17'd11688,17'd78473,17'd78474,17'd78475,17'd78476,17'd78477,17'd78478,17'd78479,17'd36729,17'd78175,17'd8139,17'd37935,17'd3828,17'd78480,17'd78481,17'd78482,17'd78483,17'd78484,17'd34498,17'd48548,17'd36301,17'd4511,17'd78485,17'd4185,17'd33533,17'd78486,17'd44009,17'd47470,17'd33992,17'd4189,17'd4189,17'd4515,17'd41612,17'd41892,17'd39471,17'd78487,17'd78488,17'd78489,17'd78489,17'd39775,17'd39775,17'd4023,17'd4023,17'd78490,17'd78491,17'd78492,17'd78493,17'd78494,17'd53795,17'd53357,17'd37565,17'd78495,17'd78496,17'd3365,17'd46590,17'd78497,17'd78498,17'd78499,17'd78500,17'd78501,17'd55562,17'd32879,17'd62335,17'd2227,17'd78502,17'd78503,17'd78503,17'd2227,17'd78412,17'd67806,17'd56218,17'd78504,17'd24664,17'd78505,17'd78506,17'd54087,17'd78507,17'd78418,17'd78508,17'd78509,17'd78270,17'd78510,17'd78422,17'd78423,17'd78511,17'd78425,17'd78425,17'd78200,17'd78512,17'd78513,17'd77629,17'd575,17'd77293,17'd77361,17'd77773,17'd76391,17'd77095,17'd78514,17'd78515,17'd78516,17'd396,17'd37170,17'd78517,17'd78518,17'd77704,17'd77028,17'd77103,17'd37447,17'd37046,17'd77170,17'd77020,17'd77240,17'd78359,17'd77364,17'd78519,17'd34668,17'd36325,17'd77234,17'd78520,17'd78521,17'd78522,17'd78523,17'd78524,17'd78354,17'd76072,17'd76309,17'd957,17'd74929,17'd76312,17'd78431,17'd78432,17'd17298,17'd770,17'd15626,17'd17789,17'd965,17'd965,17'd15240,17'd639,17'd15741,17'd74929,17'd435,17'd30046,17'd16497,17'd78525
}};
endmodule
