module images/frog2(output logic [17:0] rgb[0:39][0:39]);
assign rgb = '{
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd71709,17'd68123,17'd71706,17'd71316,17'd71710,17'd68123,17'd70856,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71710,17'd71677,17'd71348,17'd70861,17'd71711,17'd71333,17'd71712,17'd70856,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd71713,17'd71714,17'd71715,17'd71716,17'd71717,17'd71312,17'd71305,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71663,17'd71718,17'd71719,17'd71374,17'd71720,17'd71721,17'd68123,17'd68123,17'd70856,17'd70856,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd71722,17'd71430,17'd68123,17'd71709,17'd71723,17'd68123,17'd68123,17'd71724,17'd71725,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71726,17'd71589,17'd71727,17'd70867,17'd71117,17'd71728,17'd71269,17'd68123,17'd68123,17'd71729,17'd71730,17'd68123,17'd70856,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd71580,17'd71731,17'd71732,17'd12481,17'd71733,17'd71734,17'd71735,17'd71736,17'd70856,17'd71604,17'd71613,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd70873,17'd71646,17'd71737,17'd71258,17'd71189,17'd70903,17'd71738,17'd71739,17'd71740,17'd71741,17'd68123,17'd68123,17'd70862,17'd71742,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd71312,17'd71444,17'd68123,17'd64890,17'd71743,17'd71744,17'd7610,17'd71745,17'd71746,17'd71747,17'd71748,17'd71749,17'd71750,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71751,17'd71752,17'd70888,17'd71493,17'd70905,17'd70887,17'd71117,17'd6861,17'd61623,17'd71753,17'd71754,17'd71755,17'd68123,17'd71717,17'd70856,17'd70856,17'd71312,17'd70856,17'd70856,17'd70856,17'd71691,17'd52687,17'd71756,17'd71757,17'd71758,17'd71759,17'd71760,17'd71761,17'd71762,17'd71763,17'd15281,17'd68123,17'd71636,17'd68123,17'd70856,17'd71269,17'd71305,17'd71306,17'd71305,17'd71307
},
'{
17'd71764,17'd71765,17'd71766,17'd71413,17'd71189,17'd70886,17'd71767,17'd71102,17'd71768,17'd71769,17'd71228,17'd71770,17'd71771,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd71772,17'd71773,17'd68123,17'd11772,17'd71774,17'd24995,17'd71261,17'd71775,17'd71776,17'd71777,17'd71778,17'd71779,17'd71780,17'd3369,17'd71781,17'd70862,17'd71317,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71782,17'd71371,17'd71324,17'd71783,17'd71784,17'd71785,17'd71786,17'd71787,17'd71788,17'd71789,17'd71790,17'd71791,17'd71792,17'd71793,17'd71794,17'd71795,17'd71796,17'd71797,17'd57902,17'd71798,17'd71280,17'd71799,17'd43297,17'd71800,17'd71801,17'd71226,17'd71280,17'd71802,17'd71803,17'd14753,17'd71804,17'd71805,17'd70856,17'd71806,17'd68123,17'd68123,17'd71807,17'd71808,17'd71395,17'd71809
},
'{
17'd71782,17'd71320,17'd71810,17'd71811,17'd71812,17'd71813,17'd71814,17'd71473,17'd71815,17'd71816,17'd71817,17'd71818,17'd71819,17'd71820,17'd71821,17'd71822,17'd71823,17'd71824,17'd71825,17'd71826,17'd71827,17'd71828,17'd25331,17'd71829,17'd71329,17'd71830,17'd71831,17'd70867,17'd71832,17'd71833,17'd71834,17'd71835,17'd71836,17'd71837,17'd27796,17'd71838,17'd71839,17'd71840,17'd71841,17'd68123
},
'{
17'd68123,17'd70856,17'd68123,17'd68123,17'd71842,17'd71007,17'd71843,17'd70922,17'd71844,17'd71011,17'd71845,17'd71013,17'd71476,17'd71495,17'd71496,17'd71846,17'd71018,17'd71019,17'd71847,17'd71021,17'd71848,17'd71849,17'd71850,17'd71851,17'd71852,17'd71853,17'd71854,17'd71294,17'd71855,17'd71614,17'd71856,17'd59687,17'd71857,17'd71858,17'd9798,17'd71859,17'd71860,17'd71346,17'd70860,17'd71308
},
'{
17'd68123,17'd70856,17'd71861,17'd71862,17'd71863,17'd71864,17'd71865,17'd71866,17'd71867,17'd70887,17'd71510,17'd71868,17'd71039,17'd71040,17'd71869,17'd71144,17'd71870,17'd71511,17'd71073,17'd52897,17'd51878,17'd71045,17'd71046,17'd71871,17'd71872,17'd71873,17'd71874,17'd0,17'd68123,17'd71705,17'd71875,17'd71412,17'd71876,17'd71839,17'd71877,17'd71878,17'd71675,17'd71433,17'd71879,17'd71395
},
'{
17'd68123,17'd70856,17'd71880,17'd7978,17'd71055,17'd71056,17'd71881,17'd71058,17'd71059,17'd71060,17'd71061,17'd71062,17'd71037,17'd70953,17'd71062,17'd71063,17'd70887,17'd70887,17'd71063,17'd71062,17'd71063,17'd71062,17'd71037,17'd71062,17'd71064,17'd71882,17'd23759,17'd71883,17'd71884,17'd68123,17'd71885,17'd71886,17'd70857,17'd71310,17'd71640,17'd71412,17'd71887,17'd68123,17'd71700,17'd71306
},
'{
17'd68123,17'd70856,17'd68123,17'd71888,17'd35415,17'd31734,17'd61244,17'd61244,17'd71889,17'd71070,17'd71071,17'd71890,17'd71769,17'd71073,17'd71074,17'd71529,17'd71526,17'd38459,17'd71077,17'd52897,17'd71089,17'd71891,17'd71080,17'd71210,17'd71210,17'd71081,17'd71204,17'd71663,17'd71892,17'd68123,17'd71323,17'd71893,17'd71707,17'd68123,17'd71894,17'd71895,17'd71430,17'd71896,17'd71295,17'd71313
},
'{
17'd68123,17'd70856,17'd68123,17'd71897,17'd71898,17'd51878,17'd70887,17'd70887,17'd71088,17'd71059,17'd71079,17'd71079,17'd71059,17'd71868,17'd38114,17'd7487,17'd71091,17'd70887,17'd70887,17'd71899,17'd71240,17'd70906,17'd71900,17'd71901,17'd71240,17'd71902,17'd71903,17'd71437,17'd71702,17'd71598,17'd70852,17'd71904,17'd71905,17'd68123,17'd71906,17'd71907,17'd71908,17'd71909,17'd70861,17'd71313
},
'{
17'd68123,17'd70856,17'd71910,17'd71911,17'd71540,17'd71912,17'd71102,17'd70975,17'd70953,17'd71037,17'd71062,17'd71104,17'd70906,17'd71062,17'd70953,17'd71088,17'd71913,17'd71105,17'd61781,17'd71106,17'd71079,17'd24523,17'd71545,17'd12099,17'd71914,17'd71638,17'd71915,17'd71916,17'd71701,17'd68123,17'd71348,17'd71917,17'd71918,17'd71895,17'd71919,17'd71412,17'd71348,17'd71920,17'd71921,17'd71430
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd71922,17'd71923,17'd71856,17'd71767,17'd71171,17'd71062,17'd71106,17'd71119,17'd71924,17'd71041,17'd71555,17'd71122,17'd71123,17'd71556,17'd71556,17'd71925,17'd71127,17'd71926,17'd71927,17'd71130,17'd71928,17'd71929,17'd71930,17'd71931,17'd68123,17'd71721,17'd71727,17'd71932,17'd40204,17'd71933,17'd71860,17'd71934,17'd71935,17'd71935,17'd71245,17'd70881
},
'{
17'd71644,17'd71886,17'd71936,17'd71937,17'd71938,17'd71939,17'd71940,17'd14436,17'd71941,17'd71062,17'd38675,17'd71942,17'd71943,17'd71571,17'd71944,17'd71146,17'd71945,17'd46051,17'd71946,17'd71947,17'd71948,17'd71949,17'd71950,17'd8385,17'd71951,17'd71952,17'd71953,17'd71954,17'd71705,17'd71955,17'd71956,17'd65545,17'd71957,17'd5263,17'd71393,17'd71802,17'd71832,17'd71614,17'd71265,17'd71157
},
'{
17'd71958,17'd71959,17'd71960,17'd70857,17'd70944,17'd17616,17'd71961,17'd38149,17'd71962,17'd71963,17'd71964,17'd71965,17'd71175,17'd71648,17'd71966,17'd71587,17'd71590,17'd63495,17'd13300,17'd29694,17'd71967,17'd71579,17'd71968,17'd21726,17'd71969,17'd71264,17'd71970,17'd71971,17'd71859,17'd71170,17'd71972,17'd71687,17'd71973,17'd71811,17'd71331,17'd71974,17'd71832,17'd71226,17'd71323,17'd71975
},
'{
17'd71304,17'd71976,17'd71977,17'd71226,17'd71258,17'd71978,17'd44912,17'd71055,17'd71979,17'd71980,17'd71981,17'd71433,17'd70844,17'd71337,17'd71467,17'd71355,17'd71982,17'd71983,17'd71984,17'd71985,17'd71986,17'd70856,17'd71987,17'd71988,17'd71989,17'd71990,17'd71974,17'd71991,17'd71992,17'd71993,17'd71994,17'd11922,17'd68123,17'd71252,17'd71788,17'd71995,17'd71319,17'd71996,17'd71997,17'd71998
},
'{
17'd70854,17'd71319,17'd71239,17'd71999,17'd71189,17'd71088,17'd25924,17'd72000,17'd71878,17'd72001,17'd72002,17'd72003,17'd71691,17'd68123,17'd68123,17'd68123,17'd72004,17'd71324,17'd72005,17'd71691,17'd71296,17'd72006,17'd72007,17'd72008,17'd72009,17'd71832,17'd72010,17'd71992,17'd71769,17'd72011,17'd72012,17'd72013,17'd55754,17'd70830,17'd68123,17'd68123,17'd70862,17'd71318,17'd71252,17'd68123
},
'{
17'd71663,17'd71645,17'd71816,17'd71258,17'd70887,17'd71260,17'd70920,17'd72014,17'd71373,17'd72015,17'd72016,17'd72017,17'd72018,17'd70856,17'd71305,17'd71312,17'd70856,17'd70856,17'd68123,17'd68123,17'd70856,17'd72019,17'd71636,17'd72020,17'd72021,17'd54416,17'd71079,17'd72022,17'd72023,17'd72024,17'd72025,17'd68123,17'd68123,17'd68123,17'd71306,17'd70862,17'd71313,17'd71337,17'd72026,17'd68123
},
'{
17'd71323,17'd71009,17'd72027,17'd71977,17'd70886,17'd71267,17'd71430,17'd68123,17'd71719,17'd71310,17'd72028,17'd71466,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd72029,17'd72030,17'd72031,17'd72032,17'd72033,17'd72034,17'd16488,17'd71645,17'd68123,17'd72035,17'd70856,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71466,17'd70912,17'd71330,17'd72036,17'd71010,17'd72037,17'd68123,17'd71305,17'd71781,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd70854,17'd71548,17'd68123,17'd72038,17'd72039,17'd20596,17'd71702,17'd72035,17'd68123,17'd72040,17'd71536,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd72041,17'd70872,17'd71726,17'd71456,17'd68123,17'd70856,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd71426,17'd70862,17'd68123,17'd68123,17'd68123,17'd68123,17'd72042,17'd71306,17'd71296,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd71269,17'd71536,17'd71723,17'd68123,17'd68123,17'd68123,17'd68123,17'd70856,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd70856,17'd70856,17'd71305,17'd71269,17'd71312,17'd68123,17'd70856,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd71312,17'd71312,17'd71312,17'd70856,17'd71312,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
}};
endmodule
