module palette(output logic [7:0] palette[0:7][0:2]);
assign palette = '{'{8'd250,8'd250,8'd250},'{8'd0,8'd0,8'd0},'{8'd30,8'd70,8'd0},'{8'd0,8'd80,8'd240},'{8'd30,8'd120,8'd0},'{8'd60,8'd60,8'd60},'{8'd250,8'd230,8'd0},'{8'd0,8'd0,8'd0}};
endmodule
