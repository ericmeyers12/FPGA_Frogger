module images/frog4(output logic [17:0] rgb[0:39][0:39]);
assign rgb = '{
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68164,17'd68768,17'd70825,17'd69495,17'd69495,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd70825,17'd70826,17'd68599,17'd68800,17'd68164,17'd70827,17'd70828,17'd70829,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd70830,17'd70831,17'd70832,17'd70833,17'd70834,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd70835,17'd70836,17'd69433,17'd68599,17'd70837,17'd70838,17'd70839,17'd68123,17'd70840,17'd69495,17'd68123,17'd70841,17'd70842,17'd70843,17'd70844,17'd70845,17'd70829,17'd70844,17'd68340,17'd70845,17'd70841,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd70846,17'd70847,17'd70848,17'd70849,17'd70850,17'd70851,17'd70852,17'd70853,17'd70854,17'd70855,17'd70856,17'd70856,17'd70857,17'd70858,17'd70831,17'd68599,17'd70859,17'd70860,17'd70861,17'd68546,17'd68546,17'd70862,17'd69495,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd70863,17'd70864,17'd70865,17'd70866,17'd70867,17'd70868,17'd70869,17'd70870,17'd68768,17'd68546,17'd68123,17'd70871,17'd68123,17'd70872,17'd70873,17'd70874,17'd70875,17'd70876,17'd70877,17'd70878,17'd68546,17'd70879,17'd70880,17'd70880,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd70881,17'd70882,17'd70883,17'd70884,17'd70885,17'd70886,17'd70887,17'd70888,17'd13071,17'd70889,17'd70890,17'd70891,17'd68658,17'd70892,17'd70893,17'd70894,17'd70895,17'd70896,17'd70897,17'd70898,17'd70899,17'd69433,17'd70900,17'd68768,17'd69785,17'd69495,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd69495,17'd69495,17'd70901,17'd70902,17'd70903,17'd70904,17'd70905,17'd70906,17'd70907,17'd16367,17'd70908,17'd70909,17'd70910,17'd70911,17'd70912,17'd70876,17'd62182,17'd70913,17'd70914,17'd70915,17'd70916,17'd12926,17'd70917,17'd68164,17'd70918,17'd68820,17'd69495,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd69495,17'd69495,17'd70919,17'd70920,17'd70921,17'd70922,17'd70923,17'd70924,17'd70925,17'd70926,17'd70927,17'd70928,17'd70929,17'd70930,17'd70931,17'd41666,17'd70932,17'd44439,17'd70933,17'd58831,17'd70934,17'd70935,17'd70936,17'd70937,17'd70938,17'd70939,17'd69432,17'd70841,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd69495,17'd69785,17'd70940,17'd70941,17'd70942,17'd70943,17'd70944,17'd70945,17'd70946,17'd70944,17'd70947,17'd70948,17'd70949,17'd70950,17'd68546,17'd70951,17'd70884,17'd70952,17'd70953,17'd70954,17'd70927,17'd70955,17'd70956,17'd70957,17'd15185,17'd70958,17'd70959,17'd70960,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd69495,17'd68658,17'd68123,17'd68820,17'd70961,17'd70962,17'd70946,17'd70963,17'd70964,17'd70965,17'd70966,17'd70967,17'd70968,17'd70969,17'd70970,17'd70971,17'd70972,17'd70973,17'd70974,17'd70975,17'd70976,17'd70977,17'd70978,17'd20392,17'd29684,17'd70979,17'd70980,17'd70981,17'd70841,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd70982,17'd70983,17'd70984,17'd70985,17'd70986,17'd70987,17'd70988,17'd55866,17'd70989,17'd70990,17'd70991,17'd70992,17'd70993,17'd70994,17'd70995,17'd70996,17'd70997,17'd70998,17'd70999,17'd59193,17'd71000,17'd70975,17'd71001,17'd71002,17'd71003,17'd71004,17'd68123,17'd70841,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd41955,17'd71005,17'd71006,17'd71007,17'd71008,17'd71009,17'd71010,17'd71011,17'd71012,17'd71013,17'd71014,17'd71015,17'd71016,17'd71017,17'd71018,17'd71019,17'd71020,17'd71021,17'd71022,17'd71023,17'd71024,17'd71025,17'd71026,17'd71027,17'd71028,17'd71029,17'd71030,17'd68340,17'd70841,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd69495,17'd71031,17'd71032,17'd71033,17'd31153,17'd71034,17'd71035,17'd71036,17'd71037,17'd52616,17'd71038,17'd71039,17'd71040,17'd71041,17'd71042,17'd71043,17'd71044,17'd66641,17'd52897,17'd51878,17'd71045,17'd71046,17'd71047,17'd71048,17'd71049,17'd71050,17'd70941,17'd71051,17'd71052,17'd70841,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd69495,17'd71053,17'd71054,17'd71055,17'd71056,17'd71057,17'd71058,17'd71059,17'd71060,17'd71061,17'd71037,17'd71037,17'd71062,17'd71037,17'd70887,17'd70887,17'd70887,17'd71037,17'd71062,17'd71063,17'd71037,17'd71063,17'd71062,17'd71064,17'd71065,17'd13442,17'd71066,17'd71067,17'd69431,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd69495,17'd68658,17'd71068,17'd35415,17'd31734,17'd71069,17'd66236,17'd71070,17'd71070,17'd71071,17'd71072,17'd20462,17'd71073,17'd71074,17'd71075,17'd71076,17'd38459,17'd71077,17'd71078,17'd71079,17'd71044,17'd71080,17'd71080,17'd71080,17'd71081,17'd71082,17'd71083,17'd71084,17'd68768,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd69495,17'd68340,17'd71085,17'd71086,17'd71087,17'd70923,17'd70887,17'd71088,17'd71059,17'd71089,17'd71089,17'd71080,17'd71090,17'd71090,17'd71088,17'd71091,17'd70887,17'd71039,17'd71039,17'd71091,17'd70906,17'd70906,17'd71092,17'd71093,17'd71094,17'd52740,17'd71095,17'd71096,17'd71097,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd69495,17'd71098,17'd71099,17'd71100,17'd71101,17'd71102,17'd70975,17'd71103,17'd71037,17'd71037,17'd71104,17'd70887,17'd71103,17'd70954,17'd38114,17'd67539,17'd71105,17'd61781,17'd71106,17'd71089,17'd24523,17'd71107,17'd71108,17'd71109,17'd71110,17'd71111,17'd68546,17'd71112,17'd68599,17'd70841,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd71113,17'd71114,17'd71115,17'd71116,17'd71117,17'd71037,17'd71118,17'd71119,17'd71120,17'd71041,17'd71121,17'd71122,17'd71123,17'd71124,17'd71125,17'd71126,17'd71127,17'd71128,17'd71129,17'd71130,17'd71131,17'd71132,17'd61671,17'd71133,17'd71134,17'd71135,17'd70841,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd70841,17'd71136,17'd71137,17'd71138,17'd71139,17'd38544,17'd71140,17'd71141,17'd21195,17'd71142,17'd71143,17'd71144,17'd71145,17'd71146,17'd71147,17'd71148,17'd71149,17'd71150,17'd71151,17'd61648,17'd71152,17'd71153,17'd56552,17'd71154,17'd71155,17'd71156,17'd71157,17'd68340,17'd70841,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68340,17'd68123,17'd71158,17'd71159,17'd71160,17'd71161,17'd71162,17'd71163,17'd71164,17'd71038,17'd71165,17'd70876,17'd71166,17'd71167,17'd71168,17'd34312,17'd56074,17'd71000,17'd71169,17'd71170,17'd71171,17'd71172,17'd71173,17'd71174,17'd71175,17'd71176,17'd0,17'd70841,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68800,17'd69432,17'd68123,17'd68123,17'd68123,17'd71177,17'd71178,17'd71179,17'd71180,17'd71181,17'd71047,17'd71182,17'd71183,17'd71184,17'd71185,17'd71186,17'd71187,17'd71188,17'd71189,17'd70887,17'd71062,17'd71062,17'd71190,17'd71191,17'd71192,17'd71193,17'd68768,17'd68164,17'd70841,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68800,17'd69778,17'd71194,17'd71195,17'd71196,17'd71197,17'd71198,17'd71199,17'd71200,17'd71201,17'd71202,17'd71203,17'd71204,17'd71205,17'd71206,17'd71207,17'd55192,17'd71208,17'd71209,17'd71210,17'd71211,17'd71212,17'd71213,17'd71214,17'd26025,17'd69495,17'd71215,17'd71216,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd70827,17'd71217,17'd71218,17'd70923,17'd71219,17'd71220,17'd71221,17'd38413,17'd35415,17'd71222,17'd71223,17'd71224,17'd71162,17'd71225,17'd71226,17'd71227,17'd62943,17'd71228,17'd71229,17'd71230,17'd71231,17'd71232,17'd71233,17'd71234,17'd68599,17'd71235,17'd71236,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68700,17'd68700,17'd71237,17'd71238,17'd71239,17'd70904,17'd71240,17'd71091,17'd70866,17'd71241,17'd71242,17'd70850,17'd71243,17'd71244,17'd71245,17'd71246,17'd71247,17'd71248,17'd71249,17'd24034,17'd49844,17'd71250,17'd71112,17'd68820,17'd71251,17'd71252,17'd71253,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd71254,17'd71255,17'd71256,17'd71257,17'd71258,17'd71259,17'd71260,17'd71261,17'd71262,17'd71263,17'd71179,17'd68340,17'd68599,17'd49839,17'd71154,17'd71264,17'd71265,17'd71266,17'd71267,17'd71268,17'd68599,17'd68700,17'd71269,17'd68820,17'd71270,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd71271,17'd71272,17'd71273,17'd70867,17'd71274,17'd71258,17'd71267,17'd71275,17'd69495,17'd71276,17'd70831,17'd70879,17'd68658,17'd71277,17'd71278,17'd71279,17'd71280,17'd71281,17'd71282,17'd68599,17'd71283,17'd68768,17'd71284,17'd71285,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd71286,17'd71287,17'd71288,17'd71289,17'd71290,17'd70888,17'd71291,17'd68546,17'd70833,17'd69778,17'd69495,17'd71292,17'd68123,17'd68546,17'd68599,17'd68700,17'd71293,17'd71294,17'd71295,17'd68123,17'd68546,17'd68164,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd71296,17'd71297,17'd71298,17'd71299,17'd71300,17'd66404,17'd71301,17'd68123,17'd71302,17'd68123,17'd68123,17'd69495,17'd70856,17'd70841,17'd70853,17'd68768,17'd69432,17'd68546,17'd68123,17'd68340,17'd70841,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd70841,17'd69433,17'd70940,17'd70835,17'd71303,17'd68340,17'd70841,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd71084,17'd69432,17'd71251,17'd70841,17'd70841,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
},
'{
17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123
}};
endmodule
