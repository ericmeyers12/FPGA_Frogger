module images/car_right(output logic [17:0] rgb[0:79][0:39]);
assign rgb = '{
'{
17'd69201,17'd69202,17'd69203,17'd69204,17'd69205,17'd69206,17'd69206,17'd69206,17'd69207,17'd69208,17'd69209,17'd69210,17'd69210,17'd69211,17'd69212,17'd69212,17'd69212,17'd69212,17'd69212,17'd69212,17'd69212,17'd69212,17'd69212,17'd69213,17'd69213,17'd69214,17'd69215,17'd69216,17'd69217,17'd69218,17'd69218,17'd69219,17'd69220,17'd69221,17'd69222,17'd69223,17'd69224,17'd69225,17'd69226,17'd69227
},
'{
17'd69228,17'd69229,17'd69230,17'd69231,17'd69232,17'd69233,17'd69234,17'd69235,17'd69236,17'd69231,17'd69237,17'd69238,17'd69239,17'd69240,17'd69241,17'd69242,17'd69242,17'd69242,17'd69242,17'd69243,17'd69243,17'd69244,17'd69242,17'd69245,17'd69246,17'd69247,17'd69248,17'd69249,17'd69250,17'd69251,17'd69252,17'd69253,17'd69254,17'd69255,17'd69256,17'd69257,17'd69258,17'd69259,17'd69260,17'd69261
},
'{
17'd69262,17'd69263,17'd69264,17'd69265,17'd69266,17'd69267,17'd69268,17'd69269,17'd69267,17'd69269,17'd69270,17'd69271,17'd69272,17'd69273,17'd69274,17'd69275,17'd69275,17'd69275,17'd69275,17'd69275,17'd69275,17'd69275,17'd69275,17'd69276,17'd69277,17'd69278,17'd69279,17'd69280,17'd69281,17'd69282,17'd69269,17'd69269,17'd69267,17'd69267,17'd69269,17'd69269,17'd69267,17'd69283,17'd69284,17'd69285
},
'{
17'd69286,17'd69287,17'd69288,17'd69289,17'd69290,17'd69291,17'd69292,17'd69291,17'd69293,17'd69294,17'd69295,17'd69296,17'd69297,17'd69298,17'd69299,17'd69300,17'd69301,17'd69300,17'd69300,17'd69300,17'd69301,17'd69301,17'd69300,17'd69302,17'd69303,17'd69304,17'd69305,17'd69306,17'd69307,17'd69308,17'd69309,17'd69310,17'd69311,17'd69291,17'd69312,17'd69313,17'd69313,17'd69314,17'd69315,17'd69316
},
'{
17'd69317,17'd69318,17'd69319,17'd69320,17'd69320,17'd69321,17'd69322,17'd69323,17'd69324,17'd69325,17'd69326,17'd69327,17'd69328,17'd69322,17'd69321,17'd69329,17'd69329,17'd69329,17'd69329,17'd69329,17'd69329,17'd69329,17'd69330,17'd69331,17'd69332,17'd69332,17'd69333,17'd69334,17'd69335,17'd69336,17'd69337,17'd69338,17'd69339,17'd69340,17'd69339,17'd69341,17'd69341,17'd69330,17'd69342,17'd69343
},
'{
17'd69344,17'd69345,17'd69346,17'd69347,17'd69347,17'd69347,17'd69348,17'd69349,17'd69350,17'd69351,17'd69352,17'd69353,17'd69354,17'd69354,17'd69355,17'd69355,17'd69355,17'd69355,17'd69355,17'd69355,17'd69355,17'd69355,17'd69355,17'd69355,17'd69355,17'd69355,17'd69356,17'd69356,17'd69357,17'd69358,17'd69359,17'd69360,17'd69361,17'd69362,17'd69363,17'd69364,17'd69364,17'd69365,17'd69366,17'd69367
},
'{
17'd69368,17'd69369,17'd69370,17'd69371,17'd69372,17'd69372,17'd69373,17'd69374,17'd69375,17'd69376,17'd69377,17'd69378,17'd69379,17'd69379,17'd69380,17'd69381,17'd69382,17'd69380,17'd69380,17'd69382,17'd69382,17'd69380,17'd69383,17'd69382,17'd69380,17'd69384,17'd69385,17'd69378,17'd69386,17'd69387,17'd69388,17'd69389,17'd69390,17'd69370,17'd69391,17'd69392,17'd69392,17'd69393,17'd69394,17'd69395
},
'{
17'd69396,17'd69397,17'd69370,17'd69398,17'd69398,17'd69398,17'd69399,17'd69400,17'd69401,17'd69402,17'd69403,17'd69404,17'd69405,17'd69406,17'd69407,17'd69408,17'd69408,17'd69408,17'd69409,17'd69410,17'd69408,17'd69411,17'd69408,17'd69408,17'd69409,17'd69412,17'd69413,17'd69413,17'd69414,17'd69415,17'd69416,17'd69417,17'd69418,17'd69419,17'd69391,17'd69392,17'd69392,17'd69420,17'd69421,17'd69422
},
'{
17'd69423,17'd69424,17'd69425,17'd69426,17'd69426,17'd69427,17'd69373,17'd69428,17'd69429,17'd69430,17'd68546,17'd68340,17'd68599,17'd68123,17'd68700,17'd68546,17'd68123,17'd68599,17'd68658,17'd69431,17'd68599,17'd69432,17'd68123,17'd68123,17'd68599,17'd69433,17'd68340,17'd68123,17'd68599,17'd68123,17'd69434,17'd69435,17'd69436,17'd69419,17'd69437,17'd69438,17'd69437,17'd69439,17'd69440,17'd69441
},
'{
17'd69368,17'd69442,17'd69443,17'd69392,17'd69392,17'd69391,17'd69444,17'd69445,17'd69446,17'd69447,17'd68123,17'd69448,17'd69449,17'd69450,17'd69451,17'd68123,17'd6372,17'd69452,17'd69453,17'd69454,17'd69455,17'd69456,17'd69457,17'd46765,17'd68123,17'd69458,17'd69459,17'd69460,17'd69461,17'd69433,17'd69462,17'd69463,17'd69464,17'd69373,17'd69372,17'd69398,17'd69398,17'd69393,17'd69465,17'd69466
},
'{
17'd69368,17'd69467,17'd69468,17'd69392,17'd69392,17'd69391,17'd69444,17'd69445,17'd69469,17'd69470,17'd68123,17'd69471,17'd69472,17'd69473,17'd69474,17'd68123,17'd69475,17'd22901,17'd69476,17'd69477,17'd69478,17'd69479,17'd69480,17'd69481,17'd68123,17'd69482,17'd69483,17'd69484,17'd69485,17'd68658,17'd69486,17'd69487,17'd69488,17'd69373,17'd69372,17'd69398,17'd69398,17'd69489,17'd69490,17'd69491
},
'{
17'd69368,17'd69369,17'd69468,17'd69392,17'd69392,17'd69391,17'd69492,17'd69445,17'd69493,17'd69494,17'd68164,17'd68546,17'd68658,17'd68123,17'd69495,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68164,17'd68123,17'd68340,17'd68658,17'd68546,17'd69496,17'd69497,17'd69498,17'd69499,17'd69398,17'd69398,17'd69398,17'd69500,17'd69501,17'd69502
},
'{
17'd69368,17'd69503,17'd69425,17'd69372,17'd69398,17'd69372,17'd69504,17'd69505,17'd69506,17'd69507,17'd68123,17'd69508,17'd69509,17'd69510,17'd68123,17'd69511,17'd5611,17'd7827,17'd5611,17'd17505,17'd3989,17'd5611,17'd69512,17'd1935,17'd33031,17'd68123,17'd69513,17'd69514,17'd69515,17'd68658,17'd69516,17'd69517,17'd69518,17'd69519,17'd69520,17'd69392,17'd69392,17'd69521,17'd69522,17'd69523
},
'{
17'd69368,17'd69503,17'd69468,17'd69371,17'd69524,17'd69419,17'd69525,17'd69526,17'd69527,17'd69528,17'd68123,17'd69529,17'd69530,17'd69531,17'd68123,17'd69532,17'd69533,17'd69534,17'd69534,17'd69534,17'd69534,17'd69534,17'd69535,17'd69536,17'd69537,17'd68123,17'd69538,17'd69539,17'd69540,17'd68123,17'd69541,17'd69542,17'd69543,17'd69544,17'd69545,17'd69392,17'd69520,17'd69546,17'd69547,17'd69548
},
'{
17'd69423,17'd69503,17'd69468,17'd69398,17'd69372,17'd69419,17'd69549,17'd69550,17'd69551,17'd69393,17'd69552,17'd69553,17'd68164,17'd68340,17'd69554,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68820,17'd68123,17'd68546,17'd69555,17'd69556,17'd69557,17'd69420,17'd69558,17'd69559,17'd69542,17'd69392,17'd69392,17'd69560,17'd69561,17'd69562
},
'{
17'd69423,17'd69424,17'd69468,17'd69520,17'd69438,17'd69551,17'd69563,17'd69564,17'd69444,17'd69565,17'd69566,17'd69567,17'd69568,17'd69569,17'd68123,17'd69570,17'd69571,17'd69572,17'd69572,17'd69572,17'd69572,17'd69572,17'd69572,17'd69573,17'd69574,17'd68123,17'd69575,17'd69576,17'd69577,17'd69578,17'd69579,17'd69580,17'd69581,17'd69582,17'd69419,17'd69438,17'd69583,17'd69560,17'd69584,17'd69585
},
'{
17'd69396,17'd69586,17'd69370,17'd69392,17'd69392,17'd69521,17'd69587,17'd69588,17'd69419,17'd69398,17'd69589,17'd69590,17'd69591,17'd69592,17'd68123,17'd69593,17'd69594,17'd69594,17'd69594,17'd69594,17'd69594,17'd69594,17'd69595,17'd69594,17'd69596,17'd68123,17'd69597,17'd69598,17'd69599,17'd69600,17'd69601,17'd69443,17'd69558,17'd69602,17'd69499,17'd69603,17'd69398,17'd69489,17'd69604,17'd69605
},
'{
17'd69396,17'd69389,17'd69370,17'd69606,17'd69606,17'd69545,17'd69607,17'd69608,17'd69419,17'd69398,17'd69589,17'd69609,17'd68700,17'd69610,17'd68658,17'd69611,17'd69612,17'd69613,17'd69614,17'd69613,17'd69613,17'd69614,17'd69613,17'd69615,17'd69616,17'd69432,17'd69617,17'd69495,17'd69618,17'd69600,17'd69601,17'd69443,17'd69581,17'd69607,17'd69370,17'd69371,17'd69398,17'd69420,17'd69584,17'd69619
},
'{
17'd69396,17'd69389,17'd69370,17'd69392,17'd69520,17'd69620,17'd69543,17'd69621,17'd69622,17'd69398,17'd69623,17'd69624,17'd69625,17'd69626,17'd69433,17'd69627,17'd69628,17'd69629,17'd69629,17'd69629,17'd69629,17'd69629,17'd69629,17'd69630,17'd69627,17'd68546,17'd69631,17'd69632,17'd69633,17'd69600,17'd69601,17'd69634,17'd69635,17'd69636,17'd69637,17'd69638,17'd69371,17'd69420,17'd69639,17'd69640
},
'{
17'd69641,17'd69503,17'd69439,17'd69642,17'd69425,17'd69643,17'd69644,17'd69499,17'd69524,17'd69520,17'd69645,17'd69646,17'd69647,17'd69648,17'd68123,17'd69649,17'd69650,17'd69651,17'd69652,17'd69653,17'd69653,17'd69654,17'd69655,17'd69656,17'd69657,17'd68123,17'd69658,17'd69659,17'd69660,17'd69661,17'd69662,17'd69663,17'd69499,17'd69664,17'd69665,17'd69666,17'd69372,17'd69546,17'd69667,17'd69668
},
'{
17'd69669,17'd69503,17'd69670,17'd69671,17'd69492,17'd69672,17'd69673,17'd69373,17'd69371,17'd69391,17'd69674,17'd69675,17'd69676,17'd69677,17'd69432,17'd69678,17'd69679,17'd69680,17'd69679,17'd69679,17'd69679,17'd69679,17'd69680,17'd69679,17'd69681,17'd69433,17'd69682,17'd69683,17'd69684,17'd69685,17'd69686,17'd69371,17'd69372,17'd69673,17'd69687,17'd69666,17'd69371,17'd69560,17'd69688,17'd69689
},
'{
17'd69690,17'd69503,17'd69691,17'd69692,17'd69693,17'd69694,17'd69695,17'd69372,17'd69398,17'd69391,17'd69696,17'd69697,17'd69698,17'd69699,17'd69700,17'd69701,17'd69702,17'd69703,17'd69703,17'd69703,17'd69703,17'd69703,17'd69703,17'd69704,17'd69702,17'd69705,17'd69706,17'd69707,17'd69708,17'd69709,17'd69710,17'd69398,17'd69373,17'd69711,17'd69712,17'd69551,17'd69372,17'd69393,17'd69713,17'd69714
},
'{
17'd69396,17'd69563,17'd69715,17'd69716,17'd69717,17'd69718,17'd69719,17'd69720,17'd69721,17'd69722,17'd69723,17'd69724,17'd69725,17'd69726,17'd69727,17'd69728,17'd69729,17'd69730,17'd69730,17'd69730,17'd69730,17'd69730,17'd69730,17'd69729,17'd69731,17'd69732,17'd69733,17'd69734,17'd69735,17'd69736,17'd69737,17'd69738,17'd69739,17'd69740,17'd69741,17'd69742,17'd69524,17'd69370,17'd69743,17'd69744
},
'{
17'd69745,17'd69746,17'd69747,17'd69748,17'd69749,17'd69750,17'd69751,17'd69752,17'd69753,17'd69754,17'd69755,17'd69756,17'd69757,17'd69758,17'd69759,17'd69760,17'd69760,17'd69760,17'd69760,17'd69760,17'd69760,17'd69760,17'd69760,17'd69760,17'd69760,17'd69760,17'd69761,17'd69759,17'd69762,17'd69763,17'd69764,17'd69765,17'd69766,17'd69767,17'd69768,17'd69769,17'd69770,17'd69521,17'd69771,17'd69772
},
'{
17'd69773,17'd69774,17'd69775,17'd69776,17'd69777,17'd68546,17'd68164,17'd68800,17'd69778,17'd68123,17'd69779,17'd69780,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69782,17'd69780,17'd69780,17'd69783,17'd69784,17'd69433,17'd69785,17'd68800,17'd68800,17'd68768,17'd69786,17'd69787,17'd69393,17'd69788,17'd69789
},
'{
17'd69790,17'd69774,17'd69791,17'd69792,17'd69793,17'd68123,17'd69794,17'd69795,17'd69796,17'd68123,17'd69797,17'd69780,17'd69798,17'd69798,17'd69799,17'd69800,17'd69800,17'd69800,17'd69800,17'd69800,17'd69800,17'd69800,17'd69800,17'd69800,17'd69800,17'd69801,17'd69802,17'd69803,17'd69804,17'd69805,17'd68123,17'd69806,17'd69807,17'd69808,17'd69809,17'd69810,17'd69811,17'd69521,17'd69812,17'd69813
},
'{
17'd69773,17'd69814,17'd69815,17'd69816,17'd69817,17'd68123,17'd69818,17'd69819,17'd69820,17'd68123,17'd69821,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69822,17'd69822,17'd69823,17'd69782,17'd69824,17'd68123,17'd69825,17'd69826,17'd69827,17'd69809,17'd69828,17'd69696,17'd69439,17'd69829,17'd69830
},
'{
17'd69773,17'd69814,17'd69831,17'd69816,17'd69832,17'd68123,17'd69833,17'd69834,17'd69835,17'd68123,17'd69821,17'd69780,17'd69780,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69780,17'd69836,17'd69781,17'd69824,17'd68123,17'd69837,17'd69838,17'd69839,17'd69840,17'd69841,17'd69842,17'd69370,17'd69843,17'd69844
},
'{
17'd69773,17'd69814,17'd69815,17'd69845,17'd69846,17'd68123,17'd69847,17'd69848,17'd69835,17'd68123,17'd69821,17'd69780,17'd69780,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69780,17'd69836,17'd69781,17'd69824,17'd68123,17'd69837,17'd69838,17'd69849,17'd69840,17'd69841,17'd69842,17'd69850,17'd69851,17'd69852
},
'{
17'd69773,17'd69853,17'd69815,17'd69854,17'd69855,17'd68295,17'd69833,17'd69834,17'd69856,17'd68123,17'd69821,17'd69780,17'd69780,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69780,17'd69836,17'd69781,17'd69824,17'd68123,17'd69837,17'd69838,17'd69849,17'd69840,17'd69786,17'd69842,17'd69857,17'd69858,17'd69859
},
'{
17'd69860,17'd69861,17'd69862,17'd69863,17'd69864,17'd69865,17'd69866,17'd69867,17'd69868,17'd68123,17'd69869,17'd69780,17'd69780,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69780,17'd69836,17'd69781,17'd69824,17'd68123,17'd69837,17'd69838,17'd69849,17'd69870,17'd69786,17'd69696,17'd69499,17'd69871,17'd69872
},
'{
17'd69873,17'd69874,17'd69875,17'd69876,17'd69877,17'd69878,17'd69879,17'd69880,17'd69881,17'd68123,17'd69882,17'd69780,17'd69780,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69780,17'd69836,17'd69781,17'd69824,17'd68123,17'd69837,17'd69838,17'd69839,17'd69870,17'd69786,17'd69696,17'd69393,17'd69883,17'd69884
},
'{
17'd69885,17'd69886,17'd69887,17'd69888,17'd69889,17'd69890,17'd69891,17'd69892,17'd69893,17'd68123,17'd69882,17'd69780,17'd69780,17'd69823,17'd69894,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69823,17'd69894,17'd69823,17'd69781,17'd69781,17'd69781,17'd69780,17'd69823,17'd69780,17'd69824,17'd68123,17'd69837,17'd69838,17'd69849,17'd69870,17'd69786,17'd69696,17'd69420,17'd69895,17'd69896
},
'{
17'd69897,17'd69898,17'd69899,17'd69900,17'd69901,17'd69902,17'd69903,17'd69904,17'd69905,17'd68123,17'd69869,17'd69780,17'd69780,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69780,17'd69836,17'd69781,17'd69824,17'd68123,17'd69837,17'd69838,17'd69849,17'd69840,17'd69786,17'd69398,17'd69906,17'd69907,17'd69908
},
'{
17'd69909,17'd69910,17'd69911,17'd69912,17'd69913,17'd69914,17'd69915,17'd69916,17'd69917,17'd68123,17'd69869,17'd69780,17'd69780,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69780,17'd69836,17'd69781,17'd69824,17'd68123,17'd69837,17'd69838,17'd69849,17'd69870,17'd69841,17'd69918,17'd69489,17'd69919,17'd69920
},
'{
17'd69921,17'd69922,17'd69923,17'd69924,17'd69925,17'd69926,17'd69927,17'd69928,17'd69929,17'd68123,17'd69869,17'd69780,17'd69780,17'd69781,17'd69781,17'd69781,17'd69781,17'd69823,17'd69894,17'd69823,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69894,17'd69823,17'd69836,17'd69781,17'd69824,17'd68123,17'd69837,17'd69838,17'd69839,17'd69870,17'd69930,17'd69931,17'd69932,17'd69933,17'd69934
},
'{
17'd0,17'd69935,17'd69936,17'd69937,17'd69938,17'd69939,17'd69940,17'd69941,17'd69929,17'd68123,17'd69869,17'd69780,17'd69780,17'd69781,17'd69781,17'd69781,17'd69781,17'd69823,17'd69894,17'd69823,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69894,17'd69823,17'd69836,17'd69781,17'd69824,17'd68123,17'd69837,17'd69838,17'd69849,17'd69809,17'd69786,17'd69942,17'd69943,17'd0,17'd0
},
'{
17'd0,17'd69944,17'd69945,17'd69946,17'd69947,17'd69948,17'd69949,17'd69950,17'd69951,17'd68123,17'd69952,17'd69780,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69780,17'd69836,17'd69781,17'd69824,17'd68123,17'd69953,17'd69954,17'd69849,17'd69870,17'd69786,17'd69955,17'd69956,17'd0,17'd0
},
'{
17'd0,17'd69957,17'd69958,17'd69959,17'd69960,17'd69961,17'd69962,17'd69963,17'd69964,17'd68123,17'd69821,17'd69780,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69780,17'd69836,17'd69781,17'd69824,17'd68123,17'd69837,17'd69838,17'd69839,17'd69870,17'd69786,17'd69965,17'd69966,17'd0,17'd0
},
'{
17'd0,17'd69967,17'd69968,17'd69969,17'd69970,17'd69971,17'd69972,17'd69973,17'd69974,17'd68123,17'd69952,17'd69780,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69780,17'd69836,17'd69781,17'd69824,17'd68123,17'd69837,17'd69838,17'd69849,17'd69870,17'd69786,17'd69975,17'd69976,17'd0,17'd0
},
'{
17'd0,17'd69977,17'd69978,17'd69979,17'd69980,17'd69981,17'd69982,17'd69983,17'd69984,17'd68123,17'd69952,17'd69780,17'd69780,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69780,17'd69985,17'd69781,17'd69824,17'd68123,17'd69837,17'd69838,17'd69849,17'd69870,17'd69786,17'd69986,17'd69987,17'd0,17'd0
},
'{
17'd0,17'd69988,17'd69989,17'd69990,17'd69991,17'd69992,17'd69993,17'd69994,17'd69995,17'd68123,17'd69821,17'd69780,17'd69780,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69780,17'd69996,17'd69780,17'd69824,17'd68123,17'd69837,17'd69838,17'd69849,17'd69870,17'd69786,17'd69997,17'd69998,17'd0,17'd0
},
'{
17'd0,17'd69988,17'd69999,17'd70000,17'd70001,17'd70002,17'd70003,17'd70004,17'd70005,17'd68123,17'd69821,17'd69780,17'd69780,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69781,17'd69780,17'd69996,17'd69780,17'd69824,17'd68123,17'd69837,17'd69838,17'd69839,17'd69870,17'd69786,17'd70006,17'd69976,17'd0,17'd0
},
'{
17'd0,17'd70007,17'd70008,17'd70009,17'd70010,17'd70011,17'd70012,17'd70013,17'd70005,17'd68123,17'd69952,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69780,17'd69985,17'd69780,17'd69824,17'd68123,17'd69837,17'd69838,17'd69849,17'd69870,17'd69786,17'd70006,17'd70014,17'd0,17'd0
},
'{
17'd0,17'd70015,17'd70016,17'd70017,17'd70018,17'd70019,17'd70020,17'd70021,17'd70022,17'd68123,17'd69869,17'd69782,17'd70023,17'd70024,17'd70025,17'd70026,17'd70026,17'd69985,17'd69985,17'd69985,17'd69985,17'd69985,17'd69985,17'd69836,17'd70026,17'd69996,17'd69985,17'd70027,17'd69781,17'd69824,17'd68123,17'd70028,17'd69954,17'd69849,17'd69870,17'd69786,17'd70029,17'd70030,17'd0,17'd0
},
'{
17'd0,17'd70031,17'd70032,17'd70033,17'd70034,17'd70035,17'd70036,17'd70037,17'd70038,17'd68123,17'd69952,17'd70039,17'd69800,17'd69783,17'd69782,17'd69781,17'd69781,17'd69800,17'd69800,17'd69800,17'd69800,17'd69800,17'd69800,17'd69800,17'd69781,17'd69781,17'd69780,17'd70040,17'd69800,17'd69824,17'd68123,17'd69953,17'd69954,17'd69839,17'd69809,17'd70041,17'd70042,17'd69976,17'd0,17'd0
},
'{
17'd0,17'd70043,17'd70044,17'd70045,17'd70046,17'd70047,17'd70048,17'd70049,17'd69820,17'd68123,17'd69952,17'd69780,17'd70050,17'd70051,17'd70052,17'd70053,17'd70054,17'd70055,17'd70055,17'd70055,17'd70055,17'd70056,17'd70057,17'd70058,17'd70054,17'd70059,17'd70060,17'd70061,17'd69780,17'd69824,17'd68123,17'd69837,17'd69838,17'd69849,17'd69809,17'd70062,17'd70029,17'd69956,17'd0,17'd0
},
'{
17'd0,17'd70063,17'd70064,17'd70065,17'd70066,17'd70067,17'd70068,17'd70069,17'd70070,17'd68123,17'd69869,17'd70071,17'd70072,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68546,17'd70073,17'd69783,17'd69824,17'd68123,17'd70074,17'd70075,17'd70076,17'd69870,17'd70077,17'd70078,17'd70079,17'd0,17'd0
},
'{
17'd0,17'd70080,17'd70081,17'd70082,17'd70083,17'd70084,17'd70085,17'd70086,17'd70087,17'd70088,17'd70089,17'd70090,17'd70091,17'd70092,17'd70093,17'd70094,17'd70095,17'd70096,17'd70097,17'd70098,17'd70099,17'd70099,17'd70100,17'd70101,17'd70102,17'd70103,17'd70104,17'd70105,17'd70106,17'd69783,17'd70107,17'd70108,17'd70109,17'd70110,17'd69840,17'd70111,17'd70112,17'd70113,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70114,17'd70115,17'd70116,17'd62545,17'd70117,17'd70118,17'd70119,17'd70120,17'd69784,17'd70121,17'd70122,17'd70123,17'd70124,17'd70125,17'd70126,17'd70127,17'd70128,17'd70129,17'd70130,17'd70131,17'd70131,17'd70132,17'd70133,17'd70134,17'd70135,17'd70136,17'd70137,17'd69869,17'd70138,17'd70139,17'd70140,17'd70141,17'd70142,17'd70143,17'd70144,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70145,17'd70146,17'd70147,17'd70148,17'd70149,17'd70150,17'd69824,17'd70151,17'd68123,17'd70152,17'd70153,17'd70154,17'd70155,17'd70156,17'd70157,17'd70158,17'd70159,17'd70159,17'd70160,17'd70160,17'd70160,17'd70161,17'd70161,17'd70162,17'd70163,17'd70164,17'd70165,17'd68123,17'd70166,17'd69882,17'd70167,17'd68123,17'd68768,17'd70168,17'd70169,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70145,17'd70170,17'd70171,17'd70172,17'd70173,17'd70174,17'd70175,17'd70176,17'd70177,17'd70178,17'd70179,17'd70180,17'd70181,17'd70182,17'd70183,17'd70184,17'd68315,17'd70185,17'd70186,17'd70186,17'd70162,17'd70187,17'd70188,17'd70189,17'd70190,17'd70191,17'd70192,17'd70193,17'd70194,17'd70195,17'd70196,17'd70197,17'd70198,17'd70199,17'd70200,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70201,17'd70202,17'd70203,17'd70204,17'd70205,17'd70166,17'd70206,17'd68123,17'd70207,17'd70208,17'd70209,17'd70210,17'd70211,17'd70212,17'd70213,17'd70214,17'd68317,17'd70214,17'd70215,17'd70215,17'd70215,17'd70216,17'd70215,17'd70214,17'd70217,17'd70218,17'd70219,17'd70220,17'd68123,17'd70221,17'd70222,17'd70223,17'd70224,17'd70225,17'd70226,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70201,17'd70227,17'd70228,17'd70229,17'd70230,17'd70231,17'd68768,17'd70232,17'd70233,17'd70234,17'd70235,17'd70236,17'd70237,17'd70238,17'd70239,17'd70240,17'd70241,17'd70242,17'd70188,17'd70243,17'd70244,17'd70244,17'd70188,17'd70245,17'd70246,17'd70247,17'd70248,17'd70249,17'd70250,17'd68340,17'd70251,17'd69781,17'd70252,17'd70253,17'd70254,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70201,17'd70255,17'd70256,17'd70257,17'd70258,17'd70259,17'd70260,17'd70261,17'd70262,17'd70263,17'd70264,17'd70265,17'd70266,17'd70267,17'd70268,17'd70269,17'd70270,17'd70270,17'd70271,17'd70272,17'd70272,17'd70271,17'd70273,17'd70274,17'd70275,17'd70276,17'd70277,17'd70278,17'd70279,17'd70280,17'd70281,17'd70282,17'd69352,17'd70283,17'd70254,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70284,17'd70285,17'd70286,17'd70287,17'd70288,17'd70289,17'd70290,17'd70291,17'd70292,17'd70293,17'd70294,17'd70295,17'd70296,17'd70297,17'd70298,17'd70299,17'd70300,17'd70301,17'd70302,17'd70302,17'd70302,17'd70302,17'd70302,17'd70303,17'd70304,17'd70305,17'd70306,17'd70307,17'd70308,17'd70309,17'd70310,17'd70311,17'd70312,17'd69384,17'd70226,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70313,17'd70314,17'd70315,17'd70316,17'd70317,17'd70318,17'd70319,17'd70320,17'd70321,17'd70322,17'd70323,17'd70324,17'd70325,17'd70326,17'd70327,17'd70328,17'd70329,17'd70330,17'd70331,17'd70332,17'd70331,17'd70332,17'd70332,17'd70332,17'd70333,17'd70334,17'd70335,17'd70332,17'd70336,17'd70337,17'd68768,17'd70338,17'd70339,17'd70340,17'd70341,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70284,17'd70342,17'd70343,17'd70344,17'd70345,17'd70346,17'd70347,17'd70348,17'd70349,17'd70350,17'd70351,17'd70352,17'd70353,17'd70354,17'd70355,17'd70356,17'd70357,17'd70358,17'd70359,17'd70359,17'd70359,17'd70359,17'd70359,17'd70360,17'd70361,17'd70360,17'd70362,17'd70363,17'd70364,17'd70365,17'd70366,17'd70367,17'd70368,17'd70340,17'd70254,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70369,17'd70370,17'd70371,17'd70372,17'd70373,17'd70374,17'd70375,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68123,17'd68340,17'd68123,17'd70376,17'd70377,17'd70378,17'd70379,17'd70380,17'd70381,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70284,17'd70382,17'd70383,17'd70384,17'd70385,17'd70386,17'd70387,17'd70388,17'd70389,17'd70390,17'd70391,17'd70391,17'd70391,17'd70392,17'd70393,17'd70392,17'd70392,17'd70394,17'd70395,17'd70396,17'd70397,17'd70397,17'd70398,17'd70396,17'd70399,17'd70400,17'd70401,17'd70402,17'd70403,17'd70404,17'd70405,17'd69603,17'd69392,17'd70380,17'd70406,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70313,17'd70407,17'd70408,17'd70409,17'd70410,17'd70411,17'd70412,17'd70413,17'd70414,17'd70415,17'd70416,17'd70417,17'd70417,17'd70418,17'd70418,17'd70418,17'd70418,17'd70417,17'd70416,17'd70418,17'd70416,17'd70416,17'd70416,17'd70418,17'd70419,17'd70418,17'd70420,17'd70415,17'd69685,17'd70421,17'd70422,17'd70423,17'd69392,17'd70380,17'd70424,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70145,17'd70425,17'd70426,17'd70427,17'd70428,17'd70429,17'd70430,17'd70431,17'd70432,17'd70433,17'd70421,17'd70421,17'd69427,17'd69427,17'd69427,17'd69427,17'd69427,17'd69427,17'd69426,17'd69426,17'd69426,17'd69426,17'd69426,17'd70434,17'd69371,17'd69371,17'd70435,17'd69709,17'd70436,17'd70437,17'd70432,17'd70379,17'd69391,17'd70380,17'd70424,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70145,17'd70438,17'd70439,17'd70440,17'd70441,17'd70442,17'd70443,17'd70444,17'd69392,17'd69392,17'd70445,17'd70445,17'd69427,17'd69603,17'd70421,17'd70421,17'd70421,17'd69603,17'd70445,17'd70445,17'd70445,17'd70445,17'd70445,17'd69391,17'd69398,17'd69372,17'd69524,17'd69524,17'd69372,17'd69372,17'd69372,17'd69372,17'd70446,17'd70447,17'd70448,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70145,17'd70449,17'd70450,17'd70451,17'd70441,17'd70452,17'd70453,17'd70444,17'd70445,17'd69392,17'd69520,17'd69392,17'd69371,17'd69398,17'd69372,17'd69372,17'd69372,17'd69398,17'd69392,17'd69520,17'd69520,17'd69520,17'd69392,17'd69391,17'd69398,17'd69372,17'd69372,17'd69372,17'd69371,17'd69371,17'd69372,17'd69398,17'd70446,17'd70447,17'd70254,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70313,17'd70454,17'd70455,17'd70456,17'd70457,17'd70458,17'd70459,17'd70444,17'd70460,17'd69520,17'd69392,17'd69392,17'd69371,17'd69398,17'd69372,17'd69372,17'd69372,17'd69398,17'd69392,17'd69392,17'd69392,17'd69392,17'd69392,17'd69391,17'd69398,17'd69372,17'd69372,17'd69372,17'd69372,17'd69372,17'd69372,17'd69398,17'd70445,17'd70461,17'd70462,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70313,17'd70463,17'd70464,17'd70465,17'd70466,17'd70467,17'd70468,17'd70469,17'd70470,17'd69606,17'd69426,17'd70446,17'd69371,17'd69398,17'd69372,17'd69372,17'd69372,17'd69398,17'd69520,17'd70471,17'd70471,17'd70471,17'd70471,17'd69371,17'd69524,17'd69583,17'd69524,17'd69603,17'd69603,17'd69524,17'd69427,17'd69398,17'd69601,17'd69362,17'd70472,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70284,17'd70473,17'd70474,17'd70475,17'd70476,17'd70477,17'd70478,17'd70479,17'd70480,17'd70481,17'd69524,17'd69398,17'd69371,17'd69398,17'd69372,17'd69372,17'd69372,17'd69372,17'd69398,17'd69398,17'd69398,17'd69398,17'd69398,17'd69371,17'd69392,17'd69770,17'd69438,17'd69372,17'd69372,17'd69696,17'd69524,17'd69842,17'd69696,17'd70482,17'd70483,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70369,17'd70484,17'd70485,17'd70486,17'd70487,17'd70488,17'd70489,17'd70490,17'd70491,17'd70492,17'd70445,17'd69524,17'd69398,17'd69372,17'd69372,17'd69372,17'd69372,17'd69372,17'd69372,17'd69372,17'd69372,17'd69372,17'd69372,17'd69524,17'd70493,17'd70493,17'd70494,17'd69642,17'd69642,17'd70495,17'd70496,17'd70497,17'd70498,17'd69357,17'd70341,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70499,17'd70500,17'd70501,17'd70502,17'd70503,17'd70504,17'd70505,17'd70506,17'd70507,17'd70508,17'd70509,17'd70510,17'd69372,17'd69398,17'd69372,17'd69371,17'd69372,17'd69372,17'd69372,17'd69398,17'd69398,17'd69398,17'd69398,17'd69524,17'd70493,17'd70511,17'd70512,17'd70513,17'd70513,17'd70514,17'd70515,17'd70516,17'd69663,17'd70380,17'd70517,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70518,17'd70519,17'd70520,17'd70521,17'd70522,17'd70523,17'd70524,17'd70525,17'd70526,17'd70527,17'd70528,17'd70529,17'd69842,17'd70530,17'd69437,17'd69603,17'd70531,17'd70532,17'd69601,17'd69770,17'd69392,17'd69392,17'd69392,17'd69770,17'd70533,17'd70534,17'd70535,17'd70536,17'd70536,17'd70536,17'd70537,17'd70538,17'd69606,17'd69357,17'd70539,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70540,17'd70541,17'd70542,17'd70543,17'd70544,17'd70545,17'd70546,17'd70547,17'd70548,17'd70549,17'd70550,17'd70551,17'd70552,17'd69671,17'd70434,17'd69398,17'd69372,17'd69372,17'd69601,17'd70446,17'd69520,17'd69520,17'd69520,17'd70446,17'd70553,17'd70554,17'd70555,17'd70556,17'd70556,17'd70556,17'd70557,17'd70558,17'd69438,17'd70559,17'd70517,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70540,17'd70560,17'd70561,17'd70562,17'd70563,17'd70564,17'd70565,17'd70566,17'd70567,17'd70568,17'd70569,17'd70570,17'd70571,17'd70572,17'd70573,17'd70574,17'd70575,17'd69392,17'd70576,17'd69770,17'd69392,17'd69392,17'd69392,17'd70446,17'd70577,17'd70578,17'd70579,17'd70580,17'd70580,17'd70581,17'd70582,17'd70583,17'd70584,17'd70585,17'd70406,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70586,17'd70587,17'd70588,17'd70589,17'd70590,17'd70591,17'd70592,17'd70593,17'd70594,17'd70595,17'd70596,17'd70597,17'd70598,17'd70599,17'd70600,17'd70601,17'd70602,17'd70603,17'd70604,17'd70493,17'd69606,17'd69391,17'd69391,17'd70493,17'd70605,17'd70606,17'd70607,17'd70608,17'd70609,17'd70610,17'd70611,17'd70612,17'd70577,17'd70613,17'd70614,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70615,17'd70616,17'd70617,17'd70618,17'd70619,17'd70620,17'd70621,17'd70622,17'd70623,17'd70624,17'd70625,17'd70626,17'd70627,17'd70628,17'd70629,17'd70630,17'd70631,17'd70632,17'd70633,17'd70634,17'd70635,17'd69842,17'd69842,17'd69709,17'd70636,17'd70637,17'd70638,17'd70639,17'd70639,17'd70640,17'd70641,17'd70642,17'd70643,17'd69382,17'd70644,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd70645,17'd70646,17'd70647,17'd70648,17'd70649,17'd70650,17'd70651,17'd70652,17'd70653,17'd70654,17'd70655,17'd70656,17'd70657,17'd70658,17'd70659,17'd70660,17'd70660,17'd70661,17'd70662,17'd70663,17'd70664,17'd70665,17'd70666,17'd70667,17'd70668,17'd70669,17'd70670,17'd70671,17'd70672,17'd70673,17'd70674,17'd70675,17'd70676,17'd70677,17'd70678,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd0,17'd0,17'd70679,17'd70680,17'd70681,17'd70682,17'd70683,17'd70684,17'd70685,17'd70686,17'd70687,17'd70688,17'd70689,17'd70690,17'd70691,17'd70692,17'd70693,17'd70694,17'd70695,17'd70696,17'd70697,17'd70698,17'd70699,17'd70700,17'd69392,17'd70701,17'd70702,17'd70703,17'd70704,17'd70705,17'd70706,17'd70707,17'd70708,17'd70709,17'd70710,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd0,17'd0,17'd0,17'd70711,17'd70712,17'd70713,17'd70714,17'd70715,17'd70716,17'd70717,17'd70718,17'd70719,17'd70720,17'd70721,17'd70722,17'd70723,17'd70724,17'd70725,17'd70726,17'd70727,17'd70728,17'd70729,17'd69748,17'd70730,17'd70731,17'd70732,17'd70733,17'd70734,17'd70735,17'd70736,17'd70737,17'd70738,17'd70739,17'd41699,17'd70740,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd0,17'd0,17'd0,17'd70741,17'd70742,17'd70743,17'd70744,17'd70745,17'd70746,17'd70747,17'd70748,17'd70749,17'd70750,17'd70751,17'd70752,17'd70753,17'd70754,17'd70755,17'd70756,17'd70757,17'd70758,17'd70759,17'd70760,17'd70761,17'd70762,17'd70763,17'd70764,17'd70765,17'd70766,17'd70767,17'd70768,17'd70769,17'd70770,17'd0,17'd0,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd0,17'd0,17'd0,17'd0,17'd70771,17'd70772,17'd70773,17'd70774,17'd70775,17'd70776,17'd70777,17'd70778,17'd70779,17'd70780,17'd70781,17'd70782,17'd70783,17'd70784,17'd70785,17'd70786,17'd70787,17'd70788,17'd70789,17'd70790,17'd70791,17'd70792,17'd70793,17'd70794,17'd70795,17'd70796,17'd70797,17'd70798,17'd0,17'd0,17'd0,17'd0,17'd0,17'd0
},
'{
17'd0,17'd0,17'd0,17'd0,17'd0,17'd0,17'd70799,17'd70800,17'd70801,17'd70802,17'd70803,17'd70804,17'd70805,17'd70806,17'd70807,17'd70808,17'd70809,17'd70810,17'd70811,17'd50682,17'd70812,17'd70813,17'd70814,17'd70815,17'd70816,17'd70817,17'd70818,17'd6064,17'd70819,17'd70820,17'd70821,17'd70822,17'd70823,17'd70824,17'd0,17'd0,17'd0,17'd0,17'd0,17'd0
}};
endmodule
