module images/carright_sprite(output logic [5:0] rgb[0:79][0:39]);
assign rgb = '{
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd0,5'd0
},
'{
5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd9,5'd9,5'd11,5'd11,5'd0,5'd11,5'd0,5'd0,5'd11,5'd0,5'd0,5'd11,5'd0,5'd0,5'd11,5'd11,5'd9,5'd9,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0
},
'{
5'd0,5'd0,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd9,5'd9,5'd11,5'd11,5'd0,5'd11,5'd0,5'd0,5'd11,5'd0,5'd0,5'd11,5'd0,5'd0,5'd11,5'd11,5'd9,5'd9,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd10,5'd0,5'd0
},
'{
5'd0,5'd0,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd0,5'd0
},
'{
5'd0,5'd0,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd9,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd11,5'd11,5'd11,5'd11,5'd0,5'd11,5'd11,5'd0,5'd11,5'd11,5'd0,5'd11,5'd11,5'd0,5'd11,5'd11,5'd11,5'd11,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd11,5'd11,5'd11,5'd11,5'd0,5'd11,5'd11,5'd0,5'd11,5'd11,5'd0,5'd11,5'd11,5'd0,5'd11,5'd11,5'd11,5'd11,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd11,5'd11,5'd11,5'd0,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd0,5'd11,5'd11,5'd11,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd11,5'd11,5'd11,5'd0,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd0,5'd11,5'd11,5'd11,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd11,5'd11,5'd0,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd0,5'd11,5'd11,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd11,5'd11,5'd0,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd0,5'd11,5'd11,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd11,5'd0,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd0,5'd11,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd11,5'd0,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd0,5'd11,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd11,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd13,5'd13,5'd13,5'd12,5'd12,5'd11,5'd0,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd0,5'd11,5'd12,5'd12,5'd13,5'd13,5'd13,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd11,5'd11,5'd11,5'd0,5'd12,5'd0,5'd13,5'd13,5'd13,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd13,5'd13,5'd13,5'd0,5'd12,5'd0,5'd11,5'd11,5'd11
},
'{
5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd12,5'd12,5'd11,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd11,5'd12,5'd12,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12
},
'{
5'd12,5'd12,5'd12,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd11,5'd0,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd0,5'd11,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd12,5'd12,5'd12
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd0,5'd0,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd0,5'd0,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
}};
endmodule
